module configs_latches_0 (input clk, input reset,
    input [31:0] io_d_in,
    input [-1:0] io_configs_en,
    output reg [-1:0] io_configs_out);

endmodule


module configs_latches_1 (input clk, input reset,
    input [31:0] io_d_in,
    input [0:0] io_configs_en,
    output reg [31:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

endmodule


module configs_latches_2 (input clk, input reset,
    input [31:0] io_d_in,
    input [1:0] io_configs_en,
    output reg [63:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

endmodule


module configs_latches_3 (input clk, input reset,
    input [31:0] io_d_in,
    input [2:0] io_configs_en,
    output reg [95:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

endmodule


module configs_latches_4 (input clk, input reset,
    input [31:0] io_d_in,
    input [3:0] io_configs_en,
    output reg [127:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

endmodule


module configs_latches_5 (input clk, input reset,
    input [31:0] io_d_in,
    input [4:0] io_configs_en,
    output reg [159:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

endmodule


module configs_latches_6 (input clk, input reset,
    input [31:0] io_d_in,
    input [5:0] io_configs_en,
    output reg [191:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

endmodule


module configs_latches_7 (input clk, input reset,
    input [31:0] io_d_in,
    input [6:0] io_configs_en,
    output reg [223:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

endmodule


module configs_latches_8 (input clk, input reset,
    input [31:0] io_d_in,
    input [7:0] io_configs_en,
    output reg [255:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

endmodule


module configs_latches_9 (input clk, input reset,
    input [31:0] io_d_in,
    input [8:0] io_configs_en,
    output reg [287:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

endmodule


module configs_latches_10 (input clk, input reset,
    input [31:0] io_d_in,
    input [9:0] io_configs_en,
    output reg [319:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

endmodule


module configs_latches_11 (input clk, input reset,
    input [31:0] io_d_in,
    input [10:0] io_configs_en,
    output reg [351:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

endmodule


module configs_latches_12 (input clk, input reset,
    input [31:0] io_d_in,
    input [11:0] io_configs_en,
    output reg [383:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

endmodule


module configs_latches_13 (input clk, input reset,
    input [31:0] io_d_in,
    input [12:0] io_configs_en,
    output reg [415:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

endmodule


module configs_latches_14 (input clk, input reset,
    input [31:0] io_d_in,
    input [13:0] io_configs_en,
    output reg [447:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

endmodule


module configs_latches_15 (input clk, input reset,
    input [31:0] io_d_in,
    input [14:0] io_configs_en,
    output reg [479:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

endmodule


module configs_latches_16 (input clk, input reset,
    input [31:0] io_d_in,
    input [15:0] io_configs_en,
    output reg [511:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

endmodule


module configs_latches_17 (input clk, input reset,
    input [31:0] io_d_in,
    input [16:0] io_configs_en,
    output reg [543:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

endmodule


module configs_latches_18 (input clk, input reset,
    input [31:0] io_d_in,
    input [17:0] io_configs_en,
    output reg [575:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

endmodule


module configs_latches_19 (input clk, input reset,
    input [31:0] io_d_in,
    input [18:0] io_configs_en,
    output reg [607:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

endmodule


module configs_latches_20 (input clk, input reset,
    input [31:0] io_d_in,
    input [19:0] io_configs_en,
    output reg [639:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

endmodule


module configs_latches_21 (input clk, input reset,
    input [31:0] io_d_in,
    input [20:0] io_configs_en,
    output reg [671:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

endmodule


module configs_latches_22 (input clk, input reset,
    input [31:0] io_d_in,
    input [21:0] io_configs_en,
    output reg [703:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

endmodule


module configs_latches_23 (input clk, input reset,
    input [31:0] io_d_in,
    input [22:0] io_configs_en,
    output reg [735:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

endmodule


module configs_latches_24 (input clk, input reset,
    input [31:0] io_d_in,
    input [23:0] io_configs_en,
    output reg [767:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

endmodule


module configs_latches_25 (input clk, input reset,
    input [31:0] io_d_in,
    input [24:0] io_configs_en,
    output reg [799:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

endmodule


module configs_latches_26 (input clk, input reset,
    input [31:0] io_d_in,
    input [25:0] io_configs_en,
    output reg [831:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

endmodule


module configs_latches_27 (input clk, input reset,
    input [31:0] io_d_in,
    input [26:0] io_configs_en,
    output reg [863:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

endmodule


module configs_latches_28 (input clk, input reset,
    input [31:0] io_d_in,
    input [27:0] io_configs_en,
    output reg [895:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

endmodule


module configs_latches_29 (input clk, input reset,
    input [31:0] io_d_in,
    input [28:0] io_configs_en,
    output reg [927:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

endmodule


module configs_latches_30 (input clk, input reset,
    input [31:0] io_d_in,
    input [29:0] io_configs_en,
    output reg [959:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

endmodule


module configs_latches_31 (input clk, input reset,
    input [31:0] io_d_in,
    input [30:0] io_configs_en,
    output reg [991:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

endmodule


module configs_latches_32 (input clk, input reset,
    input [31:0] io_d_in,
    input [31:0] io_configs_en,
    output reg [1023:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

endmodule


module configs_latches_33 (input clk, input reset,
    input [31:0] io_d_in,
    input [32:0] io_configs_en,
    output reg [1055:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

endmodule


module configs_latches_34 (input clk, input reset,
    input [31:0] io_d_in,
    input [33:0] io_configs_en,
    output reg [1087:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

endmodule


module configs_latches_35 (input clk, input reset,
    input [31:0] io_d_in,
    input [34:0] io_configs_en,
    output reg [1119:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

endmodule


module configs_latches_36 (input clk, input reset,
    input [31:0] io_d_in,
    input [35:0] io_configs_en,
    output reg [1151:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

endmodule


module configs_latches_37 (input clk, input reset,
    input [31:0] io_d_in,
    input [36:0] io_configs_en,
    output reg [1183:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

endmodule


module configs_latches_38 (input clk, input reset,
    input [31:0] io_d_in,
    input [37:0] io_configs_en,
    output reg [1215:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

endmodule


module configs_latches_39 (input clk, input reset,
    input [31:0] io_d_in,
    input [38:0] io_configs_en,
    output reg [1247:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

endmodule


module configs_latches_40 (input clk, input reset,
    input [31:0] io_d_in,
    input [39:0] io_configs_en,
    output reg [1279:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

endmodule


module configs_latches_41 (input clk, input reset,
    input [31:0] io_d_in,
    input [40:0] io_configs_en,
    output reg [1311:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

endmodule


module configs_latches_42 (input clk, input reset,
    input [31:0] io_d_in,
    input [41:0] io_configs_en,
    output reg [1343:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

endmodule


module configs_latches_43 (input clk, input reset,
    input [31:0] io_d_in,
    input [42:0] io_configs_en,
    output reg [1375:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

endmodule


module configs_latches_44 (input clk, input reset,
    input [31:0] io_d_in,
    input [43:0] io_configs_en,
    output reg [1407:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

endmodule


module configs_latches_45 (input clk, input reset,
    input [31:0] io_d_in,
    input [44:0] io_configs_en,
    output reg [1439:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

endmodule


module configs_latches_46 (input clk, input reset,
    input [31:0] io_d_in,
    input [45:0] io_configs_en,
    output reg [1471:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

endmodule


module configs_latches_47 (input clk, input reset,
    input [31:0] io_d_in,
    input [46:0] io_configs_en,
    output reg [1503:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

endmodule


module configs_latches_48 (input clk, input reset,
    input [31:0] io_d_in,
    input [47:0] io_configs_en,
    output reg [1535:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

endmodule


module configs_latches_49 (input clk, input reset,
    input [31:0] io_d_in,
    input [48:0] io_configs_en,
    output reg [1567:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

endmodule


module configs_latches_50 (input clk, input reset,
    input [31:0] io_d_in,
    input [49:0] io_configs_en,
    output reg [1599:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

endmodule


module configs_latches_51 (input clk, input reset,
    input [31:0] io_d_in,
    input [50:0] io_configs_en,
    output reg [1631:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

endmodule


module configs_latches_52 (input clk, input reset,
    input [31:0] io_d_in,
    input [51:0] io_configs_en,
    output reg [1663:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

endmodule


module configs_latches_53 (input clk, input reset,
    input [31:0] io_d_in,
    input [52:0] io_configs_en,
    output reg [1695:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

endmodule


module configs_latches_54 (input clk, input reset,
    input [31:0] io_d_in,
    input [53:0] io_configs_en,
    output reg [1727:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

endmodule


module configs_latches_55 (input clk, input reset,
    input [31:0] io_d_in,
    input [54:0] io_configs_en,
    output reg [1759:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

endmodule


module configs_latches_56 (input clk, input reset,
    input [31:0] io_d_in,
    input [55:0] io_configs_en,
    output reg [1791:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

endmodule


module configs_latches_57 (input clk, input reset,
    input [31:0] io_d_in,
    input [56:0] io_configs_en,
    output reg [1823:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

endmodule


module configs_latches_58 (input clk, input reset,
    input [31:0] io_d_in,
    input [57:0] io_configs_en,
    output reg [1855:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

endmodule


module configs_latches_59 (input clk, input reset,
    input [31:0] io_d_in,
    input [58:0] io_configs_en,
    output reg [1887:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

endmodule


module configs_latches_60 (input clk, input reset,
    input [31:0] io_d_in,
    input [59:0] io_configs_en,
    output reg [1919:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

endmodule


module configs_latches_61 (input clk, input reset,
    input [31:0] io_d_in,
    input [60:0] io_configs_en,
    output reg [1951:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

endmodule


module configs_latches_62 (input clk, input reset,
    input [31:0] io_d_in,
    input [61:0] io_configs_en,
    output reg [1983:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

endmodule


module configs_latches_63 (input clk, input reset,
    input [31:0] io_d_in,
    input [62:0] io_configs_en,
    output reg [2015:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

endmodule


module configs_latches_64 (input clk, input reset,
    input [31:0] io_d_in,
    input [63:0] io_configs_en,
    output reg [2047:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

endmodule


module configs_latches_65 (input clk, input reset,
    input [31:0] io_d_in,
    input [64:0] io_configs_en,
    output reg [2079:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

endmodule


module configs_latches_66 (input clk, input reset,
    input [31:0] io_d_in,
    input [65:0] io_configs_en,
    output reg [2111:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

endmodule


module configs_latches_67 (input clk, input reset,
    input [31:0] io_d_in,
    input [66:0] io_configs_en,
    output reg [2143:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

endmodule


module configs_latches_68 (input clk, input reset,
    input [31:0] io_d_in,
    input [67:0] io_configs_en,
    output reg [2175:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

endmodule


module configs_latches_69 (input clk, input reset,
    input [31:0] io_d_in,
    input [68:0] io_configs_en,
    output reg [2207:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

endmodule


module configs_latches_70 (input clk, input reset,
    input [31:0] io_d_in,
    input [69:0] io_configs_en,
    output reg [2239:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

endmodule


module configs_latches_71 (input clk, input reset,
    input [31:0] io_d_in,
    input [70:0] io_configs_en,
    output reg [2271:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

endmodule


module configs_latches_72 (input clk, input reset,
    input [31:0] io_d_in,
    input [71:0] io_configs_en,
    output reg [2303:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

endmodule


module configs_latches_73 (input clk, input reset,
    input [31:0] io_d_in,
    input [72:0] io_configs_en,
    output reg [2335:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

endmodule


module configs_latches_74 (input clk, input reset,
    input [31:0] io_d_in,
    input [73:0] io_configs_en,
    output reg [2367:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

endmodule


module configs_latches_75 (input clk, input reset,
    input [31:0] io_d_in,
    input [74:0] io_configs_en,
    output reg [2399:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

endmodule


module configs_latches_76 (input clk, input reset,
    input [31:0] io_d_in,
    input [75:0] io_configs_en,
    output reg [2431:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

endmodule


module configs_latches_77 (input clk, input reset,
    input [31:0] io_d_in,
    input [76:0] io_configs_en,
    output reg [2463:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

endmodule


module configs_latches_78 (input clk, input reset,
    input [31:0] io_d_in,
    input [77:0] io_configs_en,
    output reg [2495:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

endmodule


module configs_latches_79 (input clk, input reset,
    input [31:0] io_d_in,
    input [78:0] io_configs_en,
    output reg [2527:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

endmodule


module configs_latches_80 (input clk, input reset,
    input [31:0] io_d_in,
    input [79:0] io_configs_en,
    output reg [2559:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

endmodule


module configs_latches_81 (input clk, input reset,
    input [31:0] io_d_in,
    input [80:0] io_configs_en,
    output reg [2591:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

endmodule


module configs_latches_82 (input clk, input reset,
    input [31:0] io_d_in,
    input [81:0] io_configs_en,
    output reg [2623:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

endmodule


module configs_latches_83 (input clk, input reset,
    input [31:0] io_d_in,
    input [82:0] io_configs_en,
    output reg [2655:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

endmodule


module configs_latches_84 (input clk, input reset,
    input [31:0] io_d_in,
    input [83:0] io_configs_en,
    output reg [2687:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

endmodule


module configs_latches_85 (input clk, input reset,
    input [31:0] io_d_in,
    input [84:0] io_configs_en,
    output reg [2719:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

endmodule


module configs_latches_86 (input clk, input reset,
    input [31:0] io_d_in,
    input [85:0] io_configs_en,
    output reg [2751:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

endmodule


module configs_latches_87 (input clk, input reset,
    input [31:0] io_d_in,
    input [86:0] io_configs_en,
    output reg [2783:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

endmodule


module configs_latches_88 (input clk, input reset,
    input [31:0] io_d_in,
    input [87:0] io_configs_en,
    output reg [2815:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

endmodule


module configs_latches_89 (input clk, input reset,
    input [31:0] io_d_in,
    input [88:0] io_configs_en,
    output reg [2847:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

endmodule


module configs_latches_90 (input clk, input reset,
    input [31:0] io_d_in,
    input [89:0] io_configs_en,
    output reg [2879:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

endmodule


module configs_latches_91 (input clk, input reset,
    input [31:0] io_d_in,
    input [90:0] io_configs_en,
    output reg [2911:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

endmodule


module configs_latches_92 (input clk, input reset,
    input [31:0] io_d_in,
    input [91:0] io_configs_en,
    output reg [2943:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

endmodule


module configs_latches_93 (input clk, input reset,
    input [31:0] io_d_in,
    input [92:0] io_configs_en,
    output reg [2975:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

endmodule


module configs_latches_94 (input clk, input reset,
    input [31:0] io_d_in,
    input [93:0] io_configs_en,
    output reg [3007:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

endmodule


module configs_latches_95 (input clk, input reset,
    input [31:0] io_d_in,
    input [94:0] io_configs_en,
    output reg [3039:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

    always @ (io_configs_en[94] or io_d_in)
        begin
             if (io_configs_en[94])
                  begin
                      io_configs_out[3039:3008] = io_d_in;
                  end
        end

endmodule


module configs_latches_96 (input clk, input reset,
    input [31:0] io_d_in,
    input [95:0] io_configs_en,
    output reg [3071:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

    always @ (io_configs_en[94] or io_d_in)
        begin
             if (io_configs_en[94])
                  begin
                      io_configs_out[3039:3008] = io_d_in;
                  end
        end

    always @ (io_configs_en[95] or io_d_in)
        begin
             if (io_configs_en[95])
                  begin
                      io_configs_out[3071:3040] = io_d_in;
                  end
        end

endmodule


module configs_latches_97 (input clk, input reset,
    input [31:0] io_d_in,
    input [96:0] io_configs_en,
    output reg [3103:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

    always @ (io_configs_en[94] or io_d_in)
        begin
             if (io_configs_en[94])
                  begin
                      io_configs_out[3039:3008] = io_d_in;
                  end
        end

    always @ (io_configs_en[95] or io_d_in)
        begin
             if (io_configs_en[95])
                  begin
                      io_configs_out[3071:3040] = io_d_in;
                  end
        end

    always @ (io_configs_en[96] or io_d_in)
        begin
             if (io_configs_en[96])
                  begin
                      io_configs_out[3103:3072] = io_d_in;
                  end
        end

endmodule


module configs_latches_98 (input clk, input reset,
    input [31:0] io_d_in,
    input [97:0] io_configs_en,
    output reg [3135:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

    always @ (io_configs_en[94] or io_d_in)
        begin
             if (io_configs_en[94])
                  begin
                      io_configs_out[3039:3008] = io_d_in;
                  end
        end

    always @ (io_configs_en[95] or io_d_in)
        begin
             if (io_configs_en[95])
                  begin
                      io_configs_out[3071:3040] = io_d_in;
                  end
        end

    always @ (io_configs_en[96] or io_d_in)
        begin
             if (io_configs_en[96])
                  begin
                      io_configs_out[3103:3072] = io_d_in;
                  end
        end

    always @ (io_configs_en[97] or io_d_in)
        begin
             if (io_configs_en[97])
                  begin
                      io_configs_out[3135:3104] = io_d_in;
                  end
        end

endmodule


module configs_latches_99 (input clk, input reset,
    input [31:0] io_d_in,
    input [98:0] io_configs_en,
    output reg [3167:0] io_configs_out);

    always @ (io_configs_en[0] or io_d_in)
        begin
             if (io_configs_en[0])
                  begin
                      io_configs_out[31:0] = io_d_in;
                  end
        end

    always @ (io_configs_en[1] or io_d_in)
        begin
             if (io_configs_en[1])
                  begin
                      io_configs_out[63:32] = io_d_in;
                  end
        end

    always @ (io_configs_en[2] or io_d_in)
        begin
             if (io_configs_en[2])
                  begin
                      io_configs_out[95:64] = io_d_in;
                  end
        end

    always @ (io_configs_en[3] or io_d_in)
        begin
             if (io_configs_en[3])
                  begin
                      io_configs_out[127:96] = io_d_in;
                  end
        end

    always @ (io_configs_en[4] or io_d_in)
        begin
             if (io_configs_en[4])
                  begin
                      io_configs_out[159:128] = io_d_in;
                  end
        end

    always @ (io_configs_en[5] or io_d_in)
        begin
             if (io_configs_en[5])
                  begin
                      io_configs_out[191:160] = io_d_in;
                  end
        end

    always @ (io_configs_en[6] or io_d_in)
        begin
             if (io_configs_en[6])
                  begin
                      io_configs_out[223:192] = io_d_in;
                  end
        end

    always @ (io_configs_en[7] or io_d_in)
        begin
             if (io_configs_en[7])
                  begin
                      io_configs_out[255:224] = io_d_in;
                  end
        end

    always @ (io_configs_en[8] or io_d_in)
        begin
             if (io_configs_en[8])
                  begin
                      io_configs_out[287:256] = io_d_in;
                  end
        end

    always @ (io_configs_en[9] or io_d_in)
        begin
             if (io_configs_en[9])
                  begin
                      io_configs_out[319:288] = io_d_in;
                  end
        end

    always @ (io_configs_en[10] or io_d_in)
        begin
             if (io_configs_en[10])
                  begin
                      io_configs_out[351:320] = io_d_in;
                  end
        end

    always @ (io_configs_en[11] or io_d_in)
        begin
             if (io_configs_en[11])
                  begin
                      io_configs_out[383:352] = io_d_in;
                  end
        end

    always @ (io_configs_en[12] or io_d_in)
        begin
             if (io_configs_en[12])
                  begin
                      io_configs_out[415:384] = io_d_in;
                  end
        end

    always @ (io_configs_en[13] or io_d_in)
        begin
             if (io_configs_en[13])
                  begin
                      io_configs_out[447:416] = io_d_in;
                  end
        end

    always @ (io_configs_en[14] or io_d_in)
        begin
             if (io_configs_en[14])
                  begin
                      io_configs_out[479:448] = io_d_in;
                  end
        end

    always @ (io_configs_en[15] or io_d_in)
        begin
             if (io_configs_en[15])
                  begin
                      io_configs_out[511:480] = io_d_in;
                  end
        end

    always @ (io_configs_en[16] or io_d_in)
        begin
             if (io_configs_en[16])
                  begin
                      io_configs_out[543:512] = io_d_in;
                  end
        end

    always @ (io_configs_en[17] or io_d_in)
        begin
             if (io_configs_en[17])
                  begin
                      io_configs_out[575:544] = io_d_in;
                  end
        end

    always @ (io_configs_en[18] or io_d_in)
        begin
             if (io_configs_en[18])
                  begin
                      io_configs_out[607:576] = io_d_in;
                  end
        end

    always @ (io_configs_en[19] or io_d_in)
        begin
             if (io_configs_en[19])
                  begin
                      io_configs_out[639:608] = io_d_in;
                  end
        end

    always @ (io_configs_en[20] or io_d_in)
        begin
             if (io_configs_en[20])
                  begin
                      io_configs_out[671:640] = io_d_in;
                  end
        end

    always @ (io_configs_en[21] or io_d_in)
        begin
             if (io_configs_en[21])
                  begin
                      io_configs_out[703:672] = io_d_in;
                  end
        end

    always @ (io_configs_en[22] or io_d_in)
        begin
             if (io_configs_en[22])
                  begin
                      io_configs_out[735:704] = io_d_in;
                  end
        end

    always @ (io_configs_en[23] or io_d_in)
        begin
             if (io_configs_en[23])
                  begin
                      io_configs_out[767:736] = io_d_in;
                  end
        end

    always @ (io_configs_en[24] or io_d_in)
        begin
             if (io_configs_en[24])
                  begin
                      io_configs_out[799:768] = io_d_in;
                  end
        end

    always @ (io_configs_en[25] or io_d_in)
        begin
             if (io_configs_en[25])
                  begin
                      io_configs_out[831:800] = io_d_in;
                  end
        end

    always @ (io_configs_en[26] or io_d_in)
        begin
             if (io_configs_en[26])
                  begin
                      io_configs_out[863:832] = io_d_in;
                  end
        end

    always @ (io_configs_en[27] or io_d_in)
        begin
             if (io_configs_en[27])
                  begin
                      io_configs_out[895:864] = io_d_in;
                  end
        end

    always @ (io_configs_en[28] or io_d_in)
        begin
             if (io_configs_en[28])
                  begin
                      io_configs_out[927:896] = io_d_in;
                  end
        end

    always @ (io_configs_en[29] or io_d_in)
        begin
             if (io_configs_en[29])
                  begin
                      io_configs_out[959:928] = io_d_in;
                  end
        end

    always @ (io_configs_en[30] or io_d_in)
        begin
             if (io_configs_en[30])
                  begin
                      io_configs_out[991:960] = io_d_in;
                  end
        end

    always @ (io_configs_en[31] or io_d_in)
        begin
             if (io_configs_en[31])
                  begin
                      io_configs_out[1023:992] = io_d_in;
                  end
        end

    always @ (io_configs_en[32] or io_d_in)
        begin
             if (io_configs_en[32])
                  begin
                      io_configs_out[1055:1024] = io_d_in;
                  end
        end

    always @ (io_configs_en[33] or io_d_in)
        begin
             if (io_configs_en[33])
                  begin
                      io_configs_out[1087:1056] = io_d_in;
                  end
        end

    always @ (io_configs_en[34] or io_d_in)
        begin
             if (io_configs_en[34])
                  begin
                      io_configs_out[1119:1088] = io_d_in;
                  end
        end

    always @ (io_configs_en[35] or io_d_in)
        begin
             if (io_configs_en[35])
                  begin
                      io_configs_out[1151:1120] = io_d_in;
                  end
        end

    always @ (io_configs_en[36] or io_d_in)
        begin
             if (io_configs_en[36])
                  begin
                      io_configs_out[1183:1152] = io_d_in;
                  end
        end

    always @ (io_configs_en[37] or io_d_in)
        begin
             if (io_configs_en[37])
                  begin
                      io_configs_out[1215:1184] = io_d_in;
                  end
        end

    always @ (io_configs_en[38] or io_d_in)
        begin
             if (io_configs_en[38])
                  begin
                      io_configs_out[1247:1216] = io_d_in;
                  end
        end

    always @ (io_configs_en[39] or io_d_in)
        begin
             if (io_configs_en[39])
                  begin
                      io_configs_out[1279:1248] = io_d_in;
                  end
        end

    always @ (io_configs_en[40] or io_d_in)
        begin
             if (io_configs_en[40])
                  begin
                      io_configs_out[1311:1280] = io_d_in;
                  end
        end

    always @ (io_configs_en[41] or io_d_in)
        begin
             if (io_configs_en[41])
                  begin
                      io_configs_out[1343:1312] = io_d_in;
                  end
        end

    always @ (io_configs_en[42] or io_d_in)
        begin
             if (io_configs_en[42])
                  begin
                      io_configs_out[1375:1344] = io_d_in;
                  end
        end

    always @ (io_configs_en[43] or io_d_in)
        begin
             if (io_configs_en[43])
                  begin
                      io_configs_out[1407:1376] = io_d_in;
                  end
        end

    always @ (io_configs_en[44] or io_d_in)
        begin
             if (io_configs_en[44])
                  begin
                      io_configs_out[1439:1408] = io_d_in;
                  end
        end

    always @ (io_configs_en[45] or io_d_in)
        begin
             if (io_configs_en[45])
                  begin
                      io_configs_out[1471:1440] = io_d_in;
                  end
        end

    always @ (io_configs_en[46] or io_d_in)
        begin
             if (io_configs_en[46])
                  begin
                      io_configs_out[1503:1472] = io_d_in;
                  end
        end

    always @ (io_configs_en[47] or io_d_in)
        begin
             if (io_configs_en[47])
                  begin
                      io_configs_out[1535:1504] = io_d_in;
                  end
        end

    always @ (io_configs_en[48] or io_d_in)
        begin
             if (io_configs_en[48])
                  begin
                      io_configs_out[1567:1536] = io_d_in;
                  end
        end

    always @ (io_configs_en[49] or io_d_in)
        begin
             if (io_configs_en[49])
                  begin
                      io_configs_out[1599:1568] = io_d_in;
                  end
        end

    always @ (io_configs_en[50] or io_d_in)
        begin
             if (io_configs_en[50])
                  begin
                      io_configs_out[1631:1600] = io_d_in;
                  end
        end

    always @ (io_configs_en[51] or io_d_in)
        begin
             if (io_configs_en[51])
                  begin
                      io_configs_out[1663:1632] = io_d_in;
                  end
        end

    always @ (io_configs_en[52] or io_d_in)
        begin
             if (io_configs_en[52])
                  begin
                      io_configs_out[1695:1664] = io_d_in;
                  end
        end

    always @ (io_configs_en[53] or io_d_in)
        begin
             if (io_configs_en[53])
                  begin
                      io_configs_out[1727:1696] = io_d_in;
                  end
        end

    always @ (io_configs_en[54] or io_d_in)
        begin
             if (io_configs_en[54])
                  begin
                      io_configs_out[1759:1728] = io_d_in;
                  end
        end

    always @ (io_configs_en[55] or io_d_in)
        begin
             if (io_configs_en[55])
                  begin
                      io_configs_out[1791:1760] = io_d_in;
                  end
        end

    always @ (io_configs_en[56] or io_d_in)
        begin
             if (io_configs_en[56])
                  begin
                      io_configs_out[1823:1792] = io_d_in;
                  end
        end

    always @ (io_configs_en[57] or io_d_in)
        begin
             if (io_configs_en[57])
                  begin
                      io_configs_out[1855:1824] = io_d_in;
                  end
        end

    always @ (io_configs_en[58] or io_d_in)
        begin
             if (io_configs_en[58])
                  begin
                      io_configs_out[1887:1856] = io_d_in;
                  end
        end

    always @ (io_configs_en[59] or io_d_in)
        begin
             if (io_configs_en[59])
                  begin
                      io_configs_out[1919:1888] = io_d_in;
                  end
        end

    always @ (io_configs_en[60] or io_d_in)
        begin
             if (io_configs_en[60])
                  begin
                      io_configs_out[1951:1920] = io_d_in;
                  end
        end

    always @ (io_configs_en[61] or io_d_in)
        begin
             if (io_configs_en[61])
                  begin
                      io_configs_out[1983:1952] = io_d_in;
                  end
        end

    always @ (io_configs_en[62] or io_d_in)
        begin
             if (io_configs_en[62])
                  begin
                      io_configs_out[2015:1984] = io_d_in;
                  end
        end

    always @ (io_configs_en[63] or io_d_in)
        begin
             if (io_configs_en[63])
                  begin
                      io_configs_out[2047:2016] = io_d_in;
                  end
        end

    always @ (io_configs_en[64] or io_d_in)
        begin
             if (io_configs_en[64])
                  begin
                      io_configs_out[2079:2048] = io_d_in;
                  end
        end

    always @ (io_configs_en[65] or io_d_in)
        begin
             if (io_configs_en[65])
                  begin
                      io_configs_out[2111:2080] = io_d_in;
                  end
        end

    always @ (io_configs_en[66] or io_d_in)
        begin
             if (io_configs_en[66])
                  begin
                      io_configs_out[2143:2112] = io_d_in;
                  end
        end

    always @ (io_configs_en[67] or io_d_in)
        begin
             if (io_configs_en[67])
                  begin
                      io_configs_out[2175:2144] = io_d_in;
                  end
        end

    always @ (io_configs_en[68] or io_d_in)
        begin
             if (io_configs_en[68])
                  begin
                      io_configs_out[2207:2176] = io_d_in;
                  end
        end

    always @ (io_configs_en[69] or io_d_in)
        begin
             if (io_configs_en[69])
                  begin
                      io_configs_out[2239:2208] = io_d_in;
                  end
        end

    always @ (io_configs_en[70] or io_d_in)
        begin
             if (io_configs_en[70])
                  begin
                      io_configs_out[2271:2240] = io_d_in;
                  end
        end

    always @ (io_configs_en[71] or io_d_in)
        begin
             if (io_configs_en[71])
                  begin
                      io_configs_out[2303:2272] = io_d_in;
                  end
        end

    always @ (io_configs_en[72] or io_d_in)
        begin
             if (io_configs_en[72])
                  begin
                      io_configs_out[2335:2304] = io_d_in;
                  end
        end

    always @ (io_configs_en[73] or io_d_in)
        begin
             if (io_configs_en[73])
                  begin
                      io_configs_out[2367:2336] = io_d_in;
                  end
        end

    always @ (io_configs_en[74] or io_d_in)
        begin
             if (io_configs_en[74])
                  begin
                      io_configs_out[2399:2368] = io_d_in;
                  end
        end

    always @ (io_configs_en[75] or io_d_in)
        begin
             if (io_configs_en[75])
                  begin
                      io_configs_out[2431:2400] = io_d_in;
                  end
        end

    always @ (io_configs_en[76] or io_d_in)
        begin
             if (io_configs_en[76])
                  begin
                      io_configs_out[2463:2432] = io_d_in;
                  end
        end

    always @ (io_configs_en[77] or io_d_in)
        begin
             if (io_configs_en[77])
                  begin
                      io_configs_out[2495:2464] = io_d_in;
                  end
        end

    always @ (io_configs_en[78] or io_d_in)
        begin
             if (io_configs_en[78])
                  begin
                      io_configs_out[2527:2496] = io_d_in;
                  end
        end

    always @ (io_configs_en[79] or io_d_in)
        begin
             if (io_configs_en[79])
                  begin
                      io_configs_out[2559:2528] = io_d_in;
                  end
        end

    always @ (io_configs_en[80] or io_d_in)
        begin
             if (io_configs_en[80])
                  begin
                      io_configs_out[2591:2560] = io_d_in;
                  end
        end

    always @ (io_configs_en[81] or io_d_in)
        begin
             if (io_configs_en[81])
                  begin
                      io_configs_out[2623:2592] = io_d_in;
                  end
        end

    always @ (io_configs_en[82] or io_d_in)
        begin
             if (io_configs_en[82])
                  begin
                      io_configs_out[2655:2624] = io_d_in;
                  end
        end

    always @ (io_configs_en[83] or io_d_in)
        begin
             if (io_configs_en[83])
                  begin
                      io_configs_out[2687:2656] = io_d_in;
                  end
        end

    always @ (io_configs_en[84] or io_d_in)
        begin
             if (io_configs_en[84])
                  begin
                      io_configs_out[2719:2688] = io_d_in;
                  end
        end

    always @ (io_configs_en[85] or io_d_in)
        begin
             if (io_configs_en[85])
                  begin
                      io_configs_out[2751:2720] = io_d_in;
                  end
        end

    always @ (io_configs_en[86] or io_d_in)
        begin
             if (io_configs_en[86])
                  begin
                      io_configs_out[2783:2752] = io_d_in;
                  end
        end

    always @ (io_configs_en[87] or io_d_in)
        begin
             if (io_configs_en[87])
                  begin
                      io_configs_out[2815:2784] = io_d_in;
                  end
        end

    always @ (io_configs_en[88] or io_d_in)
        begin
             if (io_configs_en[88])
                  begin
                      io_configs_out[2847:2816] = io_d_in;
                  end
        end

    always @ (io_configs_en[89] or io_d_in)
        begin
             if (io_configs_en[89])
                  begin
                      io_configs_out[2879:2848] = io_d_in;
                  end
        end

    always @ (io_configs_en[90] or io_d_in)
        begin
             if (io_configs_en[90])
                  begin
                      io_configs_out[2911:2880] = io_d_in;
                  end
        end

    always @ (io_configs_en[91] or io_d_in)
        begin
             if (io_configs_en[91])
                  begin
                      io_configs_out[2943:2912] = io_d_in;
                  end
        end

    always @ (io_configs_en[92] or io_d_in)
        begin
             if (io_configs_en[92])
                  begin
                      io_configs_out[2975:2944] = io_d_in;
                  end
        end

    always @ (io_configs_en[93] or io_d_in)
        begin
             if (io_configs_en[93])
                  begin
                      io_configs_out[3007:2976] = io_d_in;
                  end
        end

    always @ (io_configs_en[94] or io_d_in)
        begin
             if (io_configs_en[94])
                  begin
                      io_configs_out[3039:3008] = io_d_in;
                  end
        end

    always @ (io_configs_en[95] or io_d_in)
        begin
             if (io_configs_en[95])
                  begin
                      io_configs_out[3071:3040] = io_d_in;
                  end
        end

    always @ (io_configs_en[96] or io_d_in)
        begin
             if (io_configs_en[96])
                  begin
                      io_configs_out[3103:3072] = io_d_in;
                  end
        end

    always @ (io_configs_en[97] or io_d_in)
        begin
             if (io_configs_en[97])
                  begin
                      io_configs_out[3135:3104] = io_d_in;
                  end
        end

    always @ (io_configs_en[98] or io_d_in)
        begin
             if (io_configs_en[98])
                  begin
                      io_configs_out[3167:3136] = io_d_in;
                  end
        end

endmodule


