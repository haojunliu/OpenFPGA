module fpga(
    input [79:0] top_in,
    input [79:0] bot_in,
    input [79:0] left_in,
    input [79:0] right_in,
    output [79:0] top_out,
    output [79:0] bot_out,
    output [79:0] left_out,
    output [79:0] right_out,
    input [383:0] configs_in,
    input [266:0] configs_en,
    input ff_en, clock, rst
);

    // Interconnection Wire Declaration
    wire wire_25;
    wire wire_28;
    wire wire_31;
    wire wire_34;
    wire wire_37;
    wire wire_40;
    wire wire_43;
    wire wire_46;
    wire wire_73;
    wire wire_76;
    wire wire_79;
    wire wire_82;
    wire wire_85;
    wire wire_88;
    wire wire_91;
    wire wire_94;
    wire wire_121;
    wire wire_124;
    wire wire_127;
    wire wire_130;
    wire wire_133;
    wire wire_136;
    wire wire_139;
    wire wire_142;
    wire wire_169;
    wire wire_172;
    wire wire_175;
    wire wire_178;
    wire wire_181;
    wire wire_184;
    wire wire_187;
    wire wire_190;
    wire wire_217;
    wire wire_220;
    wire wire_223;
    wire wire_226;
    wire wire_229;
    wire wire_232;
    wire wire_235;
    wire wire_238;
    wire wire_265;
    wire wire_268;
    wire wire_271;
    wire wire_274;
    wire wire_277;
    wire wire_280;
    wire wire_283;
    wire wire_286;
    wire wire_313;
    wire wire_316;
    wire wire_319;
    wire wire_322;
    wire wire_325;
    wire wire_328;
    wire wire_331;
    wire wire_334;
    wire wire_361;
    wire wire_364;
    wire wire_367;
    wire wire_370;
    wire wire_373;
    wire wire_376;
    wire wire_379;
    wire wire_382;
    wire wire_409;
    wire wire_412;
    wire wire_415;
    wire wire_418;
    wire wire_421;
    wire wire_424;
    wire wire_427;
    wire wire_430;
    wire wire_457;
    wire wire_460;
    wire wire_463;
    wire wire_466;
    wire wire_469;
    wire wire_472;
    wire wire_475;
    wire wire_478;
    wire wire_505;
    wire wire_508;
    wire wire_511;
    wire wire_514;
    wire wire_517;
    wire wire_520;
    wire wire_523;
    wire wire_526;
    wire wire_561;
    wire wire_562;
    wire wire_563;
    wire wire_564;
    wire wire_565;
    wire wire_566;
    wire wire_567;
    wire wire_568;
    wire wire_603;
    wire wire_604;
    wire wire_605;
    wire wire_606;
    wire wire_607;
    wire wire_608;
    wire wire_609;
    wire wire_610;
    wire wire_645;
    wire wire_646;
    wire wire_647;
    wire wire_648;
    wire wire_649;
    wire wire_650;
    wire wire_651;
    wire wire_652;
    wire wire_687;
    wire wire_688;
    wire wire_689;
    wire wire_690;
    wire wire_691;
    wire wire_692;
    wire wire_693;
    wire wire_694;
    wire wire_729;
    wire wire_730;
    wire wire_731;
    wire wire_732;
    wire wire_733;
    wire wire_734;
    wire wire_735;
    wire wire_736;
    wire wire_771;
    wire wire_772;
    wire wire_773;
    wire wire_774;
    wire wire_775;
    wire wire_776;
    wire wire_777;
    wire wire_778;
    wire wire_813;
    wire wire_814;
    wire wire_815;
    wire wire_816;
    wire wire_817;
    wire wire_818;
    wire wire_819;
    wire wire_820;
    wire wire_855;
    wire wire_856;
    wire wire_857;
    wire wire_858;
    wire wire_859;
    wire wire_860;
    wire wire_861;
    wire wire_862;
    wire wire_897;
    wire wire_898;
    wire wire_899;
    wire wire_900;
    wire wire_901;
    wire wire_902;
    wire wire_903;
    wire wire_904;
    wire wire_939;
    wire wire_940;
    wire wire_941;
    wire wire_942;
    wire wire_943;
    wire wire_944;
    wire wire_945;
    wire wire_946;
    wire wire_973;
    wire wire_976;
    wire wire_979;
    wire wire_982;
    wire wire_985;
    wire wire_988;
    wire wire_991;
    wire wire_994;
    wire wire_1021;
    wire wire_1024;
    wire wire_1027;
    wire wire_1030;
    wire wire_1033;
    wire wire_1036;
    wire wire_1039;
    wire wire_1042;
    wire wire_1077;
    wire wire_1078;
    wire wire_1079;
    wire wire_1080;
    wire wire_1081;
    wire wire_1082;
    wire wire_1083;
    wire wire_1084;
    wire wire_1119;
    wire wire_1120;
    wire wire_1121;
    wire wire_1122;
    wire wire_1123;
    wire wire_1124;
    wire wire_1125;
    wire wire_1126;
    wire wire_1161;
    wire wire_1162;
    wire wire_1163;
    wire wire_1164;
    wire wire_1165;
    wire wire_1166;
    wire wire_1167;
    wire wire_1168;
    wire wire_1203;
    wire wire_1204;
    wire wire_1205;
    wire wire_1206;
    wire wire_1207;
    wire wire_1208;
    wire wire_1209;
    wire wire_1210;
    wire wire_1245;
    wire wire_1246;
    wire wire_1247;
    wire wire_1248;
    wire wire_1249;
    wire wire_1250;
    wire wire_1251;
    wire wire_1252;
    wire wire_1287;
    wire wire_1288;
    wire wire_1289;
    wire wire_1290;
    wire wire_1291;
    wire wire_1292;
    wire wire_1293;
    wire wire_1294;
    wire wire_1329;
    wire wire_1330;
    wire wire_1331;
    wire wire_1332;
    wire wire_1333;
    wire wire_1334;
    wire wire_1335;
    wire wire_1336;
    wire wire_1371;
    wire wire_1372;
    wire wire_1373;
    wire wire_1374;
    wire wire_1375;
    wire wire_1376;
    wire wire_1377;
    wire wire_1378;
    wire wire_1413;
    wire wire_1414;
    wire wire_1415;
    wire wire_1416;
    wire wire_1417;
    wire wire_1418;
    wire wire_1419;
    wire wire_1420;
    wire wire_1455;
    wire wire_1456;
    wire wire_1457;
    wire wire_1458;
    wire wire_1459;
    wire wire_1460;
    wire wire_1461;
    wire wire_1462;
    wire wire_1489;
    wire wire_1492;
    wire wire_1495;
    wire wire_1498;
    wire wire_1501;
    wire wire_1504;
    wire wire_1507;
    wire wire_1510;
    wire wire_1537;
    wire wire_1540;
    wire wire_1543;
    wire wire_1546;
    wire wire_1549;
    wire wire_1552;
    wire wire_1555;
    wire wire_1558;
    wire wire_1593;
    wire wire_1594;
    wire wire_1595;
    wire wire_1596;
    wire wire_1597;
    wire wire_1598;
    wire wire_1599;
    wire wire_1600;
    wire wire_1635;
    wire wire_1636;
    wire wire_1637;
    wire wire_1638;
    wire wire_1639;
    wire wire_1640;
    wire wire_1641;
    wire wire_1642;
    wire wire_1677;
    wire wire_1678;
    wire wire_1679;
    wire wire_1680;
    wire wire_1681;
    wire wire_1682;
    wire wire_1683;
    wire wire_1684;
    wire wire_1719;
    wire wire_1720;
    wire wire_1721;
    wire wire_1722;
    wire wire_1723;
    wire wire_1724;
    wire wire_1725;
    wire wire_1726;
    wire wire_1761;
    wire wire_1762;
    wire wire_1763;
    wire wire_1764;
    wire wire_1765;
    wire wire_1766;
    wire wire_1767;
    wire wire_1768;
    wire wire_1803;
    wire wire_1804;
    wire wire_1805;
    wire wire_1806;
    wire wire_1807;
    wire wire_1808;
    wire wire_1809;
    wire wire_1810;
    wire wire_1845;
    wire wire_1846;
    wire wire_1847;
    wire wire_1848;
    wire wire_1849;
    wire wire_1850;
    wire wire_1851;
    wire wire_1852;
    wire wire_1887;
    wire wire_1888;
    wire wire_1889;
    wire wire_1890;
    wire wire_1891;
    wire wire_1892;
    wire wire_1893;
    wire wire_1894;
    wire wire_1929;
    wire wire_1930;
    wire wire_1931;
    wire wire_1932;
    wire wire_1933;
    wire wire_1934;
    wire wire_1935;
    wire wire_1936;
    wire wire_1971;
    wire wire_1972;
    wire wire_1973;
    wire wire_1974;
    wire wire_1975;
    wire wire_1976;
    wire wire_1977;
    wire wire_1978;
    wire wire_2005;
    wire wire_2008;
    wire wire_2011;
    wire wire_2014;
    wire wire_2017;
    wire wire_2020;
    wire wire_2023;
    wire wire_2026;
    wire wire_2053;
    wire wire_2056;
    wire wire_2059;
    wire wire_2062;
    wire wire_2065;
    wire wire_2068;
    wire wire_2071;
    wire wire_2074;
    wire wire_2109;
    wire wire_2110;
    wire wire_2111;
    wire wire_2112;
    wire wire_2113;
    wire wire_2114;
    wire wire_2115;
    wire wire_2116;
    wire wire_2151;
    wire wire_2152;
    wire wire_2153;
    wire wire_2154;
    wire wire_2155;
    wire wire_2156;
    wire wire_2157;
    wire wire_2158;
    wire wire_2193;
    wire wire_2194;
    wire wire_2195;
    wire wire_2196;
    wire wire_2197;
    wire wire_2198;
    wire wire_2199;
    wire wire_2200;
    wire wire_2235;
    wire wire_2236;
    wire wire_2237;
    wire wire_2238;
    wire wire_2239;
    wire wire_2240;
    wire wire_2241;
    wire wire_2242;
    wire wire_2277;
    wire wire_2278;
    wire wire_2279;
    wire wire_2280;
    wire wire_2281;
    wire wire_2282;
    wire wire_2283;
    wire wire_2284;
    wire wire_2319;
    wire wire_2320;
    wire wire_2321;
    wire wire_2322;
    wire wire_2323;
    wire wire_2324;
    wire wire_2325;
    wire wire_2326;
    wire wire_2361;
    wire wire_2362;
    wire wire_2363;
    wire wire_2364;
    wire wire_2365;
    wire wire_2366;
    wire wire_2367;
    wire wire_2368;
    wire wire_2403;
    wire wire_2404;
    wire wire_2405;
    wire wire_2406;
    wire wire_2407;
    wire wire_2408;
    wire wire_2409;
    wire wire_2410;
    wire wire_2445;
    wire wire_2446;
    wire wire_2447;
    wire wire_2448;
    wire wire_2449;
    wire wire_2450;
    wire wire_2451;
    wire wire_2452;
    wire wire_2487;
    wire wire_2488;
    wire wire_2489;
    wire wire_2490;
    wire wire_2491;
    wire wire_2492;
    wire wire_2493;
    wire wire_2494;
    wire wire_2521;
    wire wire_2524;
    wire wire_2527;
    wire wire_2530;
    wire wire_2533;
    wire wire_2536;
    wire wire_2539;
    wire wire_2542;
    wire wire_2569;
    wire wire_2572;
    wire wire_2575;
    wire wire_2578;
    wire wire_2581;
    wire wire_2584;
    wire wire_2587;
    wire wire_2590;
    wire wire_2625;
    wire wire_2626;
    wire wire_2627;
    wire wire_2628;
    wire wire_2629;
    wire wire_2630;
    wire wire_2631;
    wire wire_2632;
    wire wire_2667;
    wire wire_2668;
    wire wire_2669;
    wire wire_2670;
    wire wire_2671;
    wire wire_2672;
    wire wire_2673;
    wire wire_2674;
    wire wire_2709;
    wire wire_2710;
    wire wire_2711;
    wire wire_2712;
    wire wire_2713;
    wire wire_2714;
    wire wire_2715;
    wire wire_2716;
    wire wire_2751;
    wire wire_2752;
    wire wire_2753;
    wire wire_2754;
    wire wire_2755;
    wire wire_2756;
    wire wire_2757;
    wire wire_2758;
    wire wire_2793;
    wire wire_2794;
    wire wire_2795;
    wire wire_2796;
    wire wire_2797;
    wire wire_2798;
    wire wire_2799;
    wire wire_2800;
    wire wire_2835;
    wire wire_2836;
    wire wire_2837;
    wire wire_2838;
    wire wire_2839;
    wire wire_2840;
    wire wire_2841;
    wire wire_2842;
    wire wire_2877;
    wire wire_2878;
    wire wire_2879;
    wire wire_2880;
    wire wire_2881;
    wire wire_2882;
    wire wire_2883;
    wire wire_2884;
    wire wire_2919;
    wire wire_2920;
    wire wire_2921;
    wire wire_2922;
    wire wire_2923;
    wire wire_2924;
    wire wire_2925;
    wire wire_2926;
    wire wire_2961;
    wire wire_2962;
    wire wire_2963;
    wire wire_2964;
    wire wire_2965;
    wire wire_2966;
    wire wire_2967;
    wire wire_2968;
    wire wire_3003;
    wire wire_3004;
    wire wire_3005;
    wire wire_3006;
    wire wire_3007;
    wire wire_3008;
    wire wire_3009;
    wire wire_3010;
    wire wire_3037;
    wire wire_3040;
    wire wire_3043;
    wire wire_3046;
    wire wire_3049;
    wire wire_3052;
    wire wire_3055;
    wire wire_3058;
    wire wire_3085;
    wire wire_3088;
    wire wire_3091;
    wire wire_3094;
    wire wire_3097;
    wire wire_3100;
    wire wire_3103;
    wire wire_3106;
    wire wire_3141;
    wire wire_3142;
    wire wire_3143;
    wire wire_3144;
    wire wire_3145;
    wire wire_3146;
    wire wire_3147;
    wire wire_3148;
    wire wire_3183;
    wire wire_3184;
    wire wire_3185;
    wire wire_3186;
    wire wire_3187;
    wire wire_3188;
    wire wire_3189;
    wire wire_3190;
    wire wire_3225;
    wire wire_3226;
    wire wire_3227;
    wire wire_3228;
    wire wire_3229;
    wire wire_3230;
    wire wire_3231;
    wire wire_3232;
    wire wire_3267;
    wire wire_3268;
    wire wire_3269;
    wire wire_3270;
    wire wire_3271;
    wire wire_3272;
    wire wire_3273;
    wire wire_3274;
    wire wire_3309;
    wire wire_3310;
    wire wire_3311;
    wire wire_3312;
    wire wire_3313;
    wire wire_3314;
    wire wire_3315;
    wire wire_3316;
    wire wire_3351;
    wire wire_3352;
    wire wire_3353;
    wire wire_3354;
    wire wire_3355;
    wire wire_3356;
    wire wire_3357;
    wire wire_3358;
    wire wire_3393;
    wire wire_3394;
    wire wire_3395;
    wire wire_3396;
    wire wire_3397;
    wire wire_3398;
    wire wire_3399;
    wire wire_3400;
    wire wire_3435;
    wire wire_3436;
    wire wire_3437;
    wire wire_3438;
    wire wire_3439;
    wire wire_3440;
    wire wire_3441;
    wire wire_3442;
    wire wire_3477;
    wire wire_3478;
    wire wire_3479;
    wire wire_3480;
    wire wire_3481;
    wire wire_3482;
    wire wire_3483;
    wire wire_3484;
    wire wire_3519;
    wire wire_3520;
    wire wire_3521;
    wire wire_3522;
    wire wire_3523;
    wire wire_3524;
    wire wire_3525;
    wire wire_3526;
    wire wire_3553;
    wire wire_3556;
    wire wire_3559;
    wire wire_3562;
    wire wire_3565;
    wire wire_3568;
    wire wire_3571;
    wire wire_3574;
    wire wire_3601;
    wire wire_3604;
    wire wire_3607;
    wire wire_3610;
    wire wire_3613;
    wire wire_3616;
    wire wire_3619;
    wire wire_3622;
    wire wire_3657;
    wire wire_3658;
    wire wire_3659;
    wire wire_3660;
    wire wire_3661;
    wire wire_3662;
    wire wire_3663;
    wire wire_3664;
    wire wire_3699;
    wire wire_3700;
    wire wire_3701;
    wire wire_3702;
    wire wire_3703;
    wire wire_3704;
    wire wire_3705;
    wire wire_3706;
    wire wire_3741;
    wire wire_3742;
    wire wire_3743;
    wire wire_3744;
    wire wire_3745;
    wire wire_3746;
    wire wire_3747;
    wire wire_3748;
    wire wire_3783;
    wire wire_3784;
    wire wire_3785;
    wire wire_3786;
    wire wire_3787;
    wire wire_3788;
    wire wire_3789;
    wire wire_3790;
    wire wire_3825;
    wire wire_3826;
    wire wire_3827;
    wire wire_3828;
    wire wire_3829;
    wire wire_3830;
    wire wire_3831;
    wire wire_3832;
    wire wire_3867;
    wire wire_3868;
    wire wire_3869;
    wire wire_3870;
    wire wire_3871;
    wire wire_3872;
    wire wire_3873;
    wire wire_3874;
    wire wire_3909;
    wire wire_3910;
    wire wire_3911;
    wire wire_3912;
    wire wire_3913;
    wire wire_3914;
    wire wire_3915;
    wire wire_3916;
    wire wire_3951;
    wire wire_3952;
    wire wire_3953;
    wire wire_3954;
    wire wire_3955;
    wire wire_3956;
    wire wire_3957;
    wire wire_3958;
    wire wire_3993;
    wire wire_3994;
    wire wire_3995;
    wire wire_3996;
    wire wire_3997;
    wire wire_3998;
    wire wire_3999;
    wire wire_4000;
    wire wire_4035;
    wire wire_4036;
    wire wire_4037;
    wire wire_4038;
    wire wire_4039;
    wire wire_4040;
    wire wire_4041;
    wire wire_4042;
    wire wire_4069;
    wire wire_4072;
    wire wire_4075;
    wire wire_4078;
    wire wire_4081;
    wire wire_4084;
    wire wire_4087;
    wire wire_4090;
    wire wire_4117;
    wire wire_4120;
    wire wire_4123;
    wire wire_4126;
    wire wire_4129;
    wire wire_4132;
    wire wire_4135;
    wire wire_4138;
    wire wire_4173;
    wire wire_4174;
    wire wire_4175;
    wire wire_4176;
    wire wire_4177;
    wire wire_4178;
    wire wire_4179;
    wire wire_4180;
    wire wire_4215;
    wire wire_4216;
    wire wire_4217;
    wire wire_4218;
    wire wire_4219;
    wire wire_4220;
    wire wire_4221;
    wire wire_4222;
    wire wire_4257;
    wire wire_4258;
    wire wire_4259;
    wire wire_4260;
    wire wire_4261;
    wire wire_4262;
    wire wire_4263;
    wire wire_4264;
    wire wire_4299;
    wire wire_4300;
    wire wire_4301;
    wire wire_4302;
    wire wire_4303;
    wire wire_4304;
    wire wire_4305;
    wire wire_4306;
    wire wire_4341;
    wire wire_4342;
    wire wire_4343;
    wire wire_4344;
    wire wire_4345;
    wire wire_4346;
    wire wire_4347;
    wire wire_4348;
    wire wire_4383;
    wire wire_4384;
    wire wire_4385;
    wire wire_4386;
    wire wire_4387;
    wire wire_4388;
    wire wire_4389;
    wire wire_4390;
    wire wire_4425;
    wire wire_4426;
    wire wire_4427;
    wire wire_4428;
    wire wire_4429;
    wire wire_4430;
    wire wire_4431;
    wire wire_4432;
    wire wire_4467;
    wire wire_4468;
    wire wire_4469;
    wire wire_4470;
    wire wire_4471;
    wire wire_4472;
    wire wire_4473;
    wire wire_4474;
    wire wire_4509;
    wire wire_4510;
    wire wire_4511;
    wire wire_4512;
    wire wire_4513;
    wire wire_4514;
    wire wire_4515;
    wire wire_4516;
    wire wire_4551;
    wire wire_4552;
    wire wire_4553;
    wire wire_4554;
    wire wire_4555;
    wire wire_4556;
    wire wire_4557;
    wire wire_4558;
    wire wire_4585;
    wire wire_4588;
    wire wire_4591;
    wire wire_4594;
    wire wire_4597;
    wire wire_4600;
    wire wire_4603;
    wire wire_4606;
    wire wire_4633;
    wire wire_4636;
    wire wire_4639;
    wire wire_4642;
    wire wire_4645;
    wire wire_4648;
    wire wire_4651;
    wire wire_4654;
    wire wire_4689;
    wire wire_4690;
    wire wire_4691;
    wire wire_4692;
    wire wire_4693;
    wire wire_4694;
    wire wire_4695;
    wire wire_4696;
    wire wire_4731;
    wire wire_4732;
    wire wire_4733;
    wire wire_4734;
    wire wire_4735;
    wire wire_4736;
    wire wire_4737;
    wire wire_4738;
    wire wire_4773;
    wire wire_4774;
    wire wire_4775;
    wire wire_4776;
    wire wire_4777;
    wire wire_4778;
    wire wire_4779;
    wire wire_4780;
    wire wire_4815;
    wire wire_4816;
    wire wire_4817;
    wire wire_4818;
    wire wire_4819;
    wire wire_4820;
    wire wire_4821;
    wire wire_4822;
    wire wire_4857;
    wire wire_4858;
    wire wire_4859;
    wire wire_4860;
    wire wire_4861;
    wire wire_4862;
    wire wire_4863;
    wire wire_4864;
    wire wire_4899;
    wire wire_4900;
    wire wire_4901;
    wire wire_4902;
    wire wire_4903;
    wire wire_4904;
    wire wire_4905;
    wire wire_4906;
    wire wire_4941;
    wire wire_4942;
    wire wire_4943;
    wire wire_4944;
    wire wire_4945;
    wire wire_4946;
    wire wire_4947;
    wire wire_4948;
    wire wire_4983;
    wire wire_4984;
    wire wire_4985;
    wire wire_4986;
    wire wire_4987;
    wire wire_4988;
    wire wire_4989;
    wire wire_4990;
    wire wire_5025;
    wire wire_5026;
    wire wire_5027;
    wire wire_5028;
    wire wire_5029;
    wire wire_5030;
    wire wire_5031;
    wire wire_5032;
    wire wire_5067;
    wire wire_5068;
    wire wire_5069;
    wire wire_5070;
    wire wire_5071;
    wire wire_5072;
    wire wire_5073;
    wire wire_5074;
    wire wire_5101;
    wire wire_5104;
    wire wire_5107;
    wire wire_5110;
    wire wire_5113;
    wire wire_5116;
    wire wire_5119;
    wire wire_5122;
    wire wire_5149;
    wire wire_5152;
    wire wire_5155;
    wire wire_5158;
    wire wire_5161;
    wire wire_5164;
    wire wire_5167;
    wire wire_5170;
    wire wire_5205;
    wire wire_5206;
    wire wire_5207;
    wire wire_5208;
    wire wire_5209;
    wire wire_5210;
    wire wire_5211;
    wire wire_5212;
    wire wire_5247;
    wire wire_5248;
    wire wire_5249;
    wire wire_5250;
    wire wire_5251;
    wire wire_5252;
    wire wire_5253;
    wire wire_5254;
    wire wire_5289;
    wire wire_5290;
    wire wire_5291;
    wire wire_5292;
    wire wire_5293;
    wire wire_5294;
    wire wire_5295;
    wire wire_5296;
    wire wire_5331;
    wire wire_5332;
    wire wire_5333;
    wire wire_5334;
    wire wire_5335;
    wire wire_5336;
    wire wire_5337;
    wire wire_5338;
    wire wire_5373;
    wire wire_5374;
    wire wire_5375;
    wire wire_5376;
    wire wire_5377;
    wire wire_5378;
    wire wire_5379;
    wire wire_5380;
    wire wire_5415;
    wire wire_5416;
    wire wire_5417;
    wire wire_5418;
    wire wire_5419;
    wire wire_5420;
    wire wire_5421;
    wire wire_5422;
    wire wire_5457;
    wire wire_5458;
    wire wire_5459;
    wire wire_5460;
    wire wire_5461;
    wire wire_5462;
    wire wire_5463;
    wire wire_5464;
    wire wire_5499;
    wire wire_5500;
    wire wire_5501;
    wire wire_5502;
    wire wire_5503;
    wire wire_5504;
    wire wire_5505;
    wire wire_5506;
    wire wire_5541;
    wire wire_5542;
    wire wire_5543;
    wire wire_5544;
    wire wire_5545;
    wire wire_5546;
    wire wire_5547;
    wire wire_5548;
    wire wire_5583;
    wire wire_5584;
    wire wire_5585;
    wire wire_5586;
    wire wire_5587;
    wire wire_5588;
    wire wire_5589;
    wire wire_5590;
    wire wire_5617;
    wire wire_5620;
    wire wire_5623;
    wire wire_5626;
    wire wire_5629;
    wire wire_5632;
    wire wire_5635;
    wire wire_5638;
    wire wire_5665;
    wire wire_5668;
    wire wire_5671;
    wire wire_5674;
    wire wire_5677;
    wire wire_5680;
    wire wire_5683;
    wire wire_5686;
    wire wire_5713;
    wire wire_5716;
    wire wire_5719;
    wire wire_5722;
    wire wire_5725;
    wire wire_5728;
    wire wire_5731;
    wire wire_5734;
    wire wire_5761;
    wire wire_5764;
    wire wire_5767;
    wire wire_5770;
    wire wire_5773;
    wire wire_5776;
    wire wire_5779;
    wire wire_5782;
    wire wire_5809;
    wire wire_5812;
    wire wire_5815;
    wire wire_5818;
    wire wire_5821;
    wire wire_5824;
    wire wire_5827;
    wire wire_5830;
    wire wire_5857;
    wire wire_5860;
    wire wire_5863;
    wire wire_5866;
    wire wire_5869;
    wire wire_5872;
    wire wire_5875;
    wire wire_5878;
    wire wire_5905;
    wire wire_5908;
    wire wire_5911;
    wire wire_5914;
    wire wire_5917;
    wire wire_5920;
    wire wire_5923;
    wire wire_5926;
    wire wire_5953;
    wire wire_5956;
    wire wire_5959;
    wire wire_5962;
    wire wire_5965;
    wire wire_5968;
    wire wire_5971;
    wire wire_5974;
    wire wire_6001;
    wire wire_6004;
    wire wire_6007;
    wire wire_6010;
    wire wire_6013;
    wire wire_6016;
    wire wire_6019;
    wire wire_6022;
    wire wire_6049;
    wire wire_6052;
    wire wire_6055;
    wire wire_6058;
    wire wire_6061;
    wire wire_6064;
    wire wire_6067;
    wire wire_6070;
    wire wire_6097;
    wire wire_6100;
    wire wire_6103;
    wire wire_6106;
    wire wire_6109;
    wire wire_6112;
    wire wire_6115;
    wire wire_6118;
    wire wire_6120;
    wire wire_6121;
    wire wire_6122;
    wire wire_6123;
    wire wire_6124;
    wire wire_6125;
    wire wire_6126;
    wire wire_6127;
    wire wire_6128;
    wire wire_6129;
    wire wire_6130;
    wire wire_6131;
    wire wire_6132;
    wire wire_6133;
    wire wire_6134;
    wire wire_6135;
    wire wire_6136;
    wire wire_6137;
    wire wire_6138;
    wire wire_6139;
    wire wire_6140;
    wire wire_6141;
    wire wire_6142;
    wire wire_6143;
    wire wire_6144;
    wire wire_6145;
    wire wire_6146;
    wire wire_6147;
    wire wire_6148;
    wire wire_6149;
    wire wire_6150;
    wire wire_6151;
    wire wire_6152;
    wire wire_6153;
    wire wire_6154;
    wire wire_6155;
    wire wire_6156;
    wire wire_6157;
    wire wire_6158;
    wire wire_6159;
    wire wire_6160;
    wire wire_6161;
    wire wire_6162;
    wire wire_6163;
    wire wire_6164;
    wire wire_6165;
    wire wire_6166;
    wire wire_6167;
    wire wire_6168;
    wire wire_6169;
    wire wire_6170;
    wire wire_6171;
    wire wire_6172;
    wire wire_6173;
    wire wire_6174;
    wire wire_6175;
    wire wire_6176;
    wire wire_6177;
    wire wire_6178;
    wire wire_6179;
    wire wire_6180;
    wire wire_6181;
    wire wire_6182;
    wire wire_6183;
    wire wire_6184;
    wire wire_6185;
    wire wire_6186;
    wire wire_6187;
    wire wire_6188;
    wire wire_6189;
    wire wire_6190;
    wire wire_6191;
    wire wire_6192;
    wire wire_6193;
    wire wire_6194;
    wire wire_6195;
    wire wire_6196;
    wire wire_6197;
    wire wire_6198;
    wire wire_6199;
    wire wire_6200;
    wire wire_6201;
    wire wire_6202;
    wire wire_6203;
    wire wire_6204;
    wire wire_6205;
    wire wire_6206;
    wire wire_6207;
    wire wire_6208;
    wire wire_6209;
    wire wire_6210;
    wire wire_6211;
    wire wire_6212;
    wire wire_6213;
    wire wire_6214;
    wire wire_6215;
    wire wire_6216;
    wire wire_6217;
    wire wire_6218;
    wire wire_6219;
    wire wire_6220;
    wire wire_6221;
    wire wire_6222;
    wire wire_6223;
    wire wire_6224;
    wire wire_6225;
    wire wire_6226;
    wire wire_6227;
    wire wire_6228;
    wire wire_6229;
    wire wire_6230;
    wire wire_6231;
    wire wire_6232;
    wire wire_6233;
    wire wire_6234;
    wire wire_6235;
    wire wire_6236;
    wire wire_6237;
    wire wire_6238;
    wire wire_6239;
    wire wire_6240;
    wire wire_6241;
    wire wire_6242;
    wire wire_6243;
    wire wire_6244;
    wire wire_6245;
    wire wire_6246;
    wire wire_6247;
    wire wire_6248;
    wire wire_6249;
    wire wire_6250;
    wire wire_6251;
    wire wire_6252;
    wire wire_6253;
    wire wire_6254;
    wire wire_6255;
    wire wire_6256;
    wire wire_6257;
    wire wire_6258;
    wire wire_6259;
    wire wire_6260;
    wire wire_6261;
    wire wire_6262;
    wire wire_6263;
    wire wire_6264;
    wire wire_6265;
    wire wire_6266;
    wire wire_6267;
    wire wire_6268;
    wire wire_6269;
    wire wire_6270;
    wire wire_6271;
    wire wire_6272;
    wire wire_6273;
    wire wire_6274;
    wire wire_6275;
    wire wire_6276;
    wire wire_6277;
    wire wire_6278;
    wire wire_6279;
    wire wire_6280;
    wire wire_6281;
    wire wire_6282;
    wire wire_6283;
    wire wire_6284;
    wire wire_6285;
    wire wire_6286;
    wire wire_6287;
    wire wire_6288;
    wire wire_6289;
    wire wire_6290;
    wire wire_6291;
    wire wire_6292;
    wire wire_6293;
    wire wire_6294;
    wire wire_6295;
    wire wire_6296;
    wire wire_6297;
    wire wire_6298;
    wire wire_6299;
    wire wire_6300;
    wire wire_6301;
    wire wire_6302;
    wire wire_6303;
    wire wire_6304;
    wire wire_6305;
    wire wire_6306;
    wire wire_6307;
    wire wire_6308;
    wire wire_6309;
    wire wire_6310;
    wire wire_6311;
    wire wire_6312;
    wire wire_6313;
    wire wire_6314;
    wire wire_6315;
    wire wire_6316;
    wire wire_6317;
    wire wire_6318;
    wire wire_6319;
    wire wire_6320;
    wire wire_6321;
    wire wire_6322;
    wire wire_6323;
    wire wire_6324;
    wire wire_6325;
    wire wire_6326;
    wire wire_6327;
    wire wire_6328;
    wire wire_6329;
    wire wire_6330;
    wire wire_6331;
    wire wire_6332;
    wire wire_6333;
    wire wire_6334;
    wire wire_6335;
    wire wire_6336;
    wire wire_6337;
    wire wire_6338;
    wire wire_6339;
    wire wire_6340;
    wire wire_6341;
    wire wire_6342;
    wire wire_6343;
    wire wire_6344;
    wire wire_6345;
    wire wire_6346;
    wire wire_6347;
    wire wire_6348;
    wire wire_6349;
    wire wire_6350;
    wire wire_6351;
    wire wire_6352;
    wire wire_6353;
    wire wire_6354;
    wire wire_6355;
    wire wire_6356;
    wire wire_6357;
    wire wire_6358;
    wire wire_6359;
    wire wire_6360;
    wire wire_6361;
    wire wire_6362;
    wire wire_6363;
    wire wire_6364;
    wire wire_6365;
    wire wire_6366;
    wire wire_6367;
    wire wire_6368;
    wire wire_6369;
    wire wire_6370;
    wire wire_6371;
    wire wire_6372;
    wire wire_6373;
    wire wire_6374;
    wire wire_6375;
    wire wire_6376;
    wire wire_6377;
    wire wire_6378;
    wire wire_6379;
    wire wire_6380;
    wire wire_6381;
    wire wire_6382;
    wire wire_6383;
    wire wire_6384;
    wire wire_6385;
    wire wire_6386;
    wire wire_6387;
    wire wire_6388;
    wire wire_6389;
    wire wire_6390;
    wire wire_6391;
    wire wire_6392;
    wire wire_6393;
    wire wire_6394;
    wire wire_6395;
    wire wire_6396;
    wire wire_6397;
    wire wire_6398;
    wire wire_6399;
    wire wire_6400;
    wire wire_6401;
    wire wire_6402;
    wire wire_6403;
    wire wire_6404;
    wire wire_6405;
    wire wire_6406;
    wire wire_6407;
    wire wire_6408;
    wire wire_6409;
    wire wire_6410;
    wire wire_6411;
    wire wire_6412;
    wire wire_6413;
    wire wire_6414;
    wire wire_6415;
    wire wire_6416;
    wire wire_6417;
    wire wire_6418;
    wire wire_6419;
    wire wire_6420;
    wire wire_6421;
    wire wire_6422;
    wire wire_6423;
    wire wire_6424;
    wire wire_6425;
    wire wire_6426;
    wire wire_6427;
    wire wire_6428;
    wire wire_6429;
    wire wire_6430;
    wire wire_6431;
    wire wire_6432;
    wire wire_6433;
    wire wire_6434;
    wire wire_6435;
    wire wire_6436;
    wire wire_6437;
    wire wire_6438;
    wire wire_6439;
    wire wire_6440;
    wire wire_6441;
    wire wire_6442;
    wire wire_6443;
    wire wire_6444;
    wire wire_6445;
    wire wire_6446;
    wire wire_6447;
    wire wire_6448;
    wire wire_6449;
    wire wire_6450;
    wire wire_6451;
    wire wire_6452;
    wire wire_6453;
    wire wire_6454;
    wire wire_6455;
    wire wire_6456;
    wire wire_6457;
    wire wire_6458;
    wire wire_6459;
    wire wire_6460;
    wire wire_6461;
    wire wire_6462;
    wire wire_6463;
    wire wire_6464;
    wire wire_6465;
    wire wire_6466;
    wire wire_6467;
    wire wire_6468;
    wire wire_6469;
    wire wire_6470;
    wire wire_6471;
    wire wire_6472;
    wire wire_6473;
    wire wire_6474;
    wire wire_6475;
    wire wire_6476;
    wire wire_6477;
    wire wire_6478;
    wire wire_6479;
    wire wire_6480;
    wire wire_6481;
    wire wire_6482;
    wire wire_6483;
    wire wire_6484;
    wire wire_6485;
    wire wire_6486;
    wire wire_6487;
    wire wire_6488;
    wire wire_6489;
    wire wire_6490;
    wire wire_6491;
    wire wire_6492;
    wire wire_6493;
    wire wire_6494;
    wire wire_6495;
    wire wire_6496;
    wire wire_6497;
    wire wire_6498;
    wire wire_6499;
    wire wire_6500;
    wire wire_6501;
    wire wire_6502;
    wire wire_6503;
    wire wire_6504;
    wire wire_6505;
    wire wire_6506;
    wire wire_6507;
    wire wire_6508;
    wire wire_6509;
    wire wire_6510;
    wire wire_6511;
    wire wire_6512;
    wire wire_6513;
    wire wire_6514;
    wire wire_6515;
    wire wire_6516;
    wire wire_6517;
    wire wire_6518;
    wire wire_6519;
    wire wire_6520;
    wire wire_6521;
    wire wire_6522;
    wire wire_6523;
    wire wire_6524;
    wire wire_6525;
    wire wire_6526;
    wire wire_6527;
    wire wire_6528;
    wire wire_6529;
    wire wire_6530;
    wire wire_6531;
    wire wire_6532;
    wire wire_6533;
    wire wire_6534;
    wire wire_6535;
    wire wire_6536;
    wire wire_6537;
    wire wire_6538;
    wire wire_6539;
    wire wire_6540;
    wire wire_6541;
    wire wire_6542;
    wire wire_6543;
    wire wire_6544;
    wire wire_6545;
    wire wire_6546;
    wire wire_6547;
    wire wire_6548;
    wire wire_6549;
    wire wire_6550;
    wire wire_6551;
    wire wire_6552;
    wire wire_6553;
    wire wire_6554;
    wire wire_6555;
    wire wire_6556;
    wire wire_6557;
    wire wire_6558;
    wire wire_6559;
    wire wire_6560;
    wire wire_6561;
    wire wire_6562;
    wire wire_6563;
    wire wire_6564;
    wire wire_6565;
    wire wire_6566;
    wire wire_6567;
    wire wire_6568;
    wire wire_6569;
    wire wire_6570;
    wire wire_6571;
    wire wire_6572;
    wire wire_6573;
    wire wire_6574;
    wire wire_6575;
    wire wire_6576;
    wire wire_6577;
    wire wire_6578;
    wire wire_6579;
    wire wire_6580;
    wire wire_6581;
    wire wire_6582;
    wire wire_6583;
    wire wire_6584;
    wire wire_6585;
    wire wire_6586;
    wire wire_6587;
    wire wire_6588;
    wire wire_6589;
    wire wire_6590;
    wire wire_6591;
    wire wire_6592;
    wire wire_6593;
    wire wire_6594;
    wire wire_6595;
    wire wire_6596;
    wire wire_6597;
    wire wire_6598;
    wire wire_6599;
    wire wire_6600;
    wire wire_6601;
    wire wire_6602;
    wire wire_6603;
    wire wire_6604;
    wire wire_6605;
    wire wire_6606;
    wire wire_6607;
    wire wire_6608;
    wire wire_6609;
    wire wire_6610;
    wire wire_6611;
    wire wire_6612;
    wire wire_6613;
    wire wire_6614;
    wire wire_6615;
    wire wire_6616;
    wire wire_6617;
    wire wire_6618;
    wire wire_6619;
    wire wire_6620;
    wire wire_6621;
    wire wire_6622;
    wire wire_6623;
    wire wire_6624;
    wire wire_6625;
    wire wire_6626;
    wire wire_6627;
    wire wire_6628;
    wire wire_6629;
    wire wire_6630;
    wire wire_6631;
    wire wire_6632;
    wire wire_6633;
    wire wire_6634;
    wire wire_6635;
    wire wire_6636;
    wire wire_6637;
    wire wire_6638;
    wire wire_6639;
    wire wire_6640;
    wire wire_6641;
    wire wire_6642;
    wire wire_6643;
    wire wire_6644;
    wire wire_6645;
    wire wire_6646;
    wire wire_6647;
    wire wire_6648;
    wire wire_6649;
    wire wire_6650;
    wire wire_6651;
    wire wire_6652;
    wire wire_6653;
    wire wire_6654;
    wire wire_6655;
    wire wire_6656;
    wire wire_6657;
    wire wire_6658;
    wire wire_6659;
    wire wire_6660;
    wire wire_6661;
    wire wire_6662;
    wire wire_6663;
    wire wire_6664;
    wire wire_6665;
    wire wire_6666;
    wire wire_6667;
    wire wire_6668;
    wire wire_6669;
    wire wire_6670;
    wire wire_6671;
    wire wire_6672;
    wire wire_6673;
    wire wire_6674;
    wire wire_6675;
    wire wire_6676;
    wire wire_6677;
    wire wire_6678;
    wire wire_6679;
    wire wire_6680;
    wire wire_6681;
    wire wire_6682;
    wire wire_6683;
    wire wire_6684;
    wire wire_6685;
    wire wire_6686;
    wire wire_6687;
    wire wire_6688;
    wire wire_6689;
    wire wire_6690;
    wire wire_6691;
    wire wire_6692;
    wire wire_6693;
    wire wire_6694;
    wire wire_6695;
    wire wire_6696;
    wire wire_6697;
    wire wire_6698;
    wire wire_6699;
    wire wire_6700;
    wire wire_6701;
    wire wire_6702;
    wire wire_6703;
    wire wire_6704;
    wire wire_6705;
    wire wire_6706;
    wire wire_6707;
    wire wire_6708;
    wire wire_6709;
    wire wire_6710;
    wire wire_6711;
    wire wire_6712;
    wire wire_6713;
    wire wire_6714;
    wire wire_6715;
    wire wire_6716;
    wire wire_6717;
    wire wire_6718;
    wire wire_6719;
    wire wire_6720;
    wire wire_6721;
    wire wire_6722;
    wire wire_6723;
    wire wire_6724;
    wire wire_6725;
    wire wire_6726;
    wire wire_6727;
    wire wire_6728;
    wire wire_6729;
    wire wire_6730;
    wire wire_6731;
    wire wire_6732;
    wire wire_6733;
    wire wire_6734;
    wire wire_6735;
    wire wire_6736;
    wire wire_6737;
    wire wire_6738;
    wire wire_6739;
    wire wire_6740;
    wire wire_6741;
    wire wire_6742;
    wire wire_6743;
    wire wire_6744;
    wire wire_6745;
    wire wire_6746;
    wire wire_6747;
    wire wire_6748;
    wire wire_6749;
    wire wire_6750;
    wire wire_6751;
    wire wire_6752;
    wire wire_6753;
    wire wire_6754;
    wire wire_6755;
    wire wire_6756;
    wire wire_6757;
    wire wire_6758;
    wire wire_6759;
    wire wire_6760;
    wire wire_6761;
    wire wire_6762;
    wire wire_6763;
    wire wire_6764;
    wire wire_6765;
    wire wire_6766;
    wire wire_6767;
    wire wire_6768;
    wire wire_6769;
    wire wire_6770;
    wire wire_6771;
    wire wire_6772;
    wire wire_6773;
    wire wire_6774;
    wire wire_6775;
    wire wire_6776;
    wire wire_6777;
    wire wire_6778;
    wire wire_6779;
    wire wire_6780;
    wire wire_6781;
    wire wire_6782;
    wire wire_6783;
    wire wire_6784;
    wire wire_6785;
    wire wire_6786;
    wire wire_6787;
    wire wire_6788;
    wire wire_6789;
    wire wire_6790;
    wire wire_6791;
    wire wire_6792;
    wire wire_6793;
    wire wire_6794;
    wire wire_6795;
    wire wire_6796;
    wire wire_6797;
    wire wire_6798;
    wire wire_6799;
    wire wire_6800;
    wire wire_6801;
    wire wire_6802;
    wire wire_6803;
    wire wire_6804;
    wire wire_6805;
    wire wire_6806;
    wire wire_6807;
    wire wire_6808;
    wire wire_6809;
    wire wire_6810;
    wire wire_6811;
    wire wire_6812;
    wire wire_6813;
    wire wire_6814;
    wire wire_6815;
    wire wire_6816;
    wire wire_6817;
    wire wire_6818;
    wire wire_6819;
    wire wire_6820;
    wire wire_6821;
    wire wire_6822;
    wire wire_6823;
    wire wire_6824;
    wire wire_6825;
    wire wire_6826;
    wire wire_6827;
    wire wire_6828;
    wire wire_6829;
    wire wire_6830;
    wire wire_6831;
    wire wire_6832;
    wire wire_6833;
    wire wire_6834;
    wire wire_6835;
    wire wire_6836;
    wire wire_6837;
    wire wire_6838;
    wire wire_6839;
    wire wire_6840;
    wire wire_6841;
    wire wire_6842;
    wire wire_6843;
    wire wire_6844;
    wire wire_6845;
    wire wire_6846;
    wire wire_6847;
    wire wire_6848;
    wire wire_6849;
    wire wire_6850;
    wire wire_6851;
    wire wire_6852;
    wire wire_6853;
    wire wire_6854;
    wire wire_6855;
    wire wire_6856;
    wire wire_6857;
    wire wire_6858;
    wire wire_6859;
    wire wire_6860;
    wire wire_6861;
    wire wire_6862;
    wire wire_6863;
    wire wire_6864;
    wire wire_6865;
    wire wire_6866;
    wire wire_6867;
    wire wire_6868;
    wire wire_6869;
    wire wire_6870;
    wire wire_6871;
    wire wire_6872;
    wire wire_6873;
    wire wire_6874;
    wire wire_6875;
    wire wire_6876;
    wire wire_6877;
    wire wire_6878;
    wire wire_6879;
    wire wire_6880;
    wire wire_6881;
    wire wire_6882;
    wire wire_6883;
    wire wire_6884;
    wire wire_6885;
    wire wire_6886;
    wire wire_6887;
    wire wire_6888;
    wire wire_6889;
    wire wire_6890;
    wire wire_6891;
    wire wire_6892;
    wire wire_6893;
    wire wire_6894;
    wire wire_6895;
    wire wire_6896;
    wire wire_6897;
    wire wire_6898;
    wire wire_6899;
    wire wire_6900;
    wire wire_6901;
    wire wire_6902;
    wire wire_6903;
    wire wire_6904;
    wire wire_6905;
    wire wire_6906;
    wire wire_6907;
    wire wire_6908;
    wire wire_6909;
    wire wire_6910;
    wire wire_6911;
    wire wire_6912;
    wire wire_6913;
    wire wire_6914;
    wire wire_6915;
    wire wire_6916;
    wire wire_6917;
    wire wire_6918;
    wire wire_6919;
    wire wire_6920;
    wire wire_6921;
    wire wire_6922;
    wire wire_6923;
    wire wire_6924;
    wire wire_6925;
    wire wire_6926;
    wire wire_6927;
    wire wire_6928;
    wire wire_6929;
    wire wire_6930;
    wire wire_6931;
    wire wire_6932;
    wire wire_6933;
    wire wire_6934;
    wire wire_6935;
    wire wire_6936;
    wire wire_6937;
    wire wire_6938;
    wire wire_6939;
    wire wire_6940;
    wire wire_6941;
    wire wire_6942;
    wire wire_6943;
    wire wire_6944;
    wire wire_6945;
    wire wire_6946;
    wire wire_6947;
    wire wire_6948;
    wire wire_6949;
    wire wire_6950;
    wire wire_6951;
    wire wire_6952;
    wire wire_6953;
    wire wire_6954;
    wire wire_6955;
    wire wire_6956;
    wire wire_6957;
    wire wire_6958;
    wire wire_6959;
    wire wire_6960;
    wire wire_6961;
    wire wire_6962;
    wire wire_6963;
    wire wire_6964;
    wire wire_6965;
    wire wire_6966;
    wire wire_6967;
    wire wire_6968;
    wire wire_6969;
    wire wire_6970;
    wire wire_6971;
    wire wire_6972;
    wire wire_6973;
    wire wire_6974;
    wire wire_6975;
    wire wire_6976;
    wire wire_6977;
    wire wire_6978;
    wire wire_6979;
    wire wire_6980;
    wire wire_6981;
    wire wire_6982;
    wire wire_6983;
    wire wire_6984;
    wire wire_6985;
    wire wire_6986;
    wire wire_6987;
    wire wire_6988;
    wire wire_6989;
    wire wire_6990;
    wire wire_6991;
    wire wire_6992;
    wire wire_6993;
    wire wire_6994;
    wire wire_6995;
    wire wire_6996;
    wire wire_6997;
    wire wire_6998;
    wire wire_6999;
    wire wire_7000;
    wire wire_7001;
    wire wire_7002;
    wire wire_7003;
    wire wire_7004;
    wire wire_7005;
    wire wire_7006;
    wire wire_7007;
    wire wire_7008;
    wire wire_7009;
    wire wire_7010;
    wire wire_7011;
    wire wire_7012;
    wire wire_7013;
    wire wire_7014;
    wire wire_7015;
    wire wire_7016;
    wire wire_7017;
    wire wire_7018;
    wire wire_7019;
    wire wire_7020;
    wire wire_7021;
    wire wire_7022;
    wire wire_7023;
    wire wire_7024;
    wire wire_7025;
    wire wire_7026;
    wire wire_7027;
    wire wire_7028;
    wire wire_7029;
    wire wire_7030;
    wire wire_7031;
    wire wire_7032;
    wire wire_7033;
    wire wire_7034;
    wire wire_7035;
    wire wire_7036;
    wire wire_7037;
    wire wire_7038;
    wire wire_7039;
    wire wire_7040;
    wire wire_7041;
    wire wire_7042;
    wire wire_7043;
    wire wire_7044;
    wire wire_7045;
    wire wire_7046;
    wire wire_7047;
    wire wire_7048;
    wire wire_7049;
    wire wire_7050;
    wire wire_7051;
    wire wire_7052;
    wire wire_7053;
    wire wire_7054;
    wire wire_7055;
    wire wire_7056;
    wire wire_7057;
    wire wire_7058;
    wire wire_7059;
    wire wire_7060;
    wire wire_7061;
    wire wire_7062;
    wire wire_7063;
    wire wire_7064;
    wire wire_7065;
    wire wire_7066;
    wire wire_7067;
    wire wire_7068;
    wire wire_7069;
    wire wire_7070;
    wire wire_7071;
    wire wire_7072;
    wire wire_7073;
    wire wire_7074;
    wire wire_7075;
    wire wire_7076;
    wire wire_7077;
    wire wire_7078;
    wire wire_7079;
    wire wire_7080;
    wire wire_7081;
    wire wire_7082;
    wire wire_7083;
    wire wire_7084;
    wire wire_7085;
    wire wire_7086;
    wire wire_7087;
    wire wire_7088;
    wire wire_7089;
    wire wire_7090;
    wire wire_7091;
    wire wire_7092;
    wire wire_7093;
    wire wire_7094;
    wire wire_7095;
    wire wire_7096;
    wire wire_7097;
    wire wire_7098;
    wire wire_7099;
    wire wire_7100;
    wire wire_7101;
    wire wire_7102;
    wire wire_7103;
    wire wire_7104;
    wire wire_7105;
    wire wire_7106;
    wire wire_7107;
    wire wire_7108;
    wire wire_7109;
    wire wire_7110;
    wire wire_7111;
    wire wire_7112;
    wire wire_7113;
    wire wire_7114;
    wire wire_7115;
    wire wire_7116;
    wire wire_7117;
    wire wire_7118;
    wire wire_7119;
    wire wire_7120;
    wire wire_7121;
    wire wire_7122;
    wire wire_7123;
    wire wire_7124;
    wire wire_7125;
    wire wire_7126;
    wire wire_7127;
    wire wire_7128;
    wire wire_7129;
    wire wire_7130;
    wire wire_7131;
    wire wire_7132;
    wire wire_7133;
    wire wire_7134;
    wire wire_7135;
    wire wire_7136;
    wire wire_7137;
    wire wire_7138;
    wire wire_7139;
    wire wire_7140;
    wire wire_7141;
    wire wire_7142;
    wire wire_7143;
    wire wire_7144;
    wire wire_7145;
    wire wire_7146;
    wire wire_7147;
    wire wire_7148;
    wire wire_7149;
    wire wire_7150;
    wire wire_7151;
    wire wire_7152;
    wire wire_7153;
    wire wire_7154;
    wire wire_7155;
    wire wire_7156;
    wire wire_7157;
    wire wire_7158;
    wire wire_7159;
    wire wire_7160;
    wire wire_7161;
    wire wire_7162;
    wire wire_7163;
    wire wire_7164;
    wire wire_7165;
    wire wire_7166;
    wire wire_7167;
    wire wire_7168;
    wire wire_7169;
    wire wire_7170;
    wire wire_7171;
    wire wire_7172;
    wire wire_7173;
    wire wire_7174;
    wire wire_7175;
    wire wire_7176;
    wire wire_7177;
    wire wire_7178;
    wire wire_7179;
    wire wire_7180;
    wire wire_7181;
    wire wire_7182;
    wire wire_7183;
    wire wire_7184;
    wire wire_7185;
    wire wire_7186;
    wire wire_7187;
    wire wire_7188;
    wire wire_7189;
    wire wire_7190;
    wire wire_7191;
    wire wire_7192;
    wire wire_7193;
    wire wire_7194;
    wire wire_7195;
    wire wire_7196;
    wire wire_7197;
    wire wire_7198;
    wire wire_7199;
    wire wire_7200;
    wire wire_7201;
    wire wire_7202;
    wire wire_7203;
    wire wire_7204;
    wire wire_7205;
    wire wire_7206;
    wire wire_7207;
    wire wire_7208;
    wire wire_7209;
    wire wire_7210;
    wire wire_7211;
    wire wire_7212;
    wire wire_7213;
    wire wire_7214;
    wire wire_7215;
    wire wire_7216;
    wire wire_7217;
    wire wire_7218;
    wire wire_7219;
    wire wire_7220;
    wire wire_7221;
    wire wire_7222;
    wire wire_7223;
    wire wire_7224;
    wire wire_7225;
    wire wire_7226;
    wire wire_7227;
    wire wire_7228;
    wire wire_7229;
    wire wire_7230;
    wire wire_7231;
    wire wire_7232;
    wire wire_7233;
    wire wire_7234;
    wire wire_7235;
    wire wire_7236;
    wire wire_7237;
    wire wire_7238;
    wire wire_7239;
    wire wire_7240;
    wire wire_7241;
    wire wire_7242;
    wire wire_7243;
    wire wire_7244;
    wire wire_7245;
    wire wire_7246;
    wire wire_7247;
    wire wire_7248;
    wire wire_7249;
    wire wire_7250;
    wire wire_7251;
    wire wire_7252;
    wire wire_7253;
    wire wire_7254;
    wire wire_7255;
    wire wire_7256;
    wire wire_7257;
    wire wire_7258;
    wire wire_7259;
    wire wire_7260;
    wire wire_7261;
    wire wire_7262;
    wire wire_7263;
    wire wire_7264;
    wire wire_7265;
    wire wire_7266;
    wire wire_7267;
    wire wire_7268;
    wire wire_7269;
    wire wire_7270;
    wire wire_7271;
    wire wire_7272;
    wire wire_7273;
    wire wire_7274;
    wire wire_7275;
    wire wire_7276;
    wire wire_7277;
    wire wire_7278;
    wire wire_7279;
    wire wire_7280;
    wire wire_7281;
    wire wire_7282;
    wire wire_7283;
    wire wire_7284;
    wire wire_7285;
    wire wire_7286;
    wire wire_7287;
    wire wire_7288;
    wire wire_7289;
    wire wire_7290;
    wire wire_7291;
    wire wire_7292;
    wire wire_7293;
    wire wire_7294;
    wire wire_7295;
    wire wire_7296;
    wire wire_7297;
    wire wire_7298;
    wire wire_7299;
    wire wire_7300;
    wire wire_7301;
    wire wire_7302;
    wire wire_7303;
    wire wire_7304;
    wire wire_7305;
    wire wire_7306;
    wire wire_7307;
    wire wire_7308;
    wire wire_7309;
    wire wire_7310;
    wire wire_7311;
    wire wire_7312;
    wire wire_7313;
    wire wire_7314;
    wire wire_7315;
    wire wire_7316;
    wire wire_7317;
    wire wire_7318;
    wire wire_7319;
    wire wire_7320;
    wire wire_7321;
    wire wire_7322;
    wire wire_7323;
    wire wire_7324;
    wire wire_7325;
    wire wire_7326;
    wire wire_7327;
    wire wire_7328;
    wire wire_7329;
    wire wire_7330;
    wire wire_7331;
    wire wire_7332;
    wire wire_7333;
    wire wire_7334;
    wire wire_7335;
    wire wire_7336;
    wire wire_7337;
    wire wire_7338;
    wire wire_7339;
    wire wire_7340;
    wire wire_7341;
    wire wire_7342;
    wire wire_7343;
    wire wire_7344;
    wire wire_7345;
    wire wire_7346;
    wire wire_7347;
    wire wire_7348;
    wire wire_7349;
    wire wire_7350;
    wire wire_7351;
    wire wire_7352;
    wire wire_7353;
    wire wire_7354;
    wire wire_7355;
    wire wire_7356;
    wire wire_7357;
    wire wire_7358;
    wire wire_7359;
    wire wire_7360;
    wire wire_7361;
    wire wire_7362;
    wire wire_7363;
    wire wire_7364;
    wire wire_7365;
    wire wire_7366;
    wire wire_7367;
    wire wire_7368;
    wire wire_7369;
    wire wire_7370;
    wire wire_7371;
    wire wire_7372;
    wire wire_7373;
    wire wire_7374;
    wire wire_7375;
    wire wire_7376;
    wire wire_7377;
    wire wire_7378;
    wire wire_7379;
    wire wire_7380;
    wire wire_7381;
    wire wire_7382;
    wire wire_7383;
    wire wire_7384;
    wire wire_7385;
    wire wire_7386;
    wire wire_7387;
    wire wire_7388;
    wire wire_7389;
    wire wire_7390;
    wire wire_7391;
    wire wire_7392;
    wire wire_7393;
    wire wire_7394;
    wire wire_7395;
    wire wire_7396;
    wire wire_7397;
    wire wire_7398;
    wire wire_7399;
    wire wire_7400;
    wire wire_7401;
    wire wire_7402;
    wire wire_7403;
    wire wire_7404;
    wire wire_7405;
    wire wire_7406;
    wire wire_7407;
    wire wire_7408;
    wire wire_7409;
    wire wire_7410;
    wire wire_7411;
    wire wire_7412;
    wire wire_7413;
    wire wire_7414;
    wire wire_7415;
    wire wire_7416;
    wire wire_7417;
    wire wire_7418;
    wire wire_7419;
    wire wire_7420;
    wire wire_7421;
    wire wire_7422;
    wire wire_7423;
    wire wire_7424;
    wire wire_7425;
    wire wire_7426;
    wire wire_7427;
    wire wire_7428;
    wire wire_7429;
    wire wire_7430;
    wire wire_7431;
    wire wire_7432;
    wire wire_7433;
    wire wire_7434;
    wire wire_7435;
    wire wire_7436;
    wire wire_7437;
    wire wire_7438;
    wire wire_7439;
    wire wire_7440;
    wire wire_7441;
    wire wire_7442;
    wire wire_7443;
    wire wire_7444;
    wire wire_7445;
    wire wire_7446;
    wire wire_7447;
    wire wire_7448;
    wire wire_7449;
    wire wire_7450;
    wire wire_7451;
    wire wire_7452;
    wire wire_7453;
    wire wire_7454;
    wire wire_7455;
    wire wire_7456;
    wire wire_7457;
    wire wire_7458;
    wire wire_7459;
    wire wire_7460;
    wire wire_7461;
    wire wire_7462;
    wire wire_7463;
    wire wire_7464;
    wire wire_7465;
    wire wire_7466;
    wire wire_7467;
    wire wire_7468;
    wire wire_7469;
    wire wire_7470;
    wire wire_7471;
    wire wire_7472;
    wire wire_7473;
    wire wire_7474;
    wire wire_7475;
    wire wire_7476;
    wire wire_7477;
    wire wire_7478;
    wire wire_7479;
    wire wire_7480;
    wire wire_7481;
    wire wire_7482;
    wire wire_7483;
    wire wire_7484;
    wire wire_7485;
    wire wire_7486;
    wire wire_7487;
    wire wire_7488;
    wire wire_7489;
    wire wire_7490;
    wire wire_7491;
    wire wire_7492;
    wire wire_7493;
    wire wire_7494;
    wire wire_7495;
    wire wire_7496;
    wire wire_7497;
    wire wire_7498;
    wire wire_7499;
    wire wire_7500;
    wire wire_7501;
    wire wire_7502;
    wire wire_7503;
    wire wire_7504;
    wire wire_7505;
    wire wire_7506;
    wire wire_7507;
    wire wire_7508;
    wire wire_7509;
    wire wire_7510;
    wire wire_7511;
    wire wire_7512;
    wire wire_7513;
    wire wire_7514;
    wire wire_7515;
    wire wire_7516;
    wire wire_7517;
    wire wire_7518;
    wire wire_7519;
    wire wire_7520;
    wire wire_7521;
    wire wire_7522;
    wire wire_7523;
    wire wire_7524;
    wire wire_7525;
    wire wire_7526;
    wire wire_7527;
    wire wire_7528;
    wire wire_7529;
    wire wire_7530;
    wire wire_7531;
    wire wire_7532;
    wire wire_7533;
    wire wire_7534;
    wire wire_7535;
    wire wire_7536;
    wire wire_7537;
    wire wire_7538;
    wire wire_7539;
    wire wire_7540;
    wire wire_7541;
    wire wire_7542;
    wire wire_7543;
    wire wire_7544;
    wire wire_7545;
    wire wire_7546;
    wire wire_7547;
    wire wire_7548;
    wire wire_7549;
    wire wire_7550;
    wire wire_7551;
    wire wire_7552;
    wire wire_7553;
    wire wire_7554;
    wire wire_7555;
    wire wire_7556;
    wire wire_7557;
    wire wire_7558;
    wire wire_7559;
    wire wire_7560;
    wire wire_7561;
    wire wire_7562;
    wire wire_7563;
    wire wire_7564;
    wire wire_7565;
    wire wire_7566;
    wire wire_7567;
    wire wire_7568;
    wire wire_7569;
    wire wire_7570;
    wire wire_7571;
    wire wire_7572;
    wire wire_7573;
    wire wire_7574;
    wire wire_7575;
    wire wire_7576;
    wire wire_7577;
    wire wire_7578;
    wire wire_7579;
    wire wire_7580;
    wire wire_7581;
    wire wire_7582;
    wire wire_7583;
    wire wire_7584;
    wire wire_7585;
    wire wire_7586;
    wire wire_7587;
    wire wire_7588;
    wire wire_7589;
    wire wire_7590;
    wire wire_7591;
    wire wire_7592;
    wire wire_7593;
    wire wire_7594;
    wire wire_7595;
    wire wire_7596;
    wire wire_7597;
    wire wire_7598;
    wire wire_7599;
    wire wire_7600;
    wire wire_7601;
    wire wire_7602;
    wire wire_7603;
    wire wire_7604;
    wire wire_7605;
    wire wire_7606;
    wire wire_7607;
    wire wire_7608;
    wire wire_7609;
    wire wire_7610;
    wire wire_7611;
    wire wire_7612;
    wire wire_7613;
    wire wire_7614;
    wire wire_7615;
    wire wire_7616;
    wire wire_7617;
    wire wire_7618;
    wire wire_7619;
    wire wire_7620;
    wire wire_7621;
    wire wire_7622;
    wire wire_7623;
    wire wire_7624;
    wire wire_7625;
    wire wire_7626;
    wire wire_7627;
    wire wire_7628;
    wire wire_7629;
    wire wire_7630;
    wire wire_7631;
    wire wire_7632;
    wire wire_7633;
    wire wire_7634;
    wire wire_7635;
    wire wire_7636;
    wire wire_7637;
    wire wire_7638;
    wire wire_7639;
    wire wire_7640;
    wire wire_7641;
    wire wire_7642;
    wire wire_7643;
    wire wire_7644;
    wire wire_7645;
    wire wire_7646;
    wire wire_7647;
    wire wire_7648;
    wire wire_7649;
    wire wire_7650;
    wire wire_7651;
    wire wire_7652;
    wire wire_7653;
    wire wire_7654;
    wire wire_7655;
    wire wire_7656;
    wire wire_7657;
    wire wire_7658;
    wire wire_7659;
    wire wire_7660;
    wire wire_7661;
    wire wire_7662;
    wire wire_7663;
    wire wire_7664;
    wire wire_7665;
    wire wire_7666;
    wire wire_7667;
    wire wire_7668;
    wire wire_7669;
    wire wire_7670;
    wire wire_7671;
    wire wire_7672;
    wire wire_7673;
    wire wire_7674;
    wire wire_7675;
    wire wire_7676;
    wire wire_7677;
    wire wire_7678;
    wire wire_7679;
    wire wire_7680;
    wire wire_7681;
    wire wire_7682;
    wire wire_7683;
    wire wire_7684;
    wire wire_7685;
    wire wire_7686;
    wire wire_7687;
    wire wire_7688;
    wire wire_7689;
    wire wire_7690;
    wire wire_7691;
    wire wire_7692;
    wire wire_7693;
    wire wire_7694;
    wire wire_7695;
    wire wire_7696;
    wire wire_7697;
    wire wire_7698;
    wire wire_7699;
    wire wire_7700;
    wire wire_7701;
    wire wire_7702;
    wire wire_7703;
    wire wire_7704;
    wire wire_7705;
    wire wire_7706;
    wire wire_7707;
    wire wire_7708;
    wire wire_7709;
    wire wire_7710;
    wire wire_7711;
    wire wire_7712;
    wire wire_7713;
    wire wire_7714;
    wire wire_7715;
    wire wire_7716;
    wire wire_7717;
    wire wire_7718;
    wire wire_7719;
    wire wire_7720;
    wire wire_7721;
    wire wire_7722;
    wire wire_7723;
    wire wire_7724;
    wire wire_7725;
    wire wire_7726;
    wire wire_7727;
    wire wire_7728;
    wire wire_7729;
    wire wire_7730;
    wire wire_7731;
    wire wire_7732;
    wire wire_7733;
    wire wire_7734;
    wire wire_7735;
    wire wire_7736;
    wire wire_7737;
    wire wire_7738;
    wire wire_7739;
    wire wire_7740;
    wire wire_7741;
    wire wire_7742;
    wire wire_7743;
    wire wire_7744;
    wire wire_7745;
    wire wire_7746;
    wire wire_7747;
    wire wire_7748;
    wire wire_7749;
    wire wire_7750;
    wire wire_7751;
    wire wire_7752;
    wire wire_7753;
    wire wire_7754;
    wire wire_7755;
    wire wire_7756;
    wire wire_7757;
    wire wire_7758;
    wire wire_7759;
    wire wire_7760;
    wire wire_7761;
    wire wire_7762;
    wire wire_7763;
    wire wire_7764;
    wire wire_7765;
    wire wire_7766;
    wire wire_7767;
    wire wire_7768;
    wire wire_7769;
    wire wire_7770;
    wire wire_7771;
    wire wire_7772;
    wire wire_7773;
    wire wire_7774;
    wire wire_7775;
    wire wire_7776;
    wire wire_7777;
    wire wire_7778;
    wire wire_7779;
    wire wire_7780;
    wire wire_7781;
    wire wire_7782;
    wire wire_7783;
    wire wire_7784;
    wire wire_7785;
    wire wire_7786;
    wire wire_7787;
    wire wire_7788;
    wire wire_7789;
    wire wire_7790;
    wire wire_7791;
    wire wire_7792;
    wire wire_7793;
    wire wire_7794;
    wire wire_7795;
    wire wire_7796;
    wire wire_7797;
    wire wire_7798;
    wire wire_7799;
    wire wire_7800;
    wire wire_7801;
    wire wire_7802;
    wire wire_7803;
    wire wire_7804;
    wire wire_7805;
    wire wire_7806;
    wire wire_7807;
    wire wire_7808;
    wire wire_7809;
    wire wire_7810;
    wire wire_7811;
    wire wire_7812;
    wire wire_7813;
    wire wire_7814;
    wire wire_7815;
    wire wire_7816;
    wire wire_7817;
    wire wire_7818;
    wire wire_7819;
    wire wire_7820;
    wire wire_7821;
    wire wire_7822;
    wire wire_7823;
    wire wire_7824;
    wire wire_7825;
    wire wire_7826;
    wire wire_7827;
    wire wire_7828;
    wire wire_7829;
    wire wire_7830;
    wire wire_7831;
    wire wire_7832;
    wire wire_7833;
    wire wire_7834;
    wire wire_7835;
    wire wire_7836;
    wire wire_7837;
    wire wire_7838;
    wire wire_7839;
    wire wire_7840;
    wire wire_7841;
    wire wire_7842;
    wire wire_7843;
    wire wire_7844;
    wire wire_7845;
    wire wire_7846;
    wire wire_7847;
    wire wire_7848;
    wire wire_7849;
    wire wire_7850;
    wire wire_7851;
    wire wire_7852;
    wire wire_7853;
    wire wire_7854;
    wire wire_7855;
    wire wire_7856;
    wire wire_7857;
    wire wire_7858;
    wire wire_7859;
    wire wire_7860;
    wire wire_7861;
    wire wire_7862;
    wire wire_7863;
    wire wire_7864;
    wire wire_7865;
    wire wire_7866;
    wire wire_7867;
    wire wire_7868;
    wire wire_7869;
    wire wire_7870;
    wire wire_7871;
    wire wire_7872;
    wire wire_7873;
    wire wire_7874;
    wire wire_7875;
    wire wire_7876;
    wire wire_7877;
    wire wire_7878;
    wire wire_7879;
    wire wire_7880;
    wire wire_7881;
    wire wire_7882;
    wire wire_7883;
    wire wire_7884;
    wire wire_7885;
    wire wire_7886;
    wire wire_7887;
    wire wire_7888;
    wire wire_7889;
    wire wire_7890;
    wire wire_7891;
    wire wire_7892;
    wire wire_7893;
    wire wire_7894;
    wire wire_7895;
    wire wire_7896;
    wire wire_7897;
    wire wire_7898;
    wire wire_7899;
    wire wire_7900;
    wire wire_7901;
    wire wire_7902;
    wire wire_7903;
    wire wire_7904;
    wire wire_7905;
    wire wire_7906;
    wire wire_7907;
    wire wire_7908;
    wire wire_7909;
    wire wire_7910;
    wire wire_7911;
    wire wire_7912;
    wire wire_7913;
    wire wire_7914;
    wire wire_7915;
    wire wire_7916;
    wire wire_7917;
    wire wire_7918;
    wire wire_7919;
    wire wire_7920;
    wire wire_7921;
    wire wire_7922;
    wire wire_7923;
    wire wire_7924;
    wire wire_7925;
    wire wire_7926;
    wire wire_7927;
    wire wire_7928;
    wire wire_7929;
    wire wire_7930;
    wire wire_7931;
    wire wire_7932;
    wire wire_7933;
    wire wire_7934;
    wire wire_7935;
    wire wire_7936;
    wire wire_7937;
    wire wire_7938;
    wire wire_7939;
    wire wire_7940;
    wire wire_7941;
    wire wire_7942;
    wire wire_7943;
    wire wire_7944;
    wire wire_7945;
    wire wire_7946;
    wire wire_7947;
    wire wire_7948;
    wire wire_7949;
    wire wire_7950;
    wire wire_7951;
    wire wire_7952;
    wire wire_7953;
    wire wire_7954;
    wire wire_7955;
    wire wire_7956;
    wire wire_7957;
    wire wire_7958;
    wire wire_7959;
    wire wire_7960;
    wire wire_7961;
    wire wire_7962;
    wire wire_7963;
    wire wire_7964;
    wire wire_7965;
    wire wire_7966;
    wire wire_7967;
    wire wire_7968;
    wire wire_7969;
    wire wire_7970;
    wire wire_7971;
    wire wire_7972;
    wire wire_7973;
    wire wire_7974;
    wire wire_7975;
    wire wire_7976;
    wire wire_7977;
    wire wire_7978;
    wire wire_7979;
    wire wire_7980;
    wire wire_7981;
    wire wire_7982;
    wire wire_7983;
    wire wire_7984;
    wire wire_7985;
    wire wire_7986;
    wire wire_7987;
    wire wire_7988;
    wire wire_7989;
    wire wire_7990;
    wire wire_7991;
    wire wire_7992;
    wire wire_7993;
    wire wire_7994;
    wire wire_7995;
    wire wire_7996;
    wire wire_7997;
    wire wire_7998;
    wire wire_7999;
    wire wire_8000;
    wire wire_8001;
    wire wire_8002;
    wire wire_8003;
    wire wire_8004;
    wire wire_8005;
    wire wire_8006;
    wire wire_8007;
    wire wire_8008;
    wire wire_8009;
    wire wire_8010;
    wire wire_8011;
    wire wire_8012;
    wire wire_8013;
    wire wire_8014;
    wire wire_8015;
    wire wire_8016;
    wire wire_8017;
    wire wire_8018;
    wire wire_8019;
    wire wire_8020;
    wire wire_8021;
    wire wire_8022;
    wire wire_8023;
    wire wire_8024;
    wire wire_8025;
    wire wire_8026;
    wire wire_8027;
    wire wire_8028;
    wire wire_8029;
    wire wire_8030;
    wire wire_8031;
    wire wire_8032;
    wire wire_8033;
    wire wire_8034;
    wire wire_8035;
    wire wire_8036;
    wire wire_8037;
    wire wire_8038;
    wire wire_8039;
    wire wire_8040;
    wire wire_8041;
    wire wire_8042;
    wire wire_8043;
    wire wire_8044;
    wire wire_8045;
    wire wire_8046;
    wire wire_8047;
    wire wire_8048;
    wire wire_8049;
    wire wire_8050;
    wire wire_8051;
    wire wire_8052;
    wire wire_8053;
    wire wire_8054;
    wire wire_8055;
    wire wire_8056;
    wire wire_8057;
    wire wire_8058;
    wire wire_8059;
    wire wire_8060;
    wire wire_8061;
    wire wire_8062;
    wire wire_8063;
    wire wire_8064;
    wire wire_8065;
    wire wire_8066;
    wire wire_8067;
    wire wire_8068;
    wire wire_8069;
    wire wire_8070;
    wire wire_8071;
    wire wire_8072;
    wire wire_8073;
    wire wire_8074;
    wire wire_8075;
    wire wire_8076;
    wire wire_8077;
    wire wire_8078;
    wire wire_8079;
    wire wire_8080;
    wire wire_8081;
    wire wire_8082;
    wire wire_8083;
    wire wire_8084;
    wire wire_8085;
    wire wire_8086;
    wire wire_8087;
    wire wire_8088;
    wire wire_8089;
    wire wire_8090;
    wire wire_8091;
    wire wire_8092;
    wire wire_8093;
    wire wire_8094;
    wire wire_8095;
    wire wire_8096;
    wire wire_8097;
    wire wire_8098;
    wire wire_8099;
    wire wire_8100;
    wire wire_8101;
    wire wire_8102;
    wire wire_8103;
    wire wire_8104;
    wire wire_8105;
    wire wire_8106;
    wire wire_8107;
    wire wire_8108;
    wire wire_8109;
    wire wire_8110;
    wire wire_8111;
    wire wire_8112;
    wire wire_8113;
    wire wire_8114;
    wire wire_8115;
    wire wire_8116;
    wire wire_8117;
    wire wire_8118;
    wire wire_8119;
    wire wire_8120;
    wire wire_8121;
    wire wire_8122;
    wire wire_8123;
    wire wire_8124;
    wire wire_8125;
    wire wire_8126;
    wire wire_8127;
    wire wire_8128;
    wire wire_8129;
    wire wire_8130;
    wire wire_8131;
    wire wire_8132;
    wire wire_8133;
    wire wire_8134;
    wire wire_8135;
    wire wire_8136;
    wire wire_8137;
    wire wire_8138;
    wire wire_8139;
    wire wire_8140;
    wire wire_8141;
    wire wire_8142;
    wire wire_8143;
    wire wire_8144;
    wire wire_8145;
    wire wire_8146;
    wire wire_8147;
    wire wire_8148;
    wire wire_8149;
    wire wire_8150;
    wire wire_8151;
    wire wire_8152;
    wire wire_8153;
    wire wire_8154;
    wire wire_8155;
    wire wire_8156;
    wire wire_8157;
    wire wire_8158;
    wire wire_8159;
    wire wire_8160;
    wire wire_8161;
    wire wire_8162;
    wire wire_8163;
    wire wire_8164;
    wire wire_8165;
    wire wire_8166;
    wire wire_8167;
    wire wire_8168;
    wire wire_8169;
    wire wire_8170;
    wire wire_8171;
    wire wire_8172;
    wire wire_8173;
    wire wire_8174;
    wire wire_8175;
    wire wire_8176;
    wire wire_8177;
    wire wire_8178;
    wire wire_8179;
    wire wire_8180;
    wire wire_8181;
    wire wire_8182;
    wire wire_8183;
    wire wire_8184;
    wire wire_8185;
    wire wire_8186;
    wire wire_8187;
    wire wire_8188;
    wire wire_8189;
    wire wire_8190;
    wire wire_8191;
    wire wire_8192;
    wire wire_8193;
    wire wire_8194;
    wire wire_8195;
    wire wire_8196;
    wire wire_8197;
    wire wire_8198;
    wire wire_8199;
    wire wire_8200;
    wire wire_8201;
    wire wire_8202;
    wire wire_8203;
    wire wire_8204;
    wire wire_8205;
    wire wire_8206;
    wire wire_8207;
    wire wire_8208;
    wire wire_8209;
    wire wire_8210;
    wire wire_8211;
    wire wire_8212;
    wire wire_8213;
    wire wire_8214;
    wire wire_8215;
    wire wire_8216;
    wire wire_8217;
    wire wire_8218;
    wire wire_8219;
    wire wire_8220;
    wire wire_8221;
    wire wire_8222;
    wire wire_8223;
    wire wire_8224;
    wire wire_8225;
    wire wire_8226;
    wire wire_8227;
    wire wire_8228;
    wire wire_8229;
    wire wire_8230;
    wire wire_8231;
    wire wire_8232;
    wire wire_8233;
    wire wire_8234;
    wire wire_8235;
    wire wire_8236;
    wire wire_8237;
    wire wire_8238;
    wire wire_8239;
    wire wire_8240;
    wire wire_8241;
    wire wire_8242;
    wire wire_8243;
    wire wire_8244;
    wire wire_8245;
    wire wire_8246;
    wire wire_8247;
    wire wire_8248;
    wire wire_8249;
    wire wire_8250;
    wire wire_8251;
    wire wire_8252;
    wire wire_8253;
    wire wire_8254;
    wire wire_8255;
    wire wire_8256;
    wire wire_8257;
    wire wire_8258;
    wire wire_8259;
    wire wire_8260;
    wire wire_8261;
    wire wire_8262;
    wire wire_8263;
    wire wire_8264;
    wire wire_8265;
    wire wire_8266;
    wire wire_8267;
    wire wire_8268;
    wire wire_8269;
    wire wire_8270;
    wire wire_8271;
    wire wire_8272;
    wire wire_8273;
    wire wire_8274;
    wire wire_8275;
    wire wire_8276;
    wire wire_8277;
    wire wire_8278;
    wire wire_8279;
    wire wire_8280;
    wire wire_8281;
    wire wire_8282;
    wire wire_8283;
    wire wire_8284;
    wire wire_8285;
    wire wire_8286;
    wire wire_8287;
    wire wire_8288;
    wire wire_8289;
    wire wire_8290;
    wire wire_8291;
    wire wire_8292;
    wire wire_8293;
    wire wire_8294;
    wire wire_8295;
    wire wire_8296;
    wire wire_8297;
    wire wire_8298;
    wire wire_8299;
    wire wire_8300;
    wire wire_8301;
    wire wire_8302;
    wire wire_8303;
    wire wire_8304;
    wire wire_8305;
    wire wire_8306;
    wire wire_8307;
    wire wire_8308;
    wire wire_8309;
    wire wire_8310;
    wire wire_8311;
    wire wire_8312;
    wire wire_8313;
    wire wire_8314;
    wire wire_8315;
    wire wire_8316;
    wire wire_8317;
    wire wire_8318;
    wire wire_8319;
    wire wire_8320;
    wire wire_8321;
    wire wire_8322;
    wire wire_8323;
    wire wire_8324;
    wire wire_8325;
    wire wire_8326;
    wire wire_8327;
    wire wire_8328;
    wire wire_8329;
    wire wire_8330;
    wire wire_8331;
    wire wire_8332;
    wire wire_8333;
    wire wire_8334;
    wire wire_8335;
    wire wire_8336;
    wire wire_8337;
    wire wire_8338;
    wire wire_8339;
    wire wire_8340;
    wire wire_8341;
    wire wire_8342;
    wire wire_8343;
    wire wire_8344;
    wire wire_8345;
    wire wire_8346;
    wire wire_8347;
    wire wire_8348;
    wire wire_8349;
    wire wire_8350;
    wire wire_8351;
    wire wire_8352;
    wire wire_8353;
    wire wire_8354;
    wire wire_8355;
    wire wire_8356;
    wire wire_8357;
    wire wire_8358;
    wire wire_8359;
    wire wire_8360;
    wire wire_8361;
    wire wire_8362;
    wire wire_8363;
    wire wire_8364;
    wire wire_8365;
    wire wire_8366;
    wire wire_8367;
    wire wire_8368;
    wire wire_8369;
    wire wire_8370;
    wire wire_8371;
    wire wire_8372;
    wire wire_8373;
    wire wire_8374;
    wire wire_8375;
    wire wire_8376;
    wire wire_8377;
    wire wire_8378;
    wire wire_8379;
    wire wire_8380;
    wire wire_8381;
    wire wire_8382;
    wire wire_8383;
    wire wire_8384;
    wire wire_8385;
    wire wire_8386;
    wire wire_8387;
    wire wire_8388;
    wire wire_8389;
    wire wire_8390;
    wire wire_8391;
    wire wire_8392;
    wire wire_8393;
    wire wire_8394;
    wire wire_8395;
    wire wire_8396;
    wire wire_8397;
    wire wire_8398;
    wire wire_8399;
    wire wire_8400;
    wire wire_8401;
    wire wire_8402;
    wire wire_8403;
    wire wire_8404;
    wire wire_8405;
    wire wire_8406;
    wire wire_8407;
    wire wire_8408;
    wire wire_8409;
    wire wire_8410;
    wire wire_8411;
    wire wire_8412;
    wire wire_8413;
    wire wire_8414;
    wire wire_8415;
    wire wire_8416;
    wire wire_8417;
    wire wire_8418;
    wire wire_8419;
    wire wire_8420;
    wire wire_8421;
    wire wire_8422;
    wire wire_8423;
    wire wire_8424;
    wire wire_8425;
    wire wire_8426;
    wire wire_8427;
    wire wire_8428;
    wire wire_8429;
    wire wire_8430;
    wire wire_8431;
    wire wire_8432;
    wire wire_8433;
    wire wire_8434;
    wire wire_8435;
    wire wire_8436;
    wire wire_8437;
    wire wire_8438;
    wire wire_8439;
    wire wire_8440;
    wire wire_8441;
    wire wire_8442;
    wire wire_8443;
    wire wire_8444;
    wire wire_8445;
    wire wire_8446;
    wire wire_8447;
    wire wire_8448;
    wire wire_8449;
    wire wire_8450;
    wire wire_8451;
    wire wire_8452;
    wire wire_8453;
    wire wire_8454;
    wire wire_8455;
    wire wire_8456;
    wire wire_8457;
    wire wire_8458;
    wire wire_8459;
    wire wire_8460;
    wire wire_8461;
    wire wire_8462;
    wire wire_8463;
    wire wire_8464;
    wire wire_8465;
    wire wire_8466;
    wire wire_8467;
    wire wire_8468;
    wire wire_8469;
    wire wire_8470;
    wire wire_8471;
    wire wire_8472;
    wire wire_8473;
    wire wire_8474;
    wire wire_8475;
    wire wire_8476;
    wire wire_8477;
    wire wire_8478;
    wire wire_8479;
    wire wire_8480;
    wire wire_8481;
    wire wire_8482;
    wire wire_8483;
    wire wire_8484;
    wire wire_8485;
    wire wire_8486;
    wire wire_8487;
    wire wire_8488;
    wire wire_8489;
    wire wire_8490;
    wire wire_8491;
    wire wire_8492;
    wire wire_8493;
    wire wire_8494;
    wire wire_8495;
    wire wire_8496;
    wire wire_8497;
    wire wire_8498;
    wire wire_8499;
    wire wire_8500;
    wire wire_8501;
    wire wire_8502;
    wire wire_8503;
    wire wire_8504;
    wire wire_8505;
    wire wire_8506;
    wire wire_8507;
    wire wire_8508;
    wire wire_8509;
    wire wire_8510;
    wire wire_8511;
    wire wire_8512;
    wire wire_8513;
    wire wire_8514;
    wire wire_8515;
    wire wire_8516;
    wire wire_8517;
    wire wire_8518;
    wire wire_8519;
    wire wire_8520;
    wire wire_8521;
    wire wire_8522;
    wire wire_8523;
    wire wire_8524;
    wire wire_8525;
    wire wire_8526;
    wire wire_8527;
    wire wire_8528;
    wire wire_8529;
    wire wire_8530;
    wire wire_8531;
    wire wire_8532;
    wire wire_8533;
    wire wire_8534;
    wire wire_8535;
    wire wire_8536;
    wire wire_8537;
    wire wire_8538;
    wire wire_8539;
    wire wire_8540;
    wire wire_8541;
    wire wire_8542;
    wire wire_8543;
    wire wire_8544;
    wire wire_8545;
    wire wire_8546;
    wire wire_8547;
    wire wire_8548;
    wire wire_8549;
    wire wire_8550;
    wire wire_8551;
    wire wire_8552;
    wire wire_8553;
    wire wire_8554;
    wire wire_8555;
    wire wire_8556;
    wire wire_8557;
    wire wire_8558;
    wire wire_8559;
    wire wire_8560;
    wire wire_8561;
    wire wire_8562;
    wire wire_8563;
    wire wire_8564;
    wire wire_8565;
    wire wire_8566;
    wire wire_8567;
    wire wire_8568;
    wire wire_8569;
    wire wire_8570;
    wire wire_8571;
    wire wire_8572;
    wire wire_8573;
    wire wire_8574;
    wire wire_8575;
    wire wire_8576;
    wire wire_8577;
    wire wire_8578;
    wire wire_8579;
    wire wire_8580;
    wire wire_8581;
    wire wire_8582;
    wire wire_8583;
    wire wire_8584;
    wire wire_8585;
    wire wire_8586;
    wire wire_8587;
    wire wire_8588;
    wire wire_8589;
    wire wire_8590;
    wire wire_8591;
    wire wire_8592;
    wire wire_8593;
    wire wire_8594;
    wire wire_8595;
    wire wire_8596;
    wire wire_8597;
    wire wire_8598;
    wire wire_8599;
    wire wire_8600;
    wire wire_8601;
    wire wire_8602;
    wire wire_8603;
    wire wire_8604;
    wire wire_8605;
    wire wire_8606;
    wire wire_8607;
    wire wire_8608;
    wire wire_8609;
    wire wire_8610;
    wire wire_8611;
    wire wire_8612;
    wire wire_8613;
    wire wire_8614;
    wire wire_8615;
    wire wire_8616;
    wire wire_8617;
    wire wire_8618;
    wire wire_8619;
    wire wire_8620;
    wire wire_8621;
    wire wire_8622;
    wire wire_8623;
    wire wire_8624;
    wire wire_8625;
    wire wire_8626;
    wire wire_8627;
    wire wire_8628;
    wire wire_8629;
    wire wire_8630;
    wire wire_8631;
    wire wire_8632;
    wire wire_8633;
    wire wire_8634;
    wire wire_8635;
    wire wire_8636;
    wire wire_8637;
    wire wire_8638;
    wire wire_8639;
    wire wire_8640;
    wire wire_8641;
    wire wire_8642;
    wire wire_8643;
    wire wire_8644;
    wire wire_8645;
    wire wire_8646;
    wire wire_8647;
    wire wire_8648;
    wire wire_8649;
    wire wire_8650;
    wire wire_8651;
    wire wire_8652;
    wire wire_8653;
    wire wire_8654;
    wire wire_8655;
    wire wire_8656;
    wire wire_8657;
    wire wire_8658;
    wire wire_8659;
    wire wire_8660;
    wire wire_8661;
    wire wire_8662;
    wire wire_8663;
    wire wire_8664;
    wire wire_8665;
    wire wire_8666;
    wire wire_8667;
    wire wire_8668;
    wire wire_8669;
    wire wire_8670;
    wire wire_8671;
    wire wire_8672;
    wire wire_8673;
    wire wire_8674;
    wire wire_8675;
    wire wire_8676;
    wire wire_8677;
    wire wire_8678;
    wire wire_8679;
    wire wire_8680;
    wire wire_8681;
    wire wire_8682;
    wire wire_8683;
    wire wire_8684;
    wire wire_8685;
    wire wire_8686;
    wire wire_8687;
    wire wire_8688;
    wire wire_8689;
    wire wire_8690;
    wire wire_8691;
    wire wire_8692;
    wire wire_8693;
    wire wire_8694;
    wire wire_8695;
    wire wire_8696;
    wire wire_8697;
    wire wire_8698;
    wire wire_8699;
    wire wire_8700;
    wire wire_8701;
    wire wire_8702;
    wire wire_8703;
    wire wire_8704;
    wire wire_8705;
    wire wire_8706;
    wire wire_8707;
    wire wire_8708;
    wire wire_8709;
    wire wire_8710;
    wire wire_8711;
    wire wire_8712;
    wire wire_8713;
    wire wire_8714;
    wire wire_8715;
    wire wire_8716;
    wire wire_8717;
    wire wire_8718;
    wire wire_8719;
    wire wire_8720;
    wire wire_8721;
    wire wire_8722;
    wire wire_8723;
    wire wire_8724;
    wire wire_8725;
    wire wire_8726;
    wire wire_8727;
    wire wire_8728;
    wire wire_8729;
    wire wire_8730;
    wire wire_8731;
    wire wire_8732;
    wire wire_8733;
    wire wire_8734;
    wire wire_8735;
    wire wire_8736;
    wire wire_8737;
    wire wire_8738;
    wire wire_8739;
    wire wire_8740;
    wire wire_8741;
    wire wire_8742;
    wire wire_8743;
    wire wire_8744;
    wire wire_8745;
    wire wire_8746;
    wire wire_8747;
    wire wire_8748;
    wire wire_8749;
    wire wire_8750;
    wire wire_8751;
    wire wire_8752;
    wire wire_8753;
    wire wire_8754;
    wire wire_8755;
    wire wire_8756;
    wire wire_8757;
    wire wire_8758;
    wire wire_8759;
    wire wire_8760;
    wire wire_8761;
    wire wire_8762;
    wire wire_8763;
    wire wire_8764;
    wire wire_8765;
    wire wire_8766;
    wire wire_8767;
    wire wire_8768;
    wire wire_8769;
    wire wire_8770;
    wire wire_8771;
    wire wire_8772;
    wire wire_8773;
    wire wire_8774;
    wire wire_8775;
    wire wire_8776;
    wire wire_8777;
    wire wire_8778;
    wire wire_8779;
    wire wire_8780;
    wire wire_8781;
    wire wire_8782;
    wire wire_8783;
    wire wire_8784;
    wire wire_8785;
    wire wire_8786;
    wire wire_8787;
    wire wire_8788;
    wire wire_8789;
    wire wire_8790;
    wire wire_8791;
    wire wire_8792;
    wire wire_8793;
    wire wire_8794;
    wire wire_8795;
    wire wire_8796;
    wire wire_8797;
    wire wire_8798;
    wire wire_8799;
    wire wire_8800;
    wire wire_8801;
    wire wire_8802;
    wire wire_8803;
    wire wire_8804;
    wire wire_8805;
    wire wire_8806;
    wire wire_8807;
    wire wire_8808;
    wire wire_8809;
    wire wire_8810;
    wire wire_8811;
    wire wire_8812;
    wire wire_8813;
    wire wire_8814;
    wire wire_8815;
    wire wire_8816;
    wire wire_8817;
    wire wire_8818;
    wire wire_8819;
    wire wire_8820;
    wire wire_8821;
    wire wire_8822;
    wire wire_8823;
    wire wire_8824;
    wire wire_8825;
    wire wire_8826;
    wire wire_8827;
    wire wire_8828;
    wire wire_8829;
    wire wire_8830;
    wire wire_8831;
    wire wire_8832;
    wire wire_8833;
    wire wire_8834;
    wire wire_8835;
    wire wire_8836;
    wire wire_8837;
    wire wire_8838;
    wire wire_8839;
    wire wire_8840;
    wire wire_8841;
    wire wire_8842;
    wire wire_8843;
    wire wire_8844;
    wire wire_8845;
    wire wire_8846;
    wire wire_8847;
    wire wire_8848;
    wire wire_8849;
    wire wire_8850;
    wire wire_8851;
    wire wire_8852;
    wire wire_8853;
    wire wire_8854;
    wire wire_8855;
    wire wire_8856;
    wire wire_8857;
    wire wire_8858;
    wire wire_8859;
    wire wire_8860;
    wire wire_8861;
    wire wire_8862;
    wire wire_8863;
    wire wire_8864;
    wire wire_8865;
    wire wire_8866;
    wire wire_8867;
    wire wire_8868;
    wire wire_8869;
    wire wire_8870;
    wire wire_8871;
    wire wire_8872;
    wire wire_8873;
    wire wire_8874;
    wire wire_8875;
    wire wire_8876;
    wire wire_8877;
    wire wire_8878;
    wire wire_8879;
    wire wire_8880;
    wire wire_8881;
    wire wire_8882;
    wire wire_8883;
    wire wire_8884;
    wire wire_8885;
    wire wire_8886;
    wire wire_8887;
    wire wire_8888;
    wire wire_8889;
    wire wire_8890;
    wire wire_8891;
    wire wire_8892;
    wire wire_8893;
    wire wire_8894;
    wire wire_8895;
    wire wire_8896;
    wire wire_8897;
    wire wire_8898;
    wire wire_8899;
    wire wire_8900;
    wire wire_8901;
    wire wire_8902;
    wire wire_8903;
    wire wire_8904;
    wire wire_8905;
    wire wire_8906;
    wire wire_8907;
    wire wire_8908;
    wire wire_8909;
    wire wire_8910;
    wire wire_8911;
    wire wire_8912;
    wire wire_8913;
    wire wire_8914;
    wire wire_8915;
    wire wire_8916;
    wire wire_8917;
    wire wire_8918;
    wire wire_8919;
    wire wire_8920;
    wire wire_8921;
    wire wire_8922;
    wire wire_8923;
    wire wire_8924;
    wire wire_8925;
    wire wire_8926;
    wire wire_8927;
    wire wire_8928;
    wire wire_8929;
    wire wire_8930;
    wire wire_8931;
    wire wire_8932;
    wire wire_8933;
    wire wire_8934;
    wire wire_8935;
    wire wire_8936;
    wire wire_8937;
    wire wire_8938;
    wire wire_8939;
    wire wire_8940;
    wire wire_8941;
    wire wire_8942;
    wire wire_8943;
    wire wire_8944;
    wire wire_8945;
    wire wire_8946;
    wire wire_8947;
    wire wire_8948;
    wire wire_8949;
    wire wire_8950;
    wire wire_8951;
    wire wire_8952;
    wire wire_8953;
    wire wire_8954;
    wire wire_8955;
    wire wire_8956;
    wire wire_8957;
    wire wire_8958;
    wire wire_8959;
    wire wire_8960;
    wire wire_8961;
    wire wire_8962;
    wire wire_8963;
    wire wire_8964;
    wire wire_8965;
    wire wire_8966;
    wire wire_8967;
    wire wire_8968;
    wire wire_8969;
    wire wire_8970;
    wire wire_8971;
    wire wire_8972;
    wire wire_8973;
    wire wire_8974;
    wire wire_8975;
    wire wire_8976;
    wire wire_8977;
    wire wire_8978;
    wire wire_8979;
    wire wire_8980;
    wire wire_8981;
    wire wire_8982;
    wire wire_8983;
    wire wire_8984;
    wire wire_8985;
    wire wire_8986;
    wire wire_8987;
    wire wire_8988;
    wire wire_8989;
    wire wire_8990;
    wire wire_8991;
    wire wire_8992;
    wire wire_8993;
    wire wire_8994;
    wire wire_8995;
    wire wire_8996;
    wire wire_8997;
    wire wire_8998;
    wire wire_8999;
    wire wire_9000;
    wire wire_9001;
    wire wire_9002;
    wire wire_9003;
    wire wire_9004;
    wire wire_9005;
    wire wire_9006;
    wire wire_9007;
    wire wire_9008;
    wire wire_9009;
    wire wire_9010;
    wire wire_9011;
    wire wire_9012;
    wire wire_9013;
    wire wire_9014;
    wire wire_9015;
    wire wire_9016;
    wire wire_9017;
    wire wire_9018;
    wire wire_9019;
    wire wire_9020;
    wire wire_9021;
    wire wire_9022;
    wire wire_9023;
    wire wire_9024;
    wire wire_9025;
    wire wire_9026;
    wire wire_9027;
    wire wire_9028;
    wire wire_9029;
    wire wire_9030;
    wire wire_9031;
    wire wire_9032;
    wire wire_9033;
    wire wire_9034;
    wire wire_9035;
    wire wire_9036;
    wire wire_9037;
    wire wire_9038;
    wire wire_9039;
    wire wire_9040;
    wire wire_9041;
    wire wire_9042;
    wire wire_9043;
    wire wire_9044;
    wire wire_9045;
    wire wire_9046;
    wire wire_9047;
    wire wire_9048;
    wire wire_9049;
    wire wire_9050;
    wire wire_9051;
    wire wire_9052;
    wire wire_9053;
    wire wire_9054;
    wire wire_9055;
    wire wire_9056;
    wire wire_9057;
    wire wire_9058;
    wire wire_9059;
    wire wire_9060;
    wire wire_9061;
    wire wire_9062;
    wire wire_9063;
    wire wire_9064;
    wire wire_9065;
    wire wire_9066;
    wire wire_9067;
    wire wire_9068;
    wire wire_9069;
    wire wire_9070;
    wire wire_9071;
    wire wire_9072;
    wire wire_9073;
    wire wire_9074;
    wire wire_9075;
    wire wire_9076;
    wire wire_9077;
    wire wire_9078;
    wire wire_9079;
    wire wire_9080;
    wire wire_9081;
    wire wire_9082;
    wire wire_9083;
    wire wire_9084;
    wire wire_9085;
    wire wire_9086;
    wire wire_9087;
    wire wire_9088;
    wire wire_9089;
    wire wire_9090;
    wire wire_9091;
    wire wire_9092;
    wire wire_9093;
    wire wire_9094;
    wire wire_9095;
    wire wire_9096;
    wire wire_9097;
    wire wire_9098;
    wire wire_9099;
    wire wire_9100;
    wire wire_9101;
    wire wire_9102;
    wire wire_9103;
    wire wire_9104;
    wire wire_9105;
    wire wire_9106;
    wire wire_9107;
    wire wire_9108;
    wire wire_9109;
    wire wire_9110;
    wire wire_9111;
    wire wire_9112;
    wire wire_9113;
    wire wire_9114;
    wire wire_9115;
    wire wire_9116;
    wire wire_9117;
    wire wire_9118;
    wire wire_9119;
    wire wire_9120;
    wire wire_9121;
    wire wire_9122;
    wire wire_9123;
    wire wire_9124;
    wire wire_9125;
    wire wire_9126;
    wire wire_9127;
    wire wire_9128;
    wire wire_9129;
    wire wire_9130;
    wire wire_9131;
    wire wire_9132;
    wire wire_9133;
    wire wire_9134;
    wire wire_9135;
    wire wire_9136;
    wire wire_9137;
    wire wire_9138;
    wire wire_9139;
    wire wire_9140;
    wire wire_9141;
    wire wire_9142;
    wire wire_9143;
    wire wire_9144;
    wire wire_9145;
    wire wire_9146;
    wire wire_9147;
    wire wire_9148;
    wire wire_9149;
    wire wire_9150;
    wire wire_9151;
    wire wire_9152;
    wire wire_9153;
    wire wire_9154;
    wire wire_9155;
    wire wire_9156;
    wire wire_9157;
    wire wire_9158;
    wire wire_9159;
    wire wire_9160;
    wire wire_9161;
    wire wire_9162;
    wire wire_9163;
    wire wire_9164;
    wire wire_9165;
    wire wire_9166;
    wire wire_9167;
    wire wire_9168;
    wire wire_9169;
    wire wire_9170;
    wire wire_9171;
    wire wire_9172;
    wire wire_9173;
    wire wire_9174;
    wire wire_9175;
    wire wire_9176;
    wire wire_9177;
    wire wire_9178;
    wire wire_9179;
    wire wire_9180;
    wire wire_9181;
    wire wire_9182;
    wire wire_9183;
    wire wire_9184;
    wire wire_9185;
    wire wire_9186;
    wire wire_9187;
    wire wire_9188;
    wire wire_9189;
    wire wire_9190;
    wire wire_9191;
    wire wire_9192;
    wire wire_9193;
    wire wire_9194;
    wire wire_9195;
    wire wire_9196;
    wire wire_9197;
    wire wire_9198;
    wire wire_9199;
    wire wire_9200;
    wire wire_9201;
    wire wire_9202;
    wire wire_9203;
    wire wire_9204;
    wire wire_9205;
    wire wire_9206;
    wire wire_9207;
    wire wire_9208;
    wire wire_9209;
    wire wire_9210;
    wire wire_9211;
    wire wire_9212;
    wire wire_9213;
    wire wire_9214;
    wire wire_9215;
    wire wire_9216;
    wire wire_9217;
    wire wire_9218;
    wire wire_9219;
    wire wire_9220;
    wire wire_9221;
    wire wire_9222;
    wire wire_9223;
    wire wire_9224;
    wire wire_9225;
    wire wire_9226;
    wire wire_9227;
    wire wire_9228;
    wire wire_9229;
    wire wire_9230;
    wire wire_9231;
    wire wire_9232;
    wire wire_9233;
    wire wire_9234;
    wire wire_9235;
    wire wire_9236;
    wire wire_9237;
    wire wire_9238;
    wire wire_9239;
    wire wire_9240;
    wire wire_9241;
    wire wire_9242;
    wire wire_9243;
    wire wire_9244;
    wire wire_9245;
    wire wire_9246;
    wire wire_9247;
    wire wire_9248;
    wire wire_9249;
    wire wire_9250;
    wire wire_9251;
    wire wire_9252;
    wire wire_9253;
    wire wire_9254;
    wire wire_9255;
    wire wire_9256;
    wire wire_9257;
    wire wire_9258;
    wire wire_9259;
    wire wire_9260;
    wire wire_9261;
    wire wire_9262;
    wire wire_9263;
    wire wire_9264;
    wire wire_9265;
    wire wire_9266;
    wire wire_9267;
    wire wire_9268;
    wire wire_9269;
    wire wire_9270;
    wire wire_9271;
    wire wire_9272;
    wire wire_9273;
    wire wire_9274;
    wire wire_9275;
    wire wire_9276;
    wire wire_9277;
    wire wire_9278;
    wire wire_9279;
    wire wire_9280;
    wire wire_9281;
    wire wire_9282;
    wire wire_9283;
    wire wire_9284;
    wire wire_9285;
    wire wire_9286;
    wire wire_9287;
    wire wire_9288;
    wire wire_9289;
    wire wire_9290;
    wire wire_9291;
    wire wire_9292;
    wire wire_9293;
    wire wire_9294;
    wire wire_9295;
    wire wire_9296;
    wire wire_9297;
    wire wire_9298;
    wire wire_9299;
    wire wire_9300;
    wire wire_9301;
    wire wire_9302;
    wire wire_9303;
    wire wire_9304;
    wire wire_9305;
    wire wire_9306;
    wire wire_9307;
    wire wire_9308;
    wire wire_9309;
    wire wire_9310;
    wire wire_9311;
    wire wire_9312;
    wire wire_9313;
    wire wire_9314;
    wire wire_9315;
    wire wire_9316;
    wire wire_9317;
    wire wire_9318;
    wire wire_9319;
    wire wire_9320;
    wire wire_9321;
    wire wire_9322;
    wire wire_9323;
    wire wire_9324;
    wire wire_9325;
    wire wire_9326;
    wire wire_9327;
    wire wire_9328;
    wire wire_9329;
    wire wire_9330;
    wire wire_9331;
    wire wire_9332;
    wire wire_9333;
    wire wire_9334;
    wire wire_9335;
    wire wire_9336;
    wire wire_9337;
    wire wire_9338;
    wire wire_9339;
    wire wire_9340;
    wire wire_9341;
    wire wire_9342;
    wire wire_9343;
    wire wire_9344;
    wire wire_9345;
    wire wire_9346;
    wire wire_9347;
    wire wire_9348;
    wire wire_9349;
    wire wire_9350;
    wire wire_9351;
    wire wire_9352;
    wire wire_9353;
    wire wire_9354;
    wire wire_9355;
    wire wire_9356;
    wire wire_9357;
    wire wire_9358;
    wire wire_9359;
    wire wire_9360;
    wire wire_9361;
    wire wire_9362;
    wire wire_9363;
    wire wire_9364;
    wire wire_9365;
    wire wire_9366;
    wire wire_9367;
    wire wire_9368;
    wire wire_9369;
    wire wire_9370;
    wire wire_9371;
    wire wire_9372;
    wire wire_9373;
    wire wire_9374;
    wire wire_9375;
    wire wire_9376;
    wire wire_9377;
    wire wire_9378;
    wire wire_9379;
    wire wire_9380;
    wire wire_9381;
    wire wire_9382;
    wire wire_9383;
    wire wire_9384;
    wire wire_9385;
    wire wire_9386;
    wire wire_9387;
    wire wire_9388;
    wire wire_9389;
    wire wire_9390;
    wire wire_9391;
    wire wire_9392;
    wire wire_9393;
    wire wire_9394;
    wire wire_9395;
    wire wire_9396;
    wire wire_9397;
    wire wire_9398;
    wire wire_9399;
    wire wire_9400;
    wire wire_9401;
    wire wire_9402;
    wire wire_9403;
    wire wire_9404;
    wire wire_9405;
    wire wire_9406;
    wire wire_9407;
    wire wire_9408;
    wire wire_9409;
    wire wire_9410;
    wire wire_9411;
    wire wire_9412;
    wire wire_9413;
    wire wire_9414;
    wire wire_9415;
    wire wire_9416;
    wire wire_9417;
    wire wire_9418;
    wire wire_9419;
    wire wire_9420;
    wire wire_9421;
    wire wire_9422;
    wire wire_9423;
    wire wire_9424;
    wire wire_9425;
    wire wire_9426;
    wire wire_9427;
    wire wire_9428;
    wire wire_9429;
    wire wire_9430;
    wire wire_9431;
    wire wire_9432;
    wire wire_9433;
    wire wire_9434;
    wire wire_9435;
    wire wire_9436;
    wire wire_9437;
    wire wire_9438;
    wire wire_9439;
    wire wire_9440;
    wire wire_9441;
    wire wire_9442;
    wire wire_9443;
    wire wire_9444;
    wire wire_9445;
    wire wire_9446;
    wire wire_9447;
    wire wire_9448;
    wire wire_9449;
    wire wire_9450;
    wire wire_9451;
    wire wire_9452;
    wire wire_9453;
    wire wire_9454;
    wire wire_9455;
    wire wire_9456;
    wire wire_9457;
    wire wire_9458;
    wire wire_9459;
    wire wire_9460;
    wire wire_9461;
    wire wire_9462;
    wire wire_9463;
    wire wire_9464;
    wire wire_9465;
    wire wire_9466;
    wire wire_9467;
    wire wire_9468;
    wire wire_9469;
    wire wire_9470;
    wire wire_9471;
    wire wire_9472;
    wire wire_9473;
    wire wire_9474;
    wire wire_9475;
    wire wire_9476;
    wire wire_9477;
    wire wire_9478;
    wire wire_9479;
    wire wire_9480;
    wire wire_9481;
    wire wire_9482;
    wire wire_9483;
    wire wire_9484;
    wire wire_9485;
    wire wire_9486;
    wire wire_9487;
    wire wire_9488;
    wire wire_9489;
    wire wire_9490;
    wire wire_9491;
    wire wire_9492;
    wire wire_9493;
    wire wire_9494;
    wire wire_9495;
    wire wire_9496;
    wire wire_9497;
    wire wire_9498;
    wire wire_9499;
    wire wire_9500;
    wire wire_9501;
    wire wire_9502;
    wire wire_9503;
    wire wire_9504;
    wire wire_9505;
    wire wire_9506;
    wire wire_9507;
    wire wire_9508;
    wire wire_9509;
    wire wire_9510;
    wire wire_9511;
    wire wire_9512;
    wire wire_9513;
    wire wire_9514;
    wire wire_9515;
    wire wire_9516;
    wire wire_9517;
    wire wire_9518;
    wire wire_9519;
    wire wire_9520;
    wire wire_9521;
    wire wire_9522;
    wire wire_9523;
    wire wire_9524;
    wire wire_9525;
    wire wire_9526;
    wire wire_9527;
    wire wire_9528;
    wire wire_9529;
    wire wire_9530;
    wire wire_9531;
    wire wire_9532;
    wire wire_9533;
    wire wire_9534;
    wire wire_9535;
    wire wire_9536;
    wire wire_9537;
    wire wire_9538;
    wire wire_9539;
    wire wire_9540;
    wire wire_9541;
    wire wire_9542;
    wire wire_9543;
    wire wire_9544;
    wire wire_9545;
    wire wire_9546;
    wire wire_9547;
    wire wire_9548;
    wire wire_9549;
    wire wire_9550;
    wire wire_9551;
    wire wire_9552;
    wire wire_9553;
    wire wire_9554;
    wire wire_9555;
    wire wire_9556;
    wire wire_9557;
    wire wire_9558;
    wire wire_9559;
    wire wire_9560;
    wire wire_9561;
    wire wire_9562;
    wire wire_9563;
    wire wire_9564;
    wire wire_9565;
    wire wire_9566;
    wire wire_9567;
    wire wire_9568;
    wire wire_9569;
    wire wire_9570;
    wire wire_9571;
    wire wire_9572;
    wire wire_9573;
    wire wire_9574;
    wire wire_9575;
    wire wire_9576;
    wire wire_9577;
    wire wire_9578;
    wire wire_9579;
    wire wire_9580;
    wire wire_9581;
    wire wire_9582;
    wire wire_9583;
    wire wire_9584;
    wire wire_9585;
    wire wire_9586;
    wire wire_9587;
    wire wire_9588;
    wire wire_9589;
    wire wire_9590;
    wire wire_9591;
    wire wire_9592;
    wire wire_9593;
    wire wire_9594;
    wire wire_9595;
    wire wire_9596;
    wire wire_9597;
    wire wire_9598;
    wire wire_9599;
    wire wire_9600;
    wire wire_9601;
    wire wire_9602;
    wire wire_9603;
    wire wire_9604;
    wire wire_9605;
    wire wire_9606;
    wire wire_9607;
    wire wire_9608;
    wire wire_9609;
    wire wire_9610;
    wire wire_9611;
    wire wire_9612;
    wire wire_9613;
    wire wire_9614;
    wire wire_9615;
    wire wire_9616;
    wire wire_9617;
    wire wire_9618;
    wire wire_9619;
    wire wire_9620;
    wire wire_9621;
    wire wire_9622;
    wire wire_9623;
    wire wire_9624;
    wire wire_9625;
    wire wire_9626;
    wire wire_9627;
    wire wire_9628;
    wire wire_9629;
    wire wire_9630;
    wire wire_9631;
    wire wire_9632;
    wire wire_9633;
    wire wire_9634;
    wire wire_9635;
    wire wire_9636;
    wire wire_9637;
    wire wire_9638;
    wire wire_9639;
    wire wire_9640;
    wire wire_9641;
    wire wire_9642;
    wire wire_9643;
    wire wire_9644;
    wire wire_9645;
    wire wire_9646;
    wire wire_9647;
    wire wire_9648;
    wire wire_9649;
    wire wire_9650;
    wire wire_9651;
    wire wire_9652;
    wire wire_9653;
    wire wire_9654;
    wire wire_9655;
    wire wire_9656;
    wire wire_9657;
    wire wire_9658;
    wire wire_9659;
    wire wire_9660;
    wire wire_9661;
    wire wire_9662;
    wire wire_9663;
    wire wire_9664;
    wire wire_9665;
    wire wire_9666;
    wire wire_9667;
    wire wire_9668;
    wire wire_9669;
    wire wire_9670;
    wire wire_9671;
    wire wire_9672;
    wire wire_9673;
    wire wire_9674;
    wire wire_9675;
    wire wire_9676;
    wire wire_9677;
    wire wire_9678;
    wire wire_9679;
    wire wire_9680;
    wire wire_9681;
    wire wire_9682;
    wire wire_9683;
    wire wire_9684;
    wire wire_9685;
    wire wire_9686;
    wire wire_9687;
    wire wire_9688;
    wire wire_9689;
    wire wire_9690;
    wire wire_9691;
    wire wire_9692;
    wire wire_9693;
    wire wire_9694;
    wire wire_9695;
    wire wire_9696;
    wire wire_9697;
    wire wire_9698;
    wire wire_9699;
    wire wire_9700;
    wire wire_9701;
    wire wire_9702;
    wire wire_9703;
    wire wire_9704;
    wire wire_9705;
    wire wire_9706;
    wire wire_9707;
    wire wire_9708;
    wire wire_9709;
    wire wire_9710;
    wire wire_9711;
    wire wire_9712;
    wire wire_9713;
    wire wire_9714;
    wire wire_9715;
    wire wire_9716;
    wire wire_9717;
    wire wire_9718;
    wire wire_9719;
    wire wire_9720;
    wire wire_9721;
    wire wire_9722;
    wire wire_9723;
    wire wire_9724;
    wire wire_9725;
    wire wire_9726;
    wire wire_9727;
    wire wire_9728;
    wire wire_9729;
    wire wire_9730;
    wire wire_9731;
    wire wire_9732;
    wire wire_9733;
    wire wire_9734;
    wire wire_9735;
    wire wire_9736;
    wire wire_9737;
    wire wire_9738;
    wire wire_9739;
    wire wire_9740;
    wire wire_9741;
    wire wire_9742;
    wire wire_9743;
    wire wire_9744;
    wire wire_9745;
    wire wire_9746;
    wire wire_9747;
    wire wire_9748;
    wire wire_9749;
    wire wire_9750;
    wire wire_9751;
    wire wire_9752;
    wire wire_9753;
    wire wire_9754;
    wire wire_9755;
    wire wire_9756;
    wire wire_9757;
    wire wire_9758;
    wire wire_9759;
    wire wire_9760;
    wire wire_9761;
    wire wire_9762;
    wire wire_9763;
    wire wire_9764;
    wire wire_9765;
    wire wire_9766;
    wire wire_9767;
    wire wire_9768;
    wire wire_9769;
    wire wire_9770;
    wire wire_9771;
    wire wire_9772;
    wire wire_9773;
    wire wire_9774;
    wire wire_9775;
    wire wire_9776;
    wire wire_9777;
    wire wire_9778;
    wire wire_9779;
    wire wire_9780;
    wire wire_9781;
    wire wire_9782;
    wire wire_9783;
    wire wire_9784;
    wire wire_9785;
    wire wire_9786;
    wire wire_9787;
    wire wire_9788;
    wire wire_9789;
    wire wire_9790;
    wire wire_9791;
    wire wire_9792;
    wire wire_9793;
    wire wire_9794;
    wire wire_9795;
    wire wire_9796;
    wire wire_9797;
    wire wire_9798;
    wire wire_9799;
    wire wire_9800;
    wire wire_9801;
    wire wire_9802;
    wire wire_9803;
    wire wire_9804;
    wire wire_9805;
    wire wire_9806;
    wire wire_9807;
    wire wire_9808;
    wire wire_9809;
    wire wire_9810;
    wire wire_9811;
    wire wire_9812;
    wire wire_9813;
    wire wire_9814;
    wire wire_9815;
    wire wire_9816;
    wire wire_9817;
    wire wire_9818;
    wire wire_9819;
    wire wire_9820;
    wire wire_9821;
    wire wire_9822;
    wire wire_9823;
    wire wire_9824;
    wire wire_9825;
    wire wire_9826;
    wire wire_9827;
    wire wire_9828;
    wire wire_9829;
    wire wire_9830;
    wire wire_9831;
    wire wire_9832;
    wire wire_9833;
    wire wire_9834;
    wire wire_9835;
    wire wire_9836;
    wire wire_9837;
    wire wire_9838;
    wire wire_9839;
    wire wire_9840;
    wire wire_9841;
    wire wire_9842;
    wire wire_9843;
    wire wire_9844;
    wire wire_9845;
    wire wire_9846;
    wire wire_9847;
    wire wire_9848;
    wire wire_9849;
    wire wire_9850;
    wire wire_9851;
    wire wire_9852;
    wire wire_9853;
    wire wire_9854;
    wire wire_9855;
    wire wire_9856;
    wire wire_9857;
    wire wire_9858;
    wire wire_9859;
    wire wire_9860;
    wire wire_9861;
    wire wire_9862;
    wire wire_9863;
    wire wire_9864;
    wire wire_9865;
    wire wire_9866;
    wire wire_9867;
    wire wire_9868;
    wire wire_9869;
    wire wire_9870;
    wire wire_9871;
    wire wire_9872;
    wire wire_9873;
    wire wire_9874;
    wire wire_9875;
    wire wire_9876;
    wire wire_9877;
    wire wire_9878;
    wire wire_9879;
    wire wire_9880;
    wire wire_9881;
    wire wire_9882;
    wire wire_9883;
    wire wire_9884;
    wire wire_9885;
    wire wire_9886;
    wire wire_9887;
    wire wire_9888;
    wire wire_9889;
    wire wire_9890;
    wire wire_9891;
    wire wire_9892;
    wire wire_9893;
    wire wire_9894;
    wire wire_9895;
    wire wire_9896;
    wire wire_9897;
    wire wire_9898;
    wire wire_9899;
    wire wire_9900;
    wire wire_9901;
    wire wire_9902;
    wire wire_9903;
    wire wire_9904;
    wire wire_9905;
    wire wire_9906;
    wire wire_9907;
    wire wire_9908;
    wire wire_9909;
    wire wire_9910;
    wire wire_9911;
    wire wire_9912;
    wire wire_9913;
    wire wire_9914;
    wire wire_9915;
    wire wire_9916;
    wire wire_9917;
    wire wire_9918;
    wire wire_9919;
    wire wire_9920;
    wire wire_9921;
    wire wire_9922;
    wire wire_9923;
    wire wire_9924;
    wire wire_9925;
    wire wire_9926;
    wire wire_9927;
    wire wire_9928;
    wire wire_9929;
    wire wire_9930;
    wire wire_9931;
    wire wire_9932;
    wire wire_9933;
    wire wire_9934;
    wire wire_9935;
    wire wire_9936;
    wire wire_9937;
    wire wire_9938;
    wire wire_9939;
    wire wire_9940;
    wire wire_9941;
    wire wire_9942;
    wire wire_9943;
    wire wire_9944;
    wire wire_9945;
    wire wire_9946;
    wire wire_9947;
    wire wire_9948;
    wire wire_9949;
    wire wire_9950;
    wire wire_9951;
    wire wire_9952;
    wire wire_9953;
    wire wire_9954;
    wire wire_9955;
    wire wire_9956;
    wire wire_9957;
    wire wire_9958;
    wire wire_9959;
    wire wire_9960;
    wire wire_9961;
    wire wire_9962;
    wire wire_9963;
    wire wire_9964;
    wire wire_9965;
    wire wire_9966;
    wire wire_9967;
    wire wire_9968;
    wire wire_9969;
    wire wire_9970;
    wire wire_9971;
    wire wire_9972;
    wire wire_9973;
    wire wire_9974;
    wire wire_9975;
    wire wire_9976;
    wire wire_9977;
    wire wire_9978;
    wire wire_9979;
    wire wire_9980;
    wire wire_9981;
    wire wire_9982;
    wire wire_9983;
    wire wire_9984;
    wire wire_9985;
    wire wire_9986;
    wire wire_9987;
    wire wire_9988;
    wire wire_9989;
    wire wire_9990;
    wire wire_9991;
    wire wire_9992;
    wire wire_9993;
    wire wire_9994;
    wire wire_9995;
    wire wire_9996;
    wire wire_9997;
    wire wire_9998;
    wire wire_9999;
    wire wire_10000;
    wire wire_10001;
    wire wire_10002;
    wire wire_10003;
    wire wire_10004;
    wire wire_10005;
    wire wire_10006;
    wire wire_10007;
    wire wire_10008;
    wire wire_10009;
    wire wire_10010;
    wire wire_10011;
    wire wire_10012;
    wire wire_10013;
    wire wire_10014;
    wire wire_10015;
    wire wire_10016;
    wire wire_10017;
    wire wire_10018;
    wire wire_10019;
    wire wire_10020;
    wire wire_10021;
    wire wire_10022;
    wire wire_10023;
    wire wire_10024;
    wire wire_10025;
    wire wire_10026;
    wire wire_10027;
    wire wire_10028;
    wire wire_10029;
    wire wire_10030;
    wire wire_10031;
    wire wire_10032;
    wire wire_10033;
    wire wire_10034;
    wire wire_10035;
    wire wire_10036;
    wire wire_10037;
    wire wire_10038;
    wire wire_10039;
    wire wire_10040;
    wire wire_10041;
    wire wire_10042;
    wire wire_10043;
    wire wire_10044;
    wire wire_10045;
    wire wire_10046;
    wire wire_10047;
    wire wire_10048;
    wire wire_10049;
    wire wire_10050;
    wire wire_10051;
    wire wire_10052;
    wire wire_10053;
    wire wire_10054;
    wire wire_10055;
    wire wire_10056;
    wire wire_10057;
    wire wire_10058;
    wire wire_10059;
    wire wire_10060;
    wire wire_10061;
    wire wire_10062;
    wire wire_10063;
    wire wire_10064;
    wire wire_10065;
    wire wire_10066;
    wire wire_10067;
    wire wire_10068;
    wire wire_10069;
    wire wire_10070;
    wire wire_10071;
    wire wire_10072;
    wire wire_10073;
    wire wire_10074;
    wire wire_10075;
    wire wire_10076;
    wire wire_10077;
    wire wire_10078;
    wire wire_10079;
    wire wire_10080;
    wire wire_10081;
    wire wire_10082;
    wire wire_10083;
    wire wire_10084;
    wire wire_10085;
    wire wire_10086;
    wire wire_10087;
    wire wire_10088;
    wire wire_10089;
    wire wire_10090;
    wire wire_10091;
    wire wire_10092;
    wire wire_10093;
    wire wire_10094;
    wire wire_10095;
    wire wire_10096;
    wire wire_10097;
    wire wire_10098;
    wire wire_10099;
    wire wire_10100;
    wire wire_10101;
    wire wire_10102;
    wire wire_10103;
    wire wire_10104;
    wire wire_10105;
    wire wire_10106;
    wire wire_10107;
    wire wire_10108;
    wire wire_10109;
    wire wire_10110;
    wire wire_10111;
    wire wire_10112;
    wire wire_10113;
    wire wire_10114;
    wire wire_10115;
    wire wire_10116;
    wire wire_10117;
    wire wire_10118;
    wire wire_10119;
    wire wire_10120;
    wire wire_10121;
    wire wire_10122;
    wire wire_10123;
    wire wire_10124;
    wire wire_10125;
    wire wire_10126;
    wire wire_10127;
    wire wire_10128;
    wire wire_10129;
    wire wire_10130;
    wire wire_10131;
    wire wire_10132;
    wire wire_10133;
    wire wire_10134;
    wire wire_10135;
    wire wire_10136;
    wire wire_10137;
    wire wire_10138;
    wire wire_10139;
    wire wire_10140;
    wire wire_10141;
    wire wire_10142;
    wire wire_10143;
    wire wire_10144;
    wire wire_10145;
    wire wire_10146;
    wire wire_10147;
    wire wire_10148;
    wire wire_10149;
    wire wire_10150;
    wire wire_10151;
    wire wire_10152;
    wire wire_10153;
    wire wire_10154;
    wire wire_10155;
    wire wire_10156;
    wire wire_10157;
    wire wire_10158;
    wire wire_10159;
    wire wire_10160;
    wire wire_10161;
    wire wire_10162;
    wire wire_10163;
    wire wire_10164;
    wire wire_10165;
    wire wire_10166;
    wire wire_10167;
    wire wire_10168;
    wire wire_10169;
    wire wire_10170;
    wire wire_10171;
    wire wire_10172;
    wire wire_10173;
    wire wire_10174;
    wire wire_10175;
    wire wire_10176;
    wire wire_10177;
    wire wire_10178;
    wire wire_10179;
    wire wire_10180;
    wire wire_10181;
    wire wire_10182;
    wire wire_10183;
    wire wire_10184;
    wire wire_10185;
    wire wire_10186;
    wire wire_10187;
    wire wire_10188;
    wire wire_10189;
    wire wire_10190;
    wire wire_10191;
    wire wire_10192;
    wire wire_10193;
    wire wire_10194;
    wire wire_10195;
    wire wire_10196;
    wire wire_10197;
    wire wire_10198;
    wire wire_10199;
    wire wire_10200;
    wire wire_10201;
    wire wire_10202;
    wire wire_10203;
    wire wire_10204;
    wire wire_10205;
    wire wire_10206;
    wire wire_10207;
    wire wire_10208;
    wire wire_10209;
    wire wire_10210;
    wire wire_10211;
    wire wire_10212;
    wire wire_10213;
    wire wire_10214;
    wire wire_10215;
    wire wire_10216;
    wire wire_10217;
    wire wire_10218;
    wire wire_10219;
    wire wire_10220;
    wire wire_10221;
    wire wire_10222;
    wire wire_10223;
    wire wire_10224;
    wire wire_10225;
    wire wire_10226;
    wire wire_10227;
    wire wire_10228;
    wire wire_10229;
    wire wire_10230;
    wire wire_10231;
    wire wire_10232;
    wire wire_10233;
    wire wire_10234;
    wire wire_10235;
    wire wire_10236;
    wire wire_10237;
    wire wire_10238;
    wire wire_10239;
    wire wire_10240;
    wire wire_10241;
    wire wire_10242;
    wire wire_10243;
    wire wire_10244;
    wire wire_10245;
    wire wire_10246;
    wire wire_10247;
    wire wire_10248;
    wire wire_10249;
    wire wire_10250;
    wire wire_10251;
    wire wire_10252;
    wire wire_10253;
    wire wire_10254;
    wire wire_10255;
    wire wire_10256;
    wire wire_10257;
    wire wire_10258;
    wire wire_10259;
    wire wire_10260;
    wire wire_10261;
    wire wire_10262;
    wire wire_10263;
    wire wire_10264;
    wire wire_10265;
    wire wire_10266;
    wire wire_10267;
    wire wire_10268;
    wire wire_10269;
    wire wire_10270;
    wire wire_10271;
    wire wire_10272;
    wire wire_10273;
    wire wire_10274;
    wire wire_10275;
    wire wire_10276;
    wire wire_10277;
    wire wire_10278;
    wire wire_10279;
    wire wire_10280;
    wire wire_10281;
    wire wire_10282;
    wire wire_10283;
    wire wire_10284;
    wire wire_10285;
    wire wire_10286;
    wire wire_10287;
    wire wire_10288;
    wire wire_10289;
    wire wire_10290;
    wire wire_10291;
    wire wire_10292;
    wire wire_10293;
    wire wire_10294;
    wire wire_10295;
    wire wire_10296;
    wire wire_10297;
    wire wire_10298;
    wire wire_10299;
    wire wire_10300;
    wire wire_10301;
    wire wire_10302;
    wire wire_10303;
    wire wire_10304;
    wire wire_10305;
    wire wire_10306;
    wire wire_10307;
    wire wire_10308;
    wire wire_10309;
    wire wire_10310;
    wire wire_10311;
    wire wire_10312;
    wire wire_10313;
    wire wire_10314;
    wire wire_10315;
    wire wire_10316;
    wire wire_10317;
    wire wire_10318;
    wire wire_10319;
    wire wire_10320;
    wire wire_10321;
    wire wire_10322;
    wire wire_10323;
    wire wire_10324;
    wire wire_10325;
    wire wire_10326;
    wire wire_10327;
    wire wire_10328;
    wire wire_10329;
    wire wire_10330;
    wire wire_10331;
    wire wire_10332;
    wire wire_10333;
    wire wire_10334;
    wire wire_10335;
    wire wire_10336;
    wire wire_10337;
    wire wire_10338;
    wire wire_10339;
    wire wire_10340;
    wire wire_10341;
    wire wire_10342;
    wire wire_10343;
    wire wire_10344;
    wire wire_10345;
    wire wire_10346;
    wire wire_10347;
    wire wire_10348;
    wire wire_10349;
    wire wire_10350;
    wire wire_10351;
    wire wire_10352;
    wire wire_10353;
    wire wire_10354;
    wire wire_10355;
    wire wire_10356;
    wire wire_10357;
    wire wire_10358;
    wire wire_10359;
    wire wire_10360;
    wire wire_10361;
    wire wire_10362;
    wire wire_10363;
    wire wire_10364;
    wire wire_10365;
    wire wire_10366;
    wire wire_10367;
    wire wire_10368;
    wire wire_10369;
    wire wire_10370;
    wire wire_10371;
    wire wire_10372;
    wire wire_10373;
    wire wire_10374;
    wire wire_10375;
    wire wire_10376;
    wire wire_10377;
    wire wire_10378;
    wire wire_10379;
    wire wire_10380;
    wire wire_10381;
    wire wire_10382;
    wire wire_10383;
    wire wire_10384;
    wire wire_10385;
    wire wire_10386;
    wire wire_10387;
    wire wire_10388;
    wire wire_10389;
    wire wire_10390;
    wire wire_10391;
    wire wire_10392;
    wire wire_10393;
    wire wire_10394;
    wire wire_10395;
    wire wire_10396;
    wire wire_10397;
    wire wire_10398;
    wire wire_10399;
    wire wire_10400;
    wire wire_10401;
    wire wire_10402;
    wire wire_10403;
    wire wire_10404;
    wire wire_10405;
    wire wire_10406;
    wire wire_10407;
    wire wire_10408;
    wire wire_10409;
    wire wire_10410;
    wire wire_10411;
    wire wire_10412;
    wire wire_10413;
    wire wire_10414;
    wire wire_10415;
    wire wire_10416;
    wire wire_10417;
    wire wire_10418;
    wire wire_10419;
    wire wire_10420;
    wire wire_10421;
    wire wire_10422;
    wire wire_10423;
    wire wire_10424;
    wire wire_10425;
    wire wire_10426;
    wire wire_10427;
    wire wire_10428;
    wire wire_10429;
    wire wire_10430;
    wire wire_10431;
    wire wire_10432;
    wire wire_10433;
    wire wire_10434;
    wire wire_10435;
    wire wire_10436;
    wire wire_10437;
    wire wire_10438;
    wire wire_10439;
    wire wire_10440;
    wire wire_10441;
    wire wire_10442;
    wire wire_10443;
    wire wire_10444;
    wire wire_10445;
    wire wire_10446;
    wire wire_10447;
    wire wire_10448;
    wire wire_10449;
    wire wire_10450;
    wire wire_10451;
    wire wire_10452;
    wire wire_10453;
    wire wire_10454;
    wire wire_10455;
    wire wire_10456;
    wire wire_10457;
    wire wire_10458;
    wire wire_10459;
    wire wire_10460;
    wire wire_10461;
    wire wire_10462;
    wire wire_10463;
    wire wire_10464;
    wire wire_10465;
    wire wire_10466;
    wire wire_10467;
    wire wire_10468;
    wire wire_10469;
    wire wire_10470;
    wire wire_10471;
    wire wire_10472;
    wire wire_10473;
    wire wire_10474;
    wire wire_10475;
    wire wire_10476;
    wire wire_10477;
    wire wire_10478;
    wire wire_10479;
    wire wire_10480;
    wire wire_10481;
    wire wire_10482;
    wire wire_10483;
    wire wire_10484;
    wire wire_10485;
    wire wire_10486;
    wire wire_10487;
    wire wire_10488;
    wire wire_10489;
    wire wire_10490;
    wire wire_10491;
    wire wire_10492;
    wire wire_10493;
    wire wire_10494;
    wire wire_10495;
    wire wire_10496;
    wire wire_10497;
    wire wire_10498;
    wire wire_10499;
    wire wire_10500;
    wire wire_10501;
    wire wire_10502;
    wire wire_10503;
    wire wire_10504;
    wire wire_10505;
    wire wire_10506;
    wire wire_10507;
    wire wire_10508;
    wire wire_10509;
    wire wire_10510;
    wire wire_10511;
    wire wire_10512;
    wire wire_10513;
    wire wire_10514;
    wire wire_10515;
    wire wire_10516;
    wire wire_10517;
    wire wire_10518;
    wire wire_10519;
    wire wire_10520;
    wire wire_10521;
    wire wire_10522;
    wire wire_10523;
    wire wire_10524;
    wire wire_10525;
    wire wire_10526;
    wire wire_10527;
    wire wire_10528;
    wire wire_10529;
    wire wire_10530;
    wire wire_10531;
    wire wire_10532;
    wire wire_10533;
    wire wire_10534;
    wire wire_10535;
    wire wire_10536;
    wire wire_10537;
    wire wire_10538;
    wire wire_10539;
    wire wire_10540;
    wire wire_10541;
    wire wire_10542;
    wire wire_10543;
    wire wire_10544;
    wire wire_10545;
    wire wire_10546;
    wire wire_10547;
    wire wire_10548;
    wire wire_10549;
    wire wire_10550;
    wire wire_10551;
    wire wire_10552;
    wire wire_10553;
    wire wire_10554;
    wire wire_10555;
    wire wire_10556;
    wire wire_10557;
    wire wire_10558;
    wire wire_10559;
    wire wire_10560;
    wire wire_10561;
    wire wire_10562;
    wire wire_10563;
    wire wire_10564;
    wire wire_10565;
    wire wire_10566;
    wire wire_10567;
    wire wire_10568;
    wire wire_10569;
    wire wire_10570;
    wire wire_10571;
    wire wire_10572;
    wire wire_10573;
    wire wire_10574;
    wire wire_10575;
    wire wire_10576;
    wire wire_10577;
    wire wire_10578;
    wire wire_10579;
    wire wire_10580;
    wire wire_10581;
    wire wire_10582;
    wire wire_10583;
    wire wire_10584;
    wire wire_10585;
    wire wire_10586;
    wire wire_10587;
    wire wire_10588;
    wire wire_10589;
    wire wire_10590;
    wire wire_10591;
    wire wire_10592;
    wire wire_10593;
    wire wire_10594;
    wire wire_10595;
    wire wire_10596;
    wire wire_10597;
    wire wire_10598;
    wire wire_10599;
    wire wire_10600;
    wire wire_10601;
    wire wire_10602;
    wire wire_10603;
    wire wire_10604;
    wire wire_10605;
    wire wire_10606;
    wire wire_10607;
    wire wire_10608;
    wire wire_10609;
    wire wire_10610;
    wire wire_10611;
    wire wire_10612;
    wire wire_10613;
    wire wire_10614;
    wire wire_10615;
    wire wire_10616;
    wire wire_10617;
    wire wire_10618;
    wire wire_10619;
    wire wire_10620;
    wire wire_10621;
    wire wire_10622;
    wire wire_10623;
    wire wire_10624;
    wire wire_10625;
    wire wire_10626;
    wire wire_10627;
    wire wire_10628;
    wire wire_10629;
    wire wire_10630;
    wire wire_10631;
    wire wire_10632;
    wire wire_10633;
    wire wire_10634;
    wire wire_10635;
    wire wire_10636;
    wire wire_10637;
    wire wire_10638;
    wire wire_10639;
    wire wire_10640;
    wire wire_10641;
    wire wire_10642;
    wire wire_10643;
    wire wire_10644;
    wire wire_10645;
    wire wire_10646;
    wire wire_10647;
    wire wire_10648;
    wire wire_10649;
    wire wire_10650;
    wire wire_10651;
    wire wire_10652;
    wire wire_10653;
    wire wire_10654;
    wire wire_10655;
    wire wire_10656;
    wire wire_10657;
    wire wire_10658;
    wire wire_10659;
    wire wire_10660;
    wire wire_10661;
    wire wire_10662;
    wire wire_10663;
    wire wire_10664;
    wire wire_10665;
    wire wire_10666;
    wire wire_10667;
    wire wire_10668;
    wire wire_10669;
    wire wire_10670;
    wire wire_10671;
    wire wire_10672;
    wire wire_10673;
    wire wire_10674;
    wire wire_10675;
    wire wire_10676;
    wire wire_10677;
    wire wire_10678;
    wire wire_10679;
    wire wire_10680;
    wire wire_10681;
    wire wire_10682;
    wire wire_10683;
    wire wire_10684;
    wire wire_10685;
    wire wire_10686;
    wire wire_10687;
    wire wire_10688;
    wire wire_10689;
    wire wire_10690;
    wire wire_10691;
    wire wire_10692;
    wire wire_10693;
    wire wire_10694;
    wire wire_10695;
    wire wire_10696;
    wire wire_10697;
    wire wire_10698;
    wire wire_10699;
    wire wire_10700;
    wire wire_10701;
    wire wire_10702;
    wire wire_10703;
    wire wire_10704;
    wire wire_10705;
    wire wire_10706;
    wire wire_10707;
    wire wire_10708;
    wire wire_10709;
    wire wire_10710;
    wire wire_10711;
    wire wire_10712;
    wire wire_10713;
    wire wire_10714;
    wire wire_10715;
    wire wire_10716;
    wire wire_10717;
    wire wire_10718;
    wire wire_10719;
    wire wire_10720;
    wire wire_10721;
    wire wire_10722;
    wire wire_10723;
    wire wire_10724;
    wire wire_10725;
    wire wire_10726;
    wire wire_10727;
    wire wire_10728;
    wire wire_10729;
    wire wire_10730;
    wire wire_10731;
    wire wire_10732;
    wire wire_10733;
    wire wire_10734;
    wire wire_10735;
    wire wire_10736;
    wire wire_10737;
    wire wire_10738;
    wire wire_10739;
    wire wire_10740;
    wire wire_10741;
    wire wire_10742;
    wire wire_10743;
    wire wire_10744;
    wire wire_10745;
    wire wire_10746;
    wire wire_10747;
    wire wire_10748;
    wire wire_10749;
    wire wire_10750;
    wire wire_10751;
    wire wire_10752;
    wire wire_10753;
    wire wire_10754;
    wire wire_10755;
    wire wire_10756;
    wire wire_10757;
    wire wire_10758;
    wire wire_10759;
    wire wire_10760;
    wire wire_10761;
    wire wire_10762;
    wire wire_10763;
    wire wire_10764;
    wire wire_10765;
    wire wire_10766;
    wire wire_10767;
    wire wire_10768;
    wire wire_10769;
    wire wire_10770;
    wire wire_10771;
    wire wire_10772;
    wire wire_10773;
    wire wire_10774;
    wire wire_10775;
    wire wire_10776;
    wire wire_10777;
    wire wire_10778;
    wire wire_10779;
    wire wire_10780;
    wire wire_10781;
    wire wire_10782;
    wire wire_10783;
    wire wire_10784;
    wire wire_10785;
    wire wire_10786;
    wire wire_10787;
    wire wire_10788;
    wire wire_10789;
    wire wire_10790;
    wire wire_10791;
    wire wire_10792;
    wire wire_10793;
    wire wire_10794;
    wire wire_10795;
    wire wire_10796;
    wire wire_10797;
    wire wire_10798;
    wire wire_10799;
    wire wire_10800;
    wire wire_10801;
    wire wire_10802;
    wire wire_10803;
    wire wire_10804;
    wire wire_10805;
    wire wire_10806;
    wire wire_10807;
    wire wire_10808;
    wire wire_10809;
    wire wire_10810;
    wire wire_10811;
    wire wire_10812;
    wire wire_10813;
    wire wire_10814;
    wire wire_10815;
    wire wire_10816;
    wire wire_10817;
    wire wire_10818;
    wire wire_10819;
    wire wire_10820;
    wire wire_10821;
    wire wire_10822;
    wire wire_10823;
    wire wire_10824;
    wire wire_10825;
    wire wire_10826;
    wire wire_10827;
    wire wire_10828;
    wire wire_10829;
    wire wire_10830;
    wire wire_10831;
    wire wire_10832;
    wire wire_10833;
    wire wire_10834;
    wire wire_10835;
    wire wire_10836;
    wire wire_10837;
    wire wire_10838;
    wire wire_10839;
    wire wire_10840;
    wire wire_10841;
    wire wire_10842;
    wire wire_10843;
    wire wire_10844;
    wire wire_10845;
    wire wire_10846;
    wire wire_10847;
    wire wire_10848;
    wire wire_10849;
    wire wire_10850;
    wire wire_10851;
    wire wire_10852;
    wire wire_10853;
    wire wire_10854;
    wire wire_10855;
    wire wire_10856;
    wire wire_10857;
    wire wire_10858;
    wire wire_10859;
    wire wire_10860;
    wire wire_10861;
    wire wire_10862;
    wire wire_10863;
    wire wire_10864;
    wire wire_10865;
    wire wire_10866;
    wire wire_10867;
    wire wire_10868;
    wire wire_10869;
    wire wire_10870;
    wire wire_10871;
    wire wire_10872;
    wire wire_10873;
    wire wire_10874;
    wire wire_10875;
    wire wire_10876;
    wire wire_10877;
    wire wire_10878;
    wire wire_10879;
    wire wire_10880;
    wire wire_10881;
    wire wire_10882;
    wire wire_10883;
    wire wire_10884;
    wire wire_10885;
    wire wire_10886;
    wire wire_10887;
    wire wire_10888;
    wire wire_10889;
    wire wire_10890;
    wire wire_10891;
    wire wire_10892;
    wire wire_10893;
    wire wire_10894;
    wire wire_10895;
    wire wire_10896;
    wire wire_10897;
    wire wire_10898;
    wire wire_10899;
    wire wire_10900;
    wire wire_10901;
    wire wire_10902;
    wire wire_10903;
    wire wire_10904;
    wire wire_10905;
    wire wire_10906;
    wire wire_10907;
    wire wire_10908;
    wire wire_10909;
    wire wire_10910;
    wire wire_10911;
    wire wire_10912;
    wire wire_10913;
    wire wire_10914;
    wire wire_10915;
    wire wire_10916;
    wire wire_10917;
    wire wire_10918;
    wire wire_10919;
    wire wire_10920;
    wire wire_10921;
    wire wire_10922;
    wire wire_10923;
    wire wire_10924;
    wire wire_10925;
    wire wire_10926;
    wire wire_10927;
    wire wire_10928;
    wire wire_10929;
    wire wire_10930;
    wire wire_10931;
    wire wire_10932;
    wire wire_10933;
    wire wire_10934;
    wire wire_10935;
    wire wire_10936;
    wire wire_10937;
    wire wire_10938;
    wire wire_10939;
    wire wire_10940;
    wire wire_10941;
    wire wire_10942;
    wire wire_10943;
    wire wire_10944;
    wire wire_10945;
    wire wire_10946;
    wire wire_10947;
    wire wire_10948;
    wire wire_10949;
    wire wire_10950;
    wire wire_10951;
    wire wire_10952;
    wire wire_10953;
    wire wire_10954;
    wire wire_10955;
    wire wire_10956;
    wire wire_10957;
    wire wire_10958;
    wire wire_10959;
    wire wire_10960;
    wire wire_10961;
    wire wire_10962;
    wire wire_10963;
    wire wire_10964;
    wire wire_10965;
    wire wire_10966;
    wire wire_10967;
    wire wire_10968;
    wire wire_10969;
    wire wire_10970;
    wire wire_10971;
    wire wire_10972;
    wire wire_10973;
    wire wire_10974;
    wire wire_10975;
    wire wire_10976;
    wire wire_10977;
    wire wire_10978;
    wire wire_10979;
    wire wire_10980;
    wire wire_10981;
    wire wire_10982;
    wire wire_10983;
    wire wire_10984;
    wire wire_10985;
    wire wire_10986;
    wire wire_10987;
    wire wire_10988;
    wire wire_10989;
    wire wire_10990;
    wire wire_10991;
    wire wire_10992;
    wire wire_10993;
    wire wire_10994;
    wire wire_10995;
    wire wire_10996;
    wire wire_10997;
    wire wire_10998;
    wire wire_10999;
    wire wire_11000;
    wire wire_11001;
    wire wire_11002;
    wire wire_11003;
    wire wire_11004;
    wire wire_11005;
    wire wire_11006;
    wire wire_11007;
    wire wire_11008;
    wire wire_11009;
    wire wire_11010;
    wire wire_11011;
    wire wire_11012;
    wire wire_11013;
    wire wire_11014;
    wire wire_11015;
    wire wire_11016;
    wire wire_11017;
    wire wire_11018;
    wire wire_11019;
    wire wire_11020;
    wire wire_11021;
    wire wire_11022;
    wire wire_11023;
    wire wire_11024;
    wire wire_11025;
    wire wire_11026;
    wire wire_11027;
    wire wire_11028;
    wire wire_11029;
    wire wire_11030;
    wire wire_11031;
    wire wire_11032;
    wire wire_11033;
    wire wire_11034;
    wire wire_11035;
    wire wire_11036;
    wire wire_11037;
    wire wire_11038;
    wire wire_11039;
    wire wire_11040;
    wire wire_11041;
    wire wire_11042;
    wire wire_11043;
    wire wire_11044;
    wire wire_11045;
    wire wire_11046;
    wire wire_11047;
    wire wire_11048;
    wire wire_11049;
    wire wire_11050;
    wire wire_11051;
    wire wire_11052;
    wire wire_11053;
    wire wire_11054;
    wire wire_11055;
    wire wire_11056;
    wire wire_11057;
    wire wire_11058;
    wire wire_11059;
    wire wire_11060;
    wire wire_11061;
    wire wire_11062;
    wire wire_11063;
    wire wire_11064;
    wire wire_11065;
    wire wire_11066;
    wire wire_11067;
    wire wire_11068;
    wire wire_11069;
    wire wire_11070;
    wire wire_11071;
    wire wire_11072;
    wire wire_11073;
    wire wire_11074;
    wire wire_11075;
    wire wire_11076;
    wire wire_11077;
    wire wire_11078;
    wire wire_11079;
    wire wire_11080;
    wire wire_11081;
    wire wire_11082;
    wire wire_11083;
    wire wire_11084;
    wire wire_11085;
    wire wire_11086;
    wire wire_11087;
    wire wire_11088;
    wire wire_11089;
    wire wire_11090;
    wire wire_11091;
    wire wire_11092;
    wire wire_11093;
    wire wire_11094;
    wire wire_11095;
    wire wire_11096;
    wire wire_11097;
    wire wire_11098;
    wire wire_11099;
    wire wire_11100;
    wire wire_11101;
    wire wire_11102;
    wire wire_11103;
    wire wire_11104;
    wire wire_11105;
    wire wire_11106;
    wire wire_11107;
    wire wire_11108;
    wire wire_11109;
    wire wire_11110;
    wire wire_11111;
    wire wire_11112;
    wire wire_11113;
    wire wire_11114;
    wire wire_11115;
    wire wire_11116;
    wire wire_11117;
    wire wire_11118;
    wire wire_11119;
    wire wire_11120;
    wire wire_11121;
    wire wire_11122;
    wire wire_11123;
    wire wire_11124;
    wire wire_11125;
    wire wire_11126;
    wire wire_11127;
    wire wire_11128;
    wire wire_11129;
    wire wire_11130;
    wire wire_11131;
    wire wire_11132;
    wire wire_11133;
    wire wire_11134;
    wire wire_11135;
    wire wire_11136;
    wire wire_11137;
    wire wire_11138;
    wire wire_11139;
    wire wire_11140;
    wire wire_11141;
    wire wire_11142;
    wire wire_11143;
    wire wire_11144;
    wire wire_11145;
    wire wire_11146;
    wire wire_11147;
    wire wire_11148;
    wire wire_11149;
    wire wire_11150;
    wire wire_11151;
    wire wire_11152;
    wire wire_11153;
    wire wire_11154;
    wire wire_11155;
    wire wire_11156;
    wire wire_11157;
    wire wire_11158;
    wire wire_11159;
    wire wire_11160;
    wire wire_11161;
    wire wire_11162;
    wire wire_11163;
    wire wire_11164;
    wire wire_11165;
    wire wire_11166;
    wire wire_11167;
    wire wire_11168;
    wire wire_11169;
    wire wire_11170;
    wire wire_11171;
    wire wire_11172;
    wire wire_11173;
    wire wire_11174;
    wire wire_11175;
    wire wire_11176;
    wire wire_11177;
    wire wire_11178;
    wire wire_11179;
    wire wire_11180;
    wire wire_11181;
    wire wire_11182;
    wire wire_11183;
    wire wire_11184;
    wire wire_11185;
    wire wire_11186;
    wire wire_11187;
    wire wire_11188;
    wire wire_11189;
    wire wire_11190;
    wire wire_11191;
    wire wire_11192;
    wire wire_11193;
    wire wire_11194;
    wire wire_11195;
    wire wire_11196;
    wire wire_11197;
    wire wire_11198;
    wire wire_11199;
    wire wire_11200;
    wire wire_11201;
    wire wire_11202;
    wire wire_11203;
    wire wire_11204;
    wire wire_11205;
    wire wire_11206;
    wire wire_11207;
    wire wire_11208;
    wire wire_11209;
    wire wire_11210;
    wire wire_11211;
    wire wire_11212;
    wire wire_11213;
    wire wire_11214;
    wire wire_11215;
    wire wire_11216;
    wire wire_11217;
    wire wire_11218;
    wire wire_11219;
    wire wire_11220;
    wire wire_11221;
    wire wire_11222;
    wire wire_11223;
    wire wire_11224;
    wire wire_11225;
    wire wire_11226;
    wire wire_11227;
    wire wire_11228;
    wire wire_11229;
    wire wire_11230;
    wire wire_11231;
    wire wire_11232;
    wire wire_11233;
    wire wire_11234;
    wire wire_11235;
    wire wire_11236;
    wire wire_11237;
    wire wire_11238;
    wire wire_11239;
    wire wire_11240;
    wire wire_11241;
    wire wire_11242;
    wire wire_11243;
    wire wire_11244;
    wire wire_11245;
    wire wire_11246;
    wire wire_11247;
    wire wire_11248;
    wire wire_11249;
    wire wire_11250;
    wire wire_11251;
    wire wire_11252;
    wire wire_11253;
    wire wire_11254;
    wire wire_11255;
    wire wire_11256;
    wire wire_11257;
    wire wire_11258;
    wire wire_11259;
    wire wire_11260;
    wire wire_11261;
    wire wire_11262;
    wire wire_11263;
    wire wire_11264;
    wire wire_11265;
    wire wire_11266;
    wire wire_11267;
    wire wire_11268;
    wire wire_11269;
    wire wire_11270;
    wire wire_11271;
    wire wire_11272;
    wire wire_11273;
    wire wire_11274;
    wire wire_11275;
    wire wire_11276;
    wire wire_11277;
    wire wire_11278;
    wire wire_11279;
    wire wire_11280;
    wire wire_11281;
    wire wire_11282;
    wire wire_11283;
    wire wire_11284;
    wire wire_11285;
    wire wire_11286;
    wire wire_11287;
    wire wire_11288;
    wire wire_11289;
    wire wire_11290;
    wire wire_11291;
    wire wire_11292;
    wire wire_11293;
    wire wire_11294;
    wire wire_11295;
    wire wire_11296;
    wire wire_11297;
    wire wire_11298;
    wire wire_11299;
    wire wire_11300;
    wire wire_11301;
    wire wire_11302;
    wire wire_11303;
    wire wire_11304;
    wire wire_11305;
    wire wire_11306;
    wire wire_11307;
    wire wire_11308;
    wire wire_11309;
    wire wire_11310;
    wire wire_11311;
    wire wire_11312;
    wire wire_11313;
    wire wire_11314;
    wire wire_11315;
    wire wire_11316;
    wire wire_11317;
    wire wire_11318;
    wire wire_11319;
    wire wire_11320;
    wire wire_11321;
    wire wire_11322;
    wire wire_11323;
    wire wire_11324;
    wire wire_11325;
    wire wire_11326;
    wire wire_11327;
    wire wire_11328;
    wire wire_11329;
    wire wire_11330;
    wire wire_11331;
    wire wire_11332;
    wire wire_11333;
    wire wire_11334;
    wire wire_11335;
    wire wire_11336;
    wire wire_11337;
    wire wire_11338;
    wire wire_11339;
    wire wire_11340;
    wire wire_11341;
    wire wire_11342;
    wire wire_11343;
    wire wire_11344;
    wire wire_11345;
    wire wire_11346;
    wire wire_11347;
    wire wire_11348;
    wire wire_11349;
    wire wire_11350;
    wire wire_11351;
    wire wire_11352;
    wire wire_11353;
    wire wire_11354;
    wire wire_11355;
    wire wire_11356;
    wire wire_11357;
    wire wire_11358;
    wire wire_11359;
    wire wire_11360;
    wire wire_11361;
    wire wire_11362;
    wire wire_11363;
    wire wire_11364;
    wire wire_11365;
    wire wire_11366;
    wire wire_11367;
    wire wire_11368;
    wire wire_11369;
    wire wire_11370;
    wire wire_11371;
    wire wire_11372;
    wire wire_11373;
    wire wire_11374;
    wire wire_11375;
    wire wire_11376;
    wire wire_11377;
    wire wire_11378;
    wire wire_11379;
    wire wire_11380;
    wire wire_11381;
    wire wire_11382;
    wire wire_11383;
    wire wire_11384;
    wire wire_11385;
    wire wire_11386;
    wire wire_11387;
    wire wire_11388;
    wire wire_11389;
    wire wire_11390;
    wire wire_11391;
    wire wire_11392;
    wire wire_11393;
    wire wire_11394;
    wire wire_11395;
    wire wire_11396;
    wire wire_11397;
    wire wire_11398;
    wire wire_11399;
    wire wire_11400;
    wire wire_11401;
    wire wire_11402;
    wire wire_11403;
    wire wire_11404;
    wire wire_11405;
    wire wire_11406;
    wire wire_11407;
    wire wire_11408;
    wire wire_11409;
    wire wire_11410;
    wire wire_11411;
    wire wire_11412;
    wire wire_11413;
    wire wire_11414;
    wire wire_11415;
    wire wire_11416;
    wire wire_11417;
    wire wire_11418;
    wire wire_11419;
    wire wire_11420;
    wire wire_11421;
    wire wire_11422;
    wire wire_11423;
    wire wire_11424;
    wire wire_11425;
    wire wire_11426;
    wire wire_11427;
    wire wire_11428;
    wire wire_11429;
    wire wire_11430;
    wire wire_11431;
    wire wire_11432;
    wire wire_11433;
    wire wire_11434;
    wire wire_11435;
    wire wire_11436;
    wire wire_11437;
    wire wire_11438;
    wire wire_11439;
    wire wire_11440;
    wire wire_11441;
    wire wire_11442;
    wire wire_11443;
    wire wire_11444;
    wire wire_11445;
    wire wire_11446;
    wire wire_11447;
    wire wire_11448;
    wire wire_11449;
    wire wire_11450;
    wire wire_11451;
    wire wire_11452;
    wire wire_11453;
    wire wire_11454;
    wire wire_11455;
    wire wire_11456;
    wire wire_11457;
    wire wire_11458;
    wire wire_11459;
    wire wire_11460;
    wire wire_11461;
    wire wire_11462;
    wire wire_11463;
    wire wire_11464;
    wire wire_11465;
    wire wire_11466;
    wire wire_11467;
    wire wire_11468;
    wire wire_11469;
    wire wire_11470;
    wire wire_11471;
    wire wire_11472;
    wire wire_11473;
    wire wire_11474;
    wire wire_11475;
    wire wire_11476;
    wire wire_11477;
    wire wire_11478;
    wire wire_11479;
    wire wire_11480;
    wire wire_11481;
    wire wire_11482;
    wire wire_11483;
    wire wire_11484;
    wire wire_11485;
    wire wire_11486;
    wire wire_11487;
    wire wire_11488;
    wire wire_11489;
    wire wire_11490;
    wire wire_11491;
    wire wire_11492;
    wire wire_11493;
    wire wire_11494;
    wire wire_11495;
    wire wire_11496;
    wire wire_11497;
    wire wire_11498;
    wire wire_11499;
    wire wire_11500;
    wire wire_11501;
    wire wire_11502;
    wire wire_11503;
    wire wire_11504;
    wire wire_11505;
    wire wire_11506;
    wire wire_11507;
    wire wire_11508;
    wire wire_11509;
    wire wire_11510;
    wire wire_11511;
    wire wire_11512;
    wire wire_11513;
    wire wire_11514;
    wire wire_11515;
    wire wire_11516;
    wire wire_11517;
    wire wire_11518;
    wire wire_11519;
    wire wire_11520;
    wire wire_11521;
    wire wire_11522;
    wire wire_11523;
    wire wire_11524;
    wire wire_11525;
    wire wire_11526;
    wire wire_11527;
    wire wire_11528;
    wire wire_11529;
    wire wire_11530;
    wire wire_11531;
    wire wire_11532;
    wire wire_11533;
    wire wire_11534;
    wire wire_11535;
    wire wire_11536;
    wire wire_11537;
    wire wire_11538;
    wire wire_11539;
    wire wire_11540;
    wire wire_11541;
    wire wire_11542;
    wire wire_11543;
    wire wire_11544;
    wire wire_11545;
    wire wire_11546;
    wire wire_11547;
    wire wire_11548;
    wire wire_11549;
    wire wire_11550;
    wire wire_11551;
    wire wire_11552;
    wire wire_11553;
    wire wire_11554;
    wire wire_11555;
    wire wire_11556;
    wire wire_11557;
    wire wire_11558;
    wire wire_11559;
    wire wire_11560;
    wire wire_11561;
    wire wire_11562;
    wire wire_11563;
    wire wire_11564;
    wire wire_11565;
    wire wire_11566;
    wire wire_11567;
    wire wire_11568;
    wire wire_11569;
    wire wire_11570;
    wire wire_11571;
    wire wire_11572;
    wire wire_11573;
    wire wire_11574;
    wire wire_11575;
    wire wire_11576;
    wire wire_11577;
    wire wire_11578;
    wire wire_11579;
    wire wire_11580;
    wire wire_11581;
    wire wire_11582;
    wire wire_11583;
    wire wire_11584;
    wire wire_11585;
    wire wire_11586;
    wire wire_11587;
    wire wire_11588;
    wire wire_11589;
    wire wire_11590;
    wire wire_11591;
    wire wire_11592;
    wire wire_11593;
    wire wire_11594;
    wire wire_11595;
    wire wire_11596;
    wire wire_11597;
    wire wire_11598;
    wire wire_11599;
    wire wire_11600;
    wire wire_11601;
    wire wire_11602;
    wire wire_11603;
    wire wire_11604;
    wire wire_11605;
    wire wire_11606;
    wire wire_11607;
    wire wire_11608;
    wire wire_11609;
    wire wire_11610;
    wire wire_11611;
    wire wire_11612;
    wire wire_11613;
    wire wire_11614;
    wire wire_11615;
    wire wire_11616;
    wire wire_11617;
    wire wire_11618;
    wire wire_11619;
    wire wire_11620;
    wire wire_11621;
    wire wire_11622;
    wire wire_11623;
    wire wire_11624;
    wire wire_11625;
    wire wire_11626;
    wire wire_11627;
    wire wire_11628;
    wire wire_11629;
    wire wire_11630;
    wire wire_11631;
    wire wire_11632;
    wire wire_11633;
    wire wire_11634;
    wire wire_11635;
    wire wire_11636;
    wire wire_11637;
    wire wire_11638;
    wire wire_11639;
    wire wire_11640;
    wire wire_11641;
    wire wire_11642;
    wire wire_11643;
    wire wire_11644;
    wire wire_11645;
    wire wire_11646;
    wire wire_11647;
    wire wire_11648;
    wire wire_11649;
    wire wire_11650;
    wire wire_11651;
    wire wire_11652;
    wire wire_11653;
    wire wire_11654;
    wire wire_11655;
    wire wire_11656;
    wire wire_11657;
    wire wire_11658;
    wire wire_11659;
    wire wire_11660;
    wire wire_11661;
    wire wire_11662;
    wire wire_11663;
    wire wire_11664;
    wire wire_11665;
    wire wire_11666;
    wire wire_11667;
    wire wire_11668;
    wire wire_11669;
    wire wire_11670;
    wire wire_11671;
    wire wire_11672;
    wire wire_11673;
    wire wire_11674;
    wire wire_11675;
    wire wire_11676;
    wire wire_11677;
    wire wire_11678;
    wire wire_11679;
    wire wire_11680;
    wire wire_11681;
    wire wire_11682;
    wire wire_11683;
    wire wire_11684;
    wire wire_11685;
    wire wire_11686;
    wire wire_11687;
    wire wire_11688;
    wire wire_11689;
    wire wire_11690;
    wire wire_11691;
    wire wire_11692;
    wire wire_11693;
    wire wire_11694;
    wire wire_11695;
    wire wire_11696;
    wire wire_11697;
    wire wire_11698;
    wire wire_11699;
    wire wire_11700;
    wire wire_11701;
    wire wire_11702;
    wire wire_11703;
    wire wire_11704;
    wire wire_11705;
    wire wire_11706;
    wire wire_11707;
    wire wire_11708;
    wire wire_11709;
    wire wire_11710;
    wire wire_11711;
    wire wire_11712;
    wire wire_11713;
    wire wire_11714;
    wire wire_11715;
    wire wire_11716;
    wire wire_11717;
    wire wire_11718;
    wire wire_11719;
    wire wire_11720;
    wire wire_11721;
    wire wire_11722;
    wire wire_11723;
    wire wire_11724;
    wire wire_11725;
    wire wire_11726;
    wire wire_11727;
    wire wire_11728;
    wire wire_11729;
    wire wire_11730;
    wire wire_11731;
    wire wire_11732;
    wire wire_11733;
    wire wire_11734;
    wire wire_11735;
    wire wire_11736;
    wire wire_11737;
    wire wire_11738;
    wire wire_11739;
    wire wire_11740;
    wire wire_11741;
    wire wire_11742;
    wire wire_11743;
    wire wire_11744;
    wire wire_11745;
    wire wire_11746;
    wire wire_11747;
    wire wire_11748;
    wire wire_11749;
    wire wire_11750;
    wire wire_11751;
    wire wire_11752;
    wire wire_11753;
    wire wire_11754;
    wire wire_11755;
    wire wire_11756;
    wire wire_11757;
    wire wire_11758;
    wire wire_11759;
    wire wire_11760;
    wire wire_11761;
    wire wire_11762;
    wire wire_11763;
    wire wire_11764;
    wire wire_11765;
    wire wire_11766;
    wire wire_11767;
    wire wire_11768;
    wire wire_11769;
    wire wire_11770;
    wire wire_11771;
    wire wire_11772;
    wire wire_11773;
    wire wire_11774;
    wire wire_11775;
    wire wire_11776;
    wire wire_11777;
    wire wire_11778;
    wire wire_11779;
    wire wire_11780;
    wire wire_11781;
    wire wire_11782;
    wire wire_11783;
    wire wire_11784;
    wire wire_11785;
    wire wire_11786;
    wire wire_11787;
    wire wire_11788;
    wire wire_11789;
    wire wire_11790;
    wire wire_11791;
    wire wire_11792;
    wire wire_11793;
    wire wire_11794;
    wire wire_11795;
    wire wire_11796;
    wire wire_11797;
    wire wire_11798;
    wire wire_11799;
    wire wire_11800;
    wire wire_11801;
    wire wire_11802;
    wire wire_11803;
    wire wire_11804;
    wire wire_11805;
    wire wire_11806;
    wire wire_11807;
    wire wire_11808;
    wire wire_11809;
    wire wire_11810;
    wire wire_11811;
    wire wire_11812;
    wire wire_11813;
    wire wire_11814;
    wire wire_11815;
    wire wire_11816;
    wire wire_11817;
    wire wire_11818;
    wire wire_11819;
    wire wire_11820;
    wire wire_11821;
    wire wire_11822;
    wire wire_11823;
    wire wire_11824;
    wire wire_11825;
    wire wire_11826;
    wire wire_11827;
    wire wire_11828;
    wire wire_11829;
    wire wire_11830;
    wire wire_11831;
    wire wire_11832;
    wire wire_11833;
    wire wire_11834;
    wire wire_11835;
    wire wire_11836;
    wire wire_11837;
    wire wire_11838;
    wire wire_11839;
    wire wire_11840;
    wire wire_11841;
    wire wire_11842;
    wire wire_11843;
    wire wire_11844;
    wire wire_11845;
    wire wire_11846;
    wire wire_11847;
    wire wire_11848;
    wire wire_11849;
    wire wire_11850;
    wire wire_11851;
    wire wire_11852;
    wire wire_11853;
    wire wire_11854;
    wire wire_11855;
    wire wire_11856;
    wire wire_11857;
    wire wire_11858;
    wire wire_11859;
    wire wire_11860;
    wire wire_11861;
    wire wire_11862;
    wire wire_11863;
    wire wire_11864;
    wire wire_11865;
    wire wire_11866;
    wire wire_11867;
    wire wire_11868;
    wire wire_11869;
    wire wire_11870;
    wire wire_11871;
    wire wire_11872;
    wire wire_11873;
    wire wire_11874;
    wire wire_11875;
    wire wire_11876;
    wire wire_11877;
    wire wire_11878;
    wire wire_11879;
    wire wire_11880;
    wire wire_11881;
    wire wire_11882;
    wire wire_11883;
    wire wire_11884;
    wire wire_11885;
    wire wire_11886;
    wire wire_11887;
    wire wire_11888;
    wire wire_11889;
    wire wire_11890;
    wire wire_11891;
    wire wire_11892;
    wire wire_11893;
    wire wire_11894;
    wire wire_11895;
    wire wire_11896;
    wire wire_11897;
    wire wire_11898;
    wire wire_11899;
    wire wire_11900;
    wire wire_11901;
    wire wire_11902;
    wire wire_11903;
    wire wire_11904;
    wire wire_11905;
    wire wire_11906;
    wire wire_11907;
    wire wire_11908;
    wire wire_11909;
    wire wire_11910;
    wire wire_11911;
    wire wire_11912;
    wire wire_11913;
    wire wire_11914;
    wire wire_11915;
    wire wire_11916;
    wire wire_11917;
    wire wire_11918;
    wire wire_11919;
    wire wire_11920;
    wire wire_11921;
    wire wire_11922;
    wire wire_11923;
    wire wire_11924;
    wire wire_11925;
    wire wire_11926;
    wire wire_11927;
    wire wire_11928;
    wire wire_11929;
    wire wire_11930;
    wire wire_11931;
    wire wire_11932;
    wire wire_11933;
    wire wire_11934;
    wire wire_11935;
    wire wire_11936;
    wire wire_11937;
    wire wire_11938;
    wire wire_11939;
    wire wire_11940;
    wire wire_11941;
    wire wire_11942;
    wire wire_11943;
    wire wire_11944;
    wire wire_11945;
    wire wire_11946;
    wire wire_11947;
    wire wire_11948;
    wire wire_11949;
    wire wire_11950;
    wire wire_11951;
    wire wire_11952;
    wire wire_11953;
    wire wire_11954;
    wire wire_11955;
    wire wire_11956;
    wire wire_11957;
    wire wire_11958;
    wire wire_11959;
    wire wire_11960;
    wire wire_11961;
    wire wire_11962;
    wire wire_11963;
    wire wire_11964;
    wire wire_11965;
    wire wire_11966;
    wire wire_11967;
    wire wire_11968;
    wire wire_11969;
    wire wire_11970;
    wire wire_11971;
    wire wire_11972;
    wire wire_11973;
    wire wire_11974;
    wire wire_11975;
    wire wire_11976;
    wire wire_11977;
    wire wire_11978;
    wire wire_11979;
    wire wire_11980;
    wire wire_11981;
    wire wire_11982;
    wire wire_11983;
    wire wire_11984;
    wire wire_11985;
    wire wire_11986;
    wire wire_11987;
    wire wire_11988;
    wire wire_11989;
    wire wire_11990;
    wire wire_11991;
    wire wire_11992;
    wire wire_11993;
    wire wire_11994;
    wire wire_11995;
    wire wire_11996;
    wire wire_11997;
    wire wire_11998;
    wire wire_11999;
    wire wire_12000;
    wire wire_12001;
    wire wire_12002;
    wire wire_12003;
    wire wire_12004;
    wire wire_12005;
    wire wire_12006;
    wire wire_12007;
    wire wire_12008;
    wire wire_12009;
    wire wire_12010;
    wire wire_12011;
    wire wire_12012;
    wire wire_12013;
    wire wire_12014;
    wire wire_12015;
    wire wire_12016;
    wire wire_12017;
    wire wire_12018;
    wire wire_12019;
    wire wire_12020;
    wire wire_12021;
    wire wire_12022;
    wire wire_12023;
    wire wire_12024;
    wire wire_12025;
    wire wire_12026;
    wire wire_12027;
    wire wire_12028;
    wire wire_12029;
    wire wire_12030;
    wire wire_12031;
    wire wire_12032;
    wire wire_12033;
    wire wire_12034;
    wire wire_12035;
    wire wire_12036;
    wire wire_12037;
    wire wire_12038;
    wire wire_12039;
    wire wire_12040;
    wire wire_12041;
    wire wire_12042;
    wire wire_12043;
    wire wire_12044;
    wire wire_12045;
    wire wire_12046;
    wire wire_12047;
    wire wire_12048;
    wire wire_12049;
    wire wire_12050;
    wire wire_12051;
    wire wire_12052;
    wire wire_12053;
    wire wire_12054;
    wire wire_12055;
    wire wire_12056;
    wire wire_12057;
    wire wire_12058;
    wire wire_12059;
    wire wire_12060;
    wire wire_12061;
    wire wire_12062;
    wire wire_12063;
    wire wire_12064;
    wire wire_12065;
    wire wire_12066;
    wire wire_12067;
    wire wire_12068;
    wire wire_12069;
    wire wire_12070;
    wire wire_12071;
    wire wire_12072;
    wire wire_12073;
    wire wire_12074;
    wire wire_12075;
    wire wire_12076;
    wire wire_12077;
    wire wire_12078;
    wire wire_12079;
    wire wire_12080;
    wire wire_12081;
    wire wire_12082;
    wire wire_12083;
    wire wire_12084;
    wire wire_12085;
    wire wire_12086;
    wire wire_12087;
    wire wire_12088;
    wire wire_12089;
    wire wire_12090;
    wire wire_12091;
    wire wire_12092;
    wire wire_12093;
    wire wire_12094;
    wire wire_12095;
    wire wire_12096;
    wire wire_12097;
    wire wire_12098;
    wire wire_12099;
    wire wire_12100;
    wire wire_12101;
    wire wire_12102;
    wire wire_12103;
    wire wire_12104;
    wire wire_12105;
    wire wire_12106;
    wire wire_12107;
    wire wire_12108;
    wire wire_12109;
    wire wire_12110;
    wire wire_12111;
    wire wire_12112;
    wire wire_12113;
    wire wire_12114;
    wire wire_12115;
    wire wire_12116;
    wire wire_12117;
    wire wire_12118;
    wire wire_12119;
    wire wire_12120;
    wire wire_12121;
    wire wire_12122;
    wire wire_12123;
    wire wire_12124;
    wire wire_12125;
    wire wire_12126;
    wire wire_12127;
    wire wire_12128;
    wire wire_12129;
    wire wire_12130;
    wire wire_12131;
    wire wire_12132;
    wire wire_12133;
    wire wire_12134;
    wire wire_12135;
    wire wire_12136;
    wire wire_12137;
    wire wire_12138;
    wire wire_12139;
    wire wire_12140;
    wire wire_12141;
    wire wire_12142;
    wire wire_12143;
    wire wire_12144;
    wire wire_12145;
    wire wire_12146;
    wire wire_12147;
    wire wire_12148;
    wire wire_12149;
    wire wire_12150;
    wire wire_12151;
    wire wire_12152;
    wire wire_12153;
    wire wire_12154;
    wire wire_12155;
    wire wire_12156;
    wire wire_12157;
    wire wire_12158;
    wire wire_12159;
    wire wire_12160;
    wire wire_12161;
    wire wire_12162;
    wire wire_12163;
    wire wire_12164;
    wire wire_12165;
    wire wire_12166;
    wire wire_12167;
    wire wire_12168;
    wire wire_12169;
    wire wire_12170;
    wire wire_12171;
    wire wire_12172;
    wire wire_12173;
    wire wire_12174;
    wire wire_12175;
    wire wire_12176;
    wire wire_12177;
    wire wire_12178;
    wire wire_12179;
    wire wire_12180;
    wire wire_12181;
    wire wire_12182;
    wire wire_12183;
    wire wire_12184;
    wire wire_12185;
    wire wire_12186;
    wire wire_12187;
    wire wire_12188;
    wire wire_12189;
    wire wire_12190;
    wire wire_12191;
    wire wire_12192;
    wire wire_12193;
    wire wire_12194;
    wire wire_12195;
    wire wire_12196;
    wire wire_12197;
    wire wire_12198;
    wire wire_12199;
    wire wire_12200;
    wire wire_12201;
    wire wire_12202;
    wire wire_12203;
    wire wire_12204;
    wire wire_12205;
    wire wire_12206;
    wire wire_12207;
    wire wire_12208;
    wire wire_12209;
    wire wire_12210;
    wire wire_12211;
    wire wire_12212;
    wire wire_12213;
    wire wire_12214;
    wire wire_12215;
    wire wire_12216;
    wire wire_12217;
    wire wire_12218;
    wire wire_12219;
    wire wire_12220;
    wire wire_12221;
    wire wire_12222;
    wire wire_12223;
    wire wire_12224;
    wire wire_12225;
    wire wire_12226;
    wire wire_12227;
    wire wire_12228;
    wire wire_12229;
    wire wire_12230;
    wire wire_12231;
    wire wire_12232;
    wire wire_12233;
    wire wire_12234;
    wire wire_12235;
    wire wire_12236;
    wire wire_12237;
    wire wire_12238;
    wire wire_12239;
    wire wire_12240;
    wire wire_12241;
    wire wire_12242;
    wire wire_12243;
    wire wire_12244;
    wire wire_12245;
    wire wire_12246;
    wire wire_12247;
    wire wire_12248;
    wire wire_12249;
    wire wire_12250;
    wire wire_12251;
    wire wire_12252;
    wire wire_12253;
    wire wire_12254;
    wire wire_12255;
    wire wire_12256;
    wire wire_12257;
    wire wire_12258;
    wire wire_12259;
    wire wire_12260;
    wire wire_12261;
    wire wire_12262;
    wire wire_12263;
    wire wire_12264;
    wire wire_12265;
    wire wire_12266;
    wire wire_12267;
    wire wire_12268;
    wire wire_12269;
    wire wire_12270;
    wire wire_12271;
    wire wire_12272;
    wire wire_12273;
    wire wire_12274;
    wire wire_12275;
    wire wire_12276;
    wire wire_12277;
    wire wire_12278;
    wire wire_12279;
    wire wire_12280;
    wire wire_12281;
    wire wire_12282;
    wire wire_12283;
    wire wire_12284;
    wire wire_12285;
    wire wire_12286;
    wire wire_12287;
    wire wire_12288;
    wire wire_12289;
    wire wire_12290;
    wire wire_12291;
    wire wire_12292;
    wire wire_12293;
    wire wire_12294;
    wire wire_12295;
    wire wire_12296;
    wire wire_12297;
    wire wire_12298;
    wire wire_12299;
    wire wire_12300;
    wire wire_12301;
    wire wire_12302;
    wire wire_12303;
    wire wire_12304;
    wire wire_12305;
    wire wire_12306;
    wire wire_12307;
    wire wire_12308;
    wire wire_12309;
    wire wire_12310;
    wire wire_12311;
    wire wire_12312;
    wire wire_12313;
    wire wire_12314;
    wire wire_12315;
    wire wire_12316;
    wire wire_12317;
    wire wire_12318;
    wire wire_12319;
    wire wire_12320;
    wire wire_12321;
    wire wire_12322;
    wire wire_12323;
    wire wire_12324;
    wire wire_12325;
    wire wire_12326;
    wire wire_12327;
    wire wire_12328;
    wire wire_12329;
    wire wire_12330;
    wire wire_12331;
    wire wire_12332;
    wire wire_12333;
    wire wire_12334;
    wire wire_12335;
    wire wire_12336;
    wire wire_12337;
    wire wire_12338;
    wire wire_12339;
    wire wire_12340;
    wire wire_12341;
    wire wire_12342;
    wire wire_12343;
    wire wire_12344;
    wire wire_12345;
    wire wire_12346;
    wire wire_12347;
    wire wire_12348;
    wire wire_12349;
    wire wire_12350;
    wire wire_12351;
    wire wire_12352;
    wire wire_12353;
    wire wire_12354;
    wire wire_12355;
    wire wire_12356;
    wire wire_12357;
    wire wire_12358;
    wire wire_12359;
    wire wire_12360;
    wire wire_12361;
    wire wire_12362;
    wire wire_12363;
    wire wire_12364;
    wire wire_12365;
    wire wire_12366;
    wire wire_12367;
    wire wire_12368;
    wire wire_12369;
    wire wire_12370;
    wire wire_12371;
    wire wire_12372;
    wire wire_12373;
    wire wire_12374;
    wire wire_12375;
    wire wire_12376;
    wire wire_12377;
    wire wire_12378;
    wire wire_12379;
    wire wire_12380;
    wire wire_12381;
    wire wire_12382;
    wire wire_12383;
    wire wire_12384;
    wire wire_12385;
    wire wire_12386;
    wire wire_12387;
    wire wire_12388;
    wire wire_12389;
    wire wire_12390;
    wire wire_12391;
    wire wire_12392;
    wire wire_12393;
    wire wire_12394;
    wire wire_12395;
    wire wire_12396;
    wire wire_12397;
    wire wire_12398;
    wire wire_12399;
    wire wire_12400;
    wire wire_12401;
    wire wire_12402;
    wire wire_12403;
    wire wire_12404;
    wire wire_12405;
    wire wire_12406;
    wire wire_12407;
    wire wire_12408;
    wire wire_12409;
    wire wire_12410;
    wire wire_12411;
    wire wire_12412;
    wire wire_12413;
    wire wire_12414;
    wire wire_12415;
    wire wire_12416;
    wire wire_12417;
    wire wire_12418;
    wire wire_12419;
    wire wire_12420;
    wire wire_12421;
    wire wire_12422;
    wire wire_12423;
    wire wire_12424;
    wire wire_12425;
    wire wire_12426;
    wire wire_12427;
    wire wire_12428;
    wire wire_12429;
    wire wire_12430;
    wire wire_12431;
    wire wire_12432;
    wire wire_12433;
    wire wire_12434;
    wire wire_12435;
    wire wire_12436;
    wire wire_12437;
    wire wire_12438;
    wire wire_12439;
    wire wire_12440;
    wire wire_12441;
    wire wire_12442;
    wire wire_12443;
    wire wire_12444;
    wire wire_12445;
    wire wire_12446;
    wire wire_12447;
    wire wire_12448;
    wire wire_12449;
    wire wire_12450;
    wire wire_12451;
    wire wire_12452;
    wire wire_12453;
    wire wire_12454;
    wire wire_12455;
    wire wire_12456;
    wire wire_12457;
    wire wire_12458;
    wire wire_12459;
    wire wire_12460;
    wire wire_12461;
    wire wire_12462;
    wire wire_12463;
    wire wire_12464;
    wire wire_12465;
    wire wire_12466;
    wire wire_12467;
    wire wire_12468;
    wire wire_12469;
    wire wire_12470;
    wire wire_12471;
    wire wire_12472;
    wire wire_12473;
    wire wire_12474;
    wire wire_12475;
    wire wire_12476;
    wire wire_12477;
    wire wire_12478;
    wire wire_12479;
    wire wire_12480;
    wire wire_12481;
    wire wire_12482;
    wire wire_12483;
    wire wire_12484;
    wire wire_12485;
    wire wire_12486;
    wire wire_12487;
    wire wire_12488;
    wire wire_12489;
    wire wire_12490;
    wire wire_12491;
    wire wire_12492;
    wire wire_12493;
    wire wire_12494;
    wire wire_12495;
    wire wire_12496;
    wire wire_12497;
    wire wire_12498;
    wire wire_12499;
    wire wire_12500;
    wire wire_12501;
    wire wire_12502;
    wire wire_12503;
    wire wire_12504;
    wire wire_12505;
    wire wire_12506;
    wire wire_12507;
    wire wire_12508;
    wire wire_12509;
    wire wire_12510;
    wire wire_12511;
    wire wire_12512;
    wire wire_12513;
    wire wire_12514;
    wire wire_12515;
    wire wire_12516;
    wire wire_12517;
    wire wire_12518;
    wire wire_12519;
    wire wire_12520;
    wire wire_12521;
    wire wire_12522;
    wire wire_12523;
    wire wire_12524;
    wire wire_12525;
    wire wire_12526;
    wire wire_12527;
    wire wire_12528;
    wire wire_12529;
    wire wire_12530;
    wire wire_12531;
    wire wire_12532;
    wire wire_12533;
    wire wire_12534;
    wire wire_12535;
    wire wire_12536;
    wire wire_12537;
    wire wire_12538;
    wire wire_12539;
    wire wire_12540;
    wire wire_12541;
    wire wire_12542;
    wire wire_12543;
    wire wire_12544;
    wire wire_12545;
    wire wire_12546;
    wire wire_12547;
    wire wire_12548;
    wire wire_12549;
    wire wire_12550;
    wire wire_12551;
    wire wire_12552;
    wire wire_12553;
    wire wire_12554;
    wire wire_12555;
    wire wire_12556;
    wire wire_12557;
    wire wire_12558;
    wire wire_12559;
    wire wire_12560;
    wire wire_12561;
    wire wire_12562;
    wire wire_12563;
    wire wire_12564;
    wire wire_12565;
    wire wire_12566;
    wire wire_12567;
    wire wire_12568;
    wire wire_12569;
    wire wire_12570;
    wire wire_12571;
    wire wire_12572;
    wire wire_12573;
    wire wire_12574;
    wire wire_12575;
    wire wire_12576;
    wire wire_12577;
    wire wire_12578;
    wire wire_12579;
    wire wire_12580;
    wire wire_12581;
    wire wire_12582;
    wire wire_12583;
    wire wire_12584;
    wire wire_12585;
    wire wire_12586;
    wire wire_12587;
    wire wire_12588;
    wire wire_12589;
    wire wire_12590;
    wire wire_12591;
    wire wire_12592;
    wire wire_12593;
    wire wire_12594;
    wire wire_12595;
    wire wire_12596;
    wire wire_12597;
    wire wire_12598;
    wire wire_12599;
    wire wire_12600;
    wire wire_12601;
    wire wire_12602;
    wire wire_12603;
    wire wire_12604;
    wire wire_12605;
    wire wire_12606;
    wire wire_12607;
    wire wire_12608;
    wire wire_12609;
    wire wire_12610;
    wire wire_12611;
    wire wire_12612;
    wire wire_12613;
    wire wire_12614;
    wire wire_12615;
    wire wire_12616;
    wire wire_12617;
    wire wire_12618;
    wire wire_12619;
    wire wire_12620;
    wire wire_12621;
    wire wire_12622;
    wire wire_12623;
    wire wire_12624;
    wire wire_12625;
    wire wire_12626;
    wire wire_12627;
    wire wire_12628;
    wire wire_12629;
    wire wire_12630;
    wire wire_12631;
    wire wire_12632;
    wire wire_12633;
    wire wire_12634;
    wire wire_12635;
    wire wire_12636;
    wire wire_12637;
    wire wire_12638;
    wire wire_12639;
    wire wire_12640;
    wire wire_12641;
    wire wire_12642;
    wire wire_12643;
    wire wire_12644;
    wire wire_12645;
    wire wire_12646;
    wire wire_12647;
    wire wire_12648;
    wire wire_12649;
    wire wire_12650;
    wire wire_12651;
    wire wire_12652;
    wire wire_12653;
    wire wire_12654;
    wire wire_12655;
    wire wire_12656;
    wire wire_12657;
    wire wire_12658;
    wire wire_12659;
    wire wire_12660;
    wire wire_12661;
    wire wire_12662;
    wire wire_12663;
    wire wire_12664;
    wire wire_12665;
    wire wire_12666;
    wire wire_12667;
    wire wire_12668;
    wire wire_12669;
    wire wire_12670;
    wire wire_12671;
    wire wire_12672;
    wire wire_12673;
    wire wire_12674;
    wire wire_12675;
    wire wire_12676;
    wire wire_12677;
    wire wire_12678;
    wire wire_12679;
    wire wire_12680;
    wire wire_12681;
    wire wire_12682;
    wire wire_12683;
    wire wire_12684;
    wire wire_12685;
    wire wire_12686;
    wire wire_12687;
    wire wire_12688;
    wire wire_12689;
    wire wire_12690;
    wire wire_12691;
    wire wire_12692;
    wire wire_12693;
    wire wire_12694;
    wire wire_12695;
    wire wire_12696;
    wire wire_12697;
    wire wire_12698;
    wire wire_12699;
    wire wire_12700;
    wire wire_12701;
    wire wire_12702;
    wire wire_12703;
    wire wire_12704;
    wire wire_12705;
    wire wire_12706;
    wire wire_12707;
    wire wire_12708;
    wire wire_12709;
    wire wire_12710;
    wire wire_12711;
    wire wire_12712;
    wire wire_12713;
    wire wire_12714;
    wire wire_12715;
    wire wire_12716;
    wire wire_12717;
    wire wire_12718;
    wire wire_12719;
    wire wire_12720;
    wire wire_12721;
    wire wire_12722;
    wire wire_12723;
    wire wire_12724;
    wire wire_12725;
    wire wire_12726;
    wire wire_12727;
    wire wire_12728;
    wire wire_12729;
    wire wire_12730;
    wire wire_12731;
    wire wire_12732;
    wire wire_12733;
    wire wire_12734;
    wire wire_12735;
    wire wire_12736;
    wire wire_12737;
    wire wire_12738;
    wire wire_12739;
    wire wire_12740;
    wire wire_12741;
    wire wire_12742;
    wire wire_12743;
    wire wire_12744;
    wire wire_12745;
    wire wire_12746;
    wire wire_12747;
    wire wire_12748;
    wire wire_12749;
    wire wire_12750;
    wire wire_12751;
    wire wire_12752;
    wire wire_12753;
    wire wire_12754;
    wire wire_12755;
    wire wire_12756;
    wire wire_12757;
    wire wire_12758;
    wire wire_12759;
    wire wire_12760;
    wire wire_12761;
    wire wire_12762;
    wire wire_12763;
    wire wire_12764;
    wire wire_12765;
    wire wire_12766;
    wire wire_12767;
    wire wire_12768;
    wire wire_12769;
    wire wire_12770;
    wire wire_12771;
    wire wire_12772;
    wire wire_12773;
    wire wire_12774;
    wire wire_12775;
    wire wire_12776;
    wire wire_12777;
    wire wire_12778;
    wire wire_12779;
    wire wire_12780;
    wire wire_12781;
    wire wire_12782;
    wire wire_12783;
    wire wire_12784;
    wire wire_12785;
    wire wire_12786;
    wire wire_12787;
    wire wire_12788;
    wire wire_12789;
    wire wire_12790;
    wire wire_12791;
    wire wire_12792;
    wire wire_12793;
    wire wire_12794;
    wire wire_12795;
    wire wire_12796;
    wire wire_12797;
    wire wire_12798;
    wire wire_12799;
    wire wire_12800;
    wire wire_12801;
    wire wire_12802;
    wire wire_12803;
    wire wire_12804;
    wire wire_12805;
    wire wire_12806;
    wire wire_12807;
    wire wire_12808;
    wire wire_12809;
    wire wire_12810;
    wire wire_12811;
    wire wire_12812;
    wire wire_12813;
    wire wire_12814;
    wire wire_12815;
    wire wire_12816;
    wire wire_12817;
    wire wire_12818;
    wire wire_12819;
    wire wire_12820;
    wire wire_12821;
    wire wire_12822;
    wire wire_12823;
    wire wire_12824;
    wire wire_12825;
    wire wire_12826;
    wire wire_12827;
    wire wire_12828;
    wire wire_12829;
    wire wire_12830;
    wire wire_12831;
    wire wire_12832;
    wire wire_12833;
    wire wire_12834;
    wire wire_12835;
    wire wire_12836;
    wire wire_12837;
    wire wire_12838;
    wire wire_12839;
    wire wire_12840;
    wire wire_12841;
    wire wire_12842;
    wire wire_12843;
    wire wire_12844;
    wire wire_12845;
    wire wire_12846;
    wire wire_12847;
    wire wire_12848;
    wire wire_12849;
    wire wire_12850;
    wire wire_12851;
    wire wire_12852;
    wire wire_12853;
    wire wire_12854;
    wire wire_12855;
    wire wire_12856;
    wire wire_12857;
    wire wire_12858;
    wire wire_12859;
    wire wire_12860;
    wire wire_12861;
    wire wire_12862;
    wire wire_12863;
    wire wire_12864;
    wire wire_12865;
    wire wire_12866;
    wire wire_12867;
    wire wire_12868;
    wire wire_12869;
    wire wire_12870;
    wire wire_12871;
    wire wire_12872;
    wire wire_12873;
    wire wire_12874;
    wire wire_12875;
    wire wire_12876;
    wire wire_12877;
    wire wire_12878;
    wire wire_12879;
    wire wire_12880;
    wire wire_12881;
    wire wire_12882;
    wire wire_12883;
    wire wire_12884;
    wire wire_12885;
    wire wire_12886;
    wire wire_12887;
    wire wire_12888;
    wire wire_12889;
    wire wire_12890;
    wire wire_12891;
    wire wire_12892;
    wire wire_12893;
    wire wire_12894;
    wire wire_12895;
    wire wire_12896;
    wire wire_12897;
    wire wire_12898;
    wire wire_12899;
    wire wire_12900;
    wire wire_12901;
    wire wire_12902;
    wire wire_12903;
    wire wire_12904;
    wire wire_12905;
    wire wire_12906;
    wire wire_12907;
    wire wire_12908;
    wire wire_12909;
    wire wire_12910;
    wire wire_12911;
    wire wire_12912;
    wire wire_12913;
    wire wire_12914;
    wire wire_12915;
    wire wire_12916;
    wire wire_12917;
    wire wire_12918;
    wire wire_12919;
    wire wire_12920;
    wire wire_12921;
    wire wire_12922;
    wire wire_12923;
    wire wire_12924;
    wire wire_12925;
    wire wire_12926;
    wire wire_12927;
    wire wire_12928;
    wire wire_12929;
    wire wire_12930;
    wire wire_12931;
    wire wire_12932;
    wire wire_12933;
    wire wire_12934;
    wire wire_12935;
    wire wire_12936;
    wire wire_12937;
    wire wire_12938;
    wire wire_12939;
    wire wire_12940;
    wire wire_12941;
    wire wire_12942;
    wire wire_12943;
    wire wire_12944;
    wire wire_12945;
    wire wire_12946;
    wire wire_12947;
    wire wire_12948;
    wire wire_12949;
    wire wire_12950;
    wire wire_12951;
    wire wire_12952;
    wire wire_12953;
    wire wire_12954;
    wire wire_12955;
    wire wire_12956;
    wire wire_12957;
    wire wire_12958;
    wire wire_12959;
    wire wire_12960;
    wire wire_12961;
    wire wire_12962;
    wire wire_12963;
    wire wire_12964;
    wire wire_12965;
    wire wire_12966;
    wire wire_12967;
    wire wire_12968;
    wire wire_12969;
    wire wire_12970;
    wire wire_12971;
    wire wire_12972;
    wire wire_12973;
    wire wire_12974;
    wire wire_12975;
    wire wire_12976;
    wire wire_12977;
    wire wire_12978;
    wire wire_12979;
    wire wire_12980;
    wire wire_12981;
    wire wire_12982;
    wire wire_12983;
    wire wire_12984;
    wire wire_12985;
    wire wire_12986;
    wire wire_12987;
    wire wire_12988;
    wire wire_12989;
    wire wire_12990;
    wire wire_12991;
    wire wire_12992;
    wire wire_12993;
    wire wire_12994;
    wire wire_12995;
    wire wire_12996;
    wire wire_12997;
    wire wire_12998;
    wire wire_12999;
    wire wire_13000;
    wire wire_13001;
    wire wire_13002;
    wire wire_13003;
    wire wire_13004;
    wire wire_13005;
    wire wire_13006;
    wire wire_13007;
    wire wire_13008;
    wire wire_13009;
    wire wire_13010;
    wire wire_13011;
    wire wire_13012;
    wire wire_13013;
    wire wire_13014;
    wire wire_13015;
    wire wire_13016;
    wire wire_13017;
    wire wire_13018;
    wire wire_13019;
    wire wire_13020;
    wire wire_13021;
    wire wire_13022;
    wire wire_13023;
    wire wire_13024;
    wire wire_13025;
    wire wire_13026;
    wire wire_13027;
    wire wire_13028;
    wire wire_13029;
    wire wire_13030;
    wire wire_13031;
    wire wire_13032;
    wire wire_13033;
    wire wire_13034;
    wire wire_13035;
    wire wire_13036;
    wire wire_13037;
    wire wire_13038;
    wire wire_13039;
    wire wire_13040;
    wire wire_13041;
    wire wire_13042;
    wire wire_13043;
    wire wire_13044;
    wire wire_13045;
    wire wire_13046;
    wire wire_13047;
    wire wire_13048;
    wire wire_13049;
    wire wire_13050;
    wire wire_13051;
    wire wire_13052;
    wire wire_13053;
    wire wire_13054;
    wire wire_13055;
    wire wire_13056;
    wire wire_13057;
    wire wire_13058;
    wire wire_13059;
    wire wire_13060;
    wire wire_13061;
    wire wire_13062;
    wire wire_13063;
    wire wire_13064;
    wire wire_13065;
    wire wire_13066;
    wire wire_13067;
    wire wire_13068;
    wire wire_13069;
    wire wire_13070;
    wire wire_13071;
    wire wire_13072;
    wire wire_13073;
    wire wire_13074;
    wire wire_13075;
    wire wire_13076;
    wire wire_13077;
    wire wire_13078;
    wire wire_13079;
    wire wire_13080;
    wire wire_13081;
    wire wire_13082;
    wire wire_13083;
    wire wire_13084;
    wire wire_13085;
    wire wire_13086;
    wire wire_13087;
    wire wire_13088;
    wire wire_13089;
    wire wire_13090;
    wire wire_13091;
    wire wire_13092;
    wire wire_13093;
    wire wire_13094;
    wire wire_13095;
    wire wire_13096;
    wire wire_13097;
    wire wire_13098;
    wire wire_13099;
    wire wire_13100;
    wire wire_13101;
    wire wire_13102;
    wire wire_13103;
    wire wire_13104;
    wire wire_13105;
    wire wire_13106;
    wire wire_13107;
    wire wire_13108;
    wire wire_13109;
    wire wire_13110;
    wire wire_13111;
    wire wire_13112;
    wire wire_13113;
    wire wire_13114;
    wire wire_13115;
    wire wire_13116;
    wire wire_13117;
    wire wire_13118;
    wire wire_13119;
    wire wire_13120;
    wire wire_13121;
    wire wire_13122;
    wire wire_13123;
    wire wire_13124;
    wire wire_13125;
    wire wire_13126;
    wire wire_13127;
    wire wire_13128;
    wire wire_13129;
    wire wire_13130;
    wire wire_13131;
    wire wire_13132;
    wire wire_13133;
    wire wire_13134;
    wire wire_13135;
    wire wire_13136;
    wire wire_13137;
    wire wire_13138;
    wire wire_13139;
    wire wire_13140;
    wire wire_13141;
    wire wire_13142;
    wire wire_13143;
    wire wire_13144;
    wire wire_13145;
    wire wire_13146;
    wire wire_13147;
    wire wire_13148;
    wire wire_13149;
    wire wire_13150;
    wire wire_13151;
    wire wire_13152;
    wire wire_13153;
    wire wire_13154;
    wire wire_13155;
    wire wire_13156;
    wire wire_13157;
    wire wire_13158;
    wire wire_13159;
    wire wire_13160;
    wire wire_13161;
    wire wire_13162;
    wire wire_13163;
    wire wire_13164;
    wire wire_13165;
    wire wire_13166;
    wire wire_13167;
    wire wire_13168;
    wire wire_13169;
    wire wire_13170;
    wire wire_13171;
    wire wire_13172;
    wire wire_13173;
    wire wire_13174;
    wire wire_13175;
    wire wire_13176;
    wire wire_13177;
    wire wire_13178;
    wire wire_13179;
    wire wire_13180;
    wire wire_13181;
    wire wire_13182;
    wire wire_13183;
    wire wire_13184;
    wire wire_13185;
    wire wire_13186;
    wire wire_13187;
    wire wire_13188;
    wire wire_13189;
    wire wire_13190;
    wire wire_13191;
    wire wire_13192;
    wire wire_13193;
    wire wire_13194;
    wire wire_13195;
    wire wire_13196;
    wire wire_13197;
    wire wire_13198;
    wire wire_13199;
    wire wire_13200;
    wire wire_13201;
    wire wire_13202;
    wire wire_13203;
    wire wire_13204;
    wire wire_13205;
    wire wire_13206;
    wire wire_13207;
    wire wire_13208;
    wire wire_13209;
    wire wire_13210;
    wire wire_13211;
    wire wire_13212;
    wire wire_13213;
    wire wire_13214;
    wire wire_13215;
    wire wire_13216;
    wire wire_13217;
    wire wire_13218;
    wire wire_13219;
    wire wire_13220;
    wire wire_13221;
    wire wire_13222;
    wire wire_13223;
    wire wire_13224;
    wire wire_13225;
    wire wire_13226;
    wire wire_13227;
    wire wire_13228;
    wire wire_13229;
    wire wire_13230;
    wire wire_13231;
    wire wire_13232;
    wire wire_13233;
    wire wire_13234;
    wire wire_13235;
    wire wire_13236;
    wire wire_13237;
    wire wire_13238;
    wire wire_13239;
    wire wire_13240;
    wire wire_13241;
    wire wire_13242;
    wire wire_13243;
    wire wire_13244;
    wire wire_13245;
    wire wire_13246;
    wire wire_13247;
    wire wire_13248;
    wire wire_13249;
    wire wire_13250;
    wire wire_13251;
    wire wire_13252;
    wire wire_13253;
    wire wire_13254;
    wire wire_13255;
    wire wire_13256;
    wire wire_13257;
    wire wire_13258;
    wire wire_13259;
    wire wire_13260;
    wire wire_13261;
    wire wire_13262;
    wire wire_13263;
    wire wire_13264;
    wire wire_13265;
    wire wire_13266;
    wire wire_13267;
    wire wire_13268;
    wire wire_13269;
    wire wire_13270;
    wire wire_13271;
    wire wire_13272;
    wire wire_13273;
    wire wire_13274;
    wire wire_13275;
    wire wire_13276;
    wire wire_13277;
    wire wire_13278;
    wire wire_13279;
    wire wire_13280;
    wire wire_13281;
    wire wire_13282;
    wire wire_13283;
    wire wire_13284;
    wire wire_13285;
    wire wire_13286;
    wire wire_13287;
    wire wire_13288;
    wire wire_13289;
    wire wire_13290;
    wire wire_13291;
    wire wire_13292;
    wire wire_13293;
    wire wire_13294;
    wire wire_13295;
    wire wire_13296;
    wire wire_13297;
    wire wire_13298;
    wire wire_13299;
    wire wire_13300;
    wire wire_13301;
    wire wire_13302;
    wire wire_13303;
    wire wire_13304;
    wire wire_13305;
    wire wire_13306;
    wire wire_13307;
    wire wire_13308;
    wire wire_13309;
    wire wire_13310;
    wire wire_13311;
    wire wire_13312;
    wire wire_13313;
    wire wire_13314;
    wire wire_13315;
    wire wire_13316;
    wire wire_13317;
    wire wire_13318;
    wire wire_13319;
    wire wire_13320;
    wire wire_13321;
    wire wire_13322;
    wire wire_13323;
    wire wire_13324;
    wire wire_13325;
    wire wire_13326;
    wire wire_13327;
    wire wire_13328;
    wire wire_13329;
    wire wire_13330;
    wire wire_13331;
    wire wire_13332;
    wire wire_13333;
    wire wire_13334;
    wire wire_13335;
    wire wire_13336;
    wire wire_13337;
    wire wire_13338;
    wire wire_13339;
    wire wire_13340;
    wire wire_13341;
    wire wire_13342;
    wire wire_13343;
    wire wire_13344;
    wire wire_13345;
    wire wire_13346;
    wire wire_13347;
    wire wire_13348;
    wire wire_13349;
    wire wire_13350;
    wire wire_13351;
    wire wire_13352;
    wire wire_13353;
    wire wire_13354;
    wire wire_13355;
    wire wire_13356;
    wire wire_13357;
    wire wire_13358;
    wire wire_13359;
    wire wire_13360;
    wire wire_13361;
    wire wire_13362;
    wire wire_13363;
    wire wire_13364;
    wire wire_13365;
    wire wire_13366;
    wire wire_13367;
    wire wire_13368;
    wire wire_13369;
    wire wire_13370;
    wire wire_13371;
    wire wire_13372;
    wire wire_13373;
    wire wire_13374;
    wire wire_13375;
    wire wire_13376;
    wire wire_13377;
    wire wire_13378;
    wire wire_13379;
    wire wire_13380;
    wire wire_13381;
    wire wire_13382;
    wire wire_13383;
    wire wire_13384;
    wire wire_13385;
    wire wire_13386;
    wire wire_13387;
    wire wire_13388;
    wire wire_13389;
    wire wire_13390;
    wire wire_13391;
    wire wire_13392;
    wire wire_13393;
    wire wire_13394;
    wire wire_13395;
    wire wire_13396;
    wire wire_13397;
    wire wire_13398;
    wire wire_13399;
    wire wire_13400;
    wire wire_13401;
    wire wire_13402;
    wire wire_13403;
    wire wire_13404;
    wire wire_13405;
    wire wire_13406;
    wire wire_13407;
    wire wire_13408;
    wire wire_13409;
    wire wire_13410;
    wire wire_13411;
    wire wire_13412;
    wire wire_13413;
    wire wire_13414;
    wire wire_13415;
    wire wire_13416;
    wire wire_13417;
    wire wire_13418;
    wire wire_13419;
    wire wire_13420;
    wire wire_13421;
    wire wire_13422;
    wire wire_13423;
    wire wire_13424;
    wire wire_13425;
    wire wire_13426;
    wire wire_13427;
    wire wire_13428;
    wire wire_13429;
    wire wire_13430;
    wire wire_13431;
    wire wire_13432;
    wire wire_13433;
    wire wire_13434;
    wire wire_13435;
    wire wire_13436;
    wire wire_13437;
    wire wire_13438;
    wire wire_13439;
    wire wire_13440;
    wire wire_13441;
    wire wire_13442;
    wire wire_13443;
    wire wire_13444;
    wire wire_13445;
    wire wire_13446;
    wire wire_13447;
    wire wire_13448;
    wire wire_13449;
    wire wire_13450;
    wire wire_13451;
    wire wire_13452;
    wire wire_13453;
    wire wire_13454;
    wire wire_13455;
    wire wire_13456;
    wire wire_13457;
    wire wire_13458;
    wire wire_13459;
    wire wire_13460;
    wire wire_13461;
    wire wire_13462;
    wire wire_13463;
    wire wire_13464;
    wire wire_13465;
    wire wire_13466;
    wire wire_13467;
    wire wire_13468;
    wire wire_13469;
    wire wire_13470;
    wire wire_13471;
    wire wire_13472;
    wire wire_13473;
    wire wire_13474;
    wire wire_13475;
    wire wire_13476;
    wire wire_13477;
    wire wire_13478;
    wire wire_13479;
    wire wire_13480;
    wire wire_13481;
    wire wire_13482;
    wire wire_13483;
    wire wire_13484;
    wire wire_13485;
    wire wire_13486;
    wire wire_13487;
    wire wire_13488;
    wire wire_13489;
    wire wire_13490;
    wire wire_13491;
    wire wire_13492;
    wire wire_13493;
    wire wire_13494;
    wire wire_13495;
    wire wire_13496;
    wire wire_13497;
    wire wire_13498;
    wire wire_13499;
    wire wire_13500;
    wire wire_13501;
    wire wire_13502;
    wire wire_13503;
    wire wire_13504;
    wire wire_13505;
    wire wire_13506;
    wire wire_13507;
    wire wire_13508;
    wire wire_13509;
    wire wire_13510;
    wire wire_13511;
    wire wire_13512;
    wire wire_13513;
    wire wire_13514;
    wire wire_13515;
    wire wire_13516;
    wire wire_13517;
    wire wire_13518;
    wire wire_13519;
    wire wire_13520;
    wire wire_13521;
    wire wire_13522;
    wire wire_13523;
    wire wire_13524;
    wire wire_13525;
    wire wire_13526;
    wire wire_13527;
    wire wire_13528;
    wire wire_13529;
    wire wire_13530;
    wire wire_13531;
    wire wire_13532;
    wire wire_13533;
    wire wire_13534;
    wire wire_13535;
    wire wire_13536;
    wire wire_13537;
    wire wire_13538;
    wire wire_13539;
    wire wire_13540;
    wire wire_13541;
    wire wire_13542;
    wire wire_13543;
    wire wire_13544;
    wire wire_13545;
    wire wire_13546;
    wire wire_13547;
    wire wire_13548;
    wire wire_13549;
    wire wire_13550;
    wire wire_13551;
    wire wire_13552;
    wire wire_13553;
    wire wire_13554;
    wire wire_13555;
    wire wire_13556;
    wire wire_13557;
    wire wire_13558;
    wire wire_13559;
    wire wire_13560;
    wire wire_13561;
    wire wire_13562;
    wire wire_13563;
    wire wire_13564;
    wire wire_13565;
    wire wire_13566;
    wire wire_13567;
    wire wire_13568;
    wire wire_13569;
    wire wire_13570;
    wire wire_13571;
    wire wire_13572;
    wire wire_13573;
    wire wire_13574;
    wire wire_13575;
    wire wire_13576;
    wire wire_13577;
    wire wire_13578;
    wire wire_13579;
    wire wire_13580;
    wire wire_13581;
    wire wire_13582;
    wire wire_13583;
    wire wire_13584;
    wire wire_13585;
    wire wire_13586;
    wire wire_13587;
    wire wire_13588;
    wire wire_13589;
    wire wire_13590;
    wire wire_13591;
    wire wire_13592;
    wire wire_13593;
    wire wire_13594;
    wire wire_13595;
    wire wire_13596;
    wire wire_13597;
    wire wire_13598;
    wire wire_13599;
    wire wire_13600;
    wire wire_13601;
    wire wire_13602;
    wire wire_13603;
    wire wire_13604;
    wire wire_13605;
    wire wire_13606;
    wire wire_13607;
    wire wire_13608;
    wire wire_13609;
    wire wire_13610;
    wire wire_13611;
    wire wire_13612;
    wire wire_13613;
    wire wire_13614;
    wire wire_13615;
    wire wire_13616;
    wire wire_13617;
    wire wire_13618;
    wire wire_13619;
    wire wire_13620;
    wire wire_13621;
    wire wire_13622;
    wire wire_13623;
    wire wire_13624;
    wire wire_13625;
    wire wire_13626;
    wire wire_13627;
    wire wire_13628;
    wire wire_13629;
    wire wire_13630;
    wire wire_13631;
    wire wire_13632;
    wire wire_13633;
    wire wire_13634;
    wire wire_13635;
    wire wire_13636;
    wire wire_13637;
    wire wire_13638;
    wire wire_13639;
    wire wire_13640;
    wire wire_13641;
    wire wire_13642;
    wire wire_13643;
    wire wire_13644;
    wire wire_13645;
    wire wire_13646;
    wire wire_13647;
    wire wire_13648;
    wire wire_13649;
    wire wire_13650;
    wire wire_13651;
    wire wire_13652;
    wire wire_13653;
    wire wire_13654;
    wire wire_13655;
    wire wire_13656;
    wire wire_13657;
    wire wire_13658;
    wire wire_13659;
    wire wire_13660;
    wire wire_13661;
    wire wire_13662;
    wire wire_13663;
    wire wire_13664;
    wire wire_13665;
    wire wire_13666;
    wire wire_13667;
    wire wire_13668;
    wire wire_13669;
    wire wire_13670;
    wire wire_13671;
    wire wire_13672;
    wire wire_13673;
    wire wire_13674;
    wire wire_13675;
    wire wire_13676;
    wire wire_13677;
    wire wire_13678;
    wire wire_13679;
    wire wire_13680;
    wire wire_13681;
    wire wire_13682;
    wire wire_13683;
    wire wire_13684;
    wire wire_13685;
    wire wire_13686;
    wire wire_13687;
    wire wire_13688;
    wire wire_13689;
    wire wire_13690;
    wire wire_13691;
    wire wire_13692;
    wire wire_13693;
    wire wire_13694;
    wire wire_13695;
    wire wire_13696;
    wire wire_13697;
    wire wire_13698;
    wire wire_13699;
    wire wire_13700;
    wire wire_13701;
    wire wire_13702;
    wire wire_13703;
    wire wire_13704;
    wire wire_13705;
    wire wire_13706;
    wire wire_13707;
    wire wire_13708;
    wire wire_13709;
    wire wire_13710;
    wire wire_13711;
    wire wire_13712;
    wire wire_13713;
    wire wire_13714;
    wire wire_13715;
    wire wire_13716;
    wire wire_13717;
    wire wire_13718;
    wire wire_13719;
    wire wire_13720;
    wire wire_13721;
    wire wire_13722;
    wire wire_13723;
    wire wire_13724;
    wire wire_13725;
    wire wire_13726;
    wire wire_13727;
    wire wire_13728;
    wire wire_13729;
    wire wire_13730;
    wire wire_13731;
    wire wire_13732;
    wire wire_13733;
    wire wire_13734;
    wire wire_13735;
    wire wire_13736;
    wire wire_13737;
    wire wire_13738;
    wire wire_13739;
    wire wire_13740;
    wire wire_13741;
    wire wire_13742;
    wire wire_13743;
    wire wire_13744;
    wire wire_13745;
    wire wire_13746;
    wire wire_13747;
    wire wire_13748;
    wire wire_13749;
    wire wire_13750;
    wire wire_13751;
    wire wire_13752;
    wire wire_13753;
    wire wire_13754;
    wire wire_13755;
    wire wire_13756;
    wire wire_13757;
    wire wire_13758;
    wire wire_13759;
    wire wire_13760;
    wire wire_13761;
    wire wire_13762;
    wire wire_13763;
    wire wire_13764;
    wire wire_13765;
    wire wire_13766;
    wire wire_13767;
    wire wire_13768;
    wire wire_13769;
    wire wire_13770;
    wire wire_13771;
    wire wire_13772;
    wire wire_13773;
    wire wire_13774;
    wire wire_13775;
    wire wire_13776;
    wire wire_13777;
    wire wire_13778;
    wire wire_13779;
    wire wire_13780;
    wire wire_13781;
    wire wire_13782;
    wire wire_13783;
    wire wire_13784;
    wire wire_13785;
    wire wire_13786;
    wire wire_13787;
    wire wire_13788;
    wire wire_13789;
    wire wire_13790;
    wire wire_13791;
    wire wire_13792;
    wire wire_13793;
    wire wire_13794;
    wire wire_13795;
    wire wire_13796;
    wire wire_13797;
    wire wire_13798;
    wire wire_13799;
    wire wire_13800;
    wire wire_13801;
    wire wire_13802;
    wire wire_13803;
    wire wire_13804;
    wire wire_13805;
    wire wire_13806;
    wire wire_13807;
    wire wire_13808;
    wire wire_13809;
    wire wire_13810;
    wire wire_13811;
    wire wire_13812;
    wire wire_13813;
    wire wire_13814;
    wire wire_13815;
    wire wire_13816;
    wire wire_13817;
    wire wire_13818;
    wire wire_13819;
    wire wire_13820;
    wire wire_13821;
    wire wire_13822;
    wire wire_13823;
    wire wire_13824;
    wire wire_13825;
    wire wire_13826;
    wire wire_13827;
    wire wire_13828;
    wire wire_13829;
    wire wire_13830;
    wire wire_13831;
    wire wire_13832;
    wire wire_13833;
    wire wire_13834;
    wire wire_13835;
    wire wire_13836;
    wire wire_13837;
    wire wire_13838;
    wire wire_13839;
    wire wire_13840;
    wire wire_13841;
    wire wire_13842;
    wire wire_13843;
    wire wire_13844;
    wire wire_13845;
    wire wire_13846;
    wire wire_13847;
    wire wire_13848;
    wire wire_13849;
    wire wire_13850;
    wire wire_13851;
    wire wire_13852;
    wire wire_13853;
    wire wire_13854;
    wire wire_13855;
    wire wire_13856;
    wire wire_13857;
    wire wire_13858;
    wire wire_13859;
    wire wire_13860;
    wire wire_13861;
    wire wire_13862;
    wire wire_13863;
    wire wire_13864;
    wire wire_13865;
    wire wire_13866;
    wire wire_13867;
    wire wire_13868;
    wire wire_13869;
    wire wire_13870;
    wire wire_13871;
    wire wire_13872;
    wire wire_13873;
    wire wire_13874;
    wire wire_13875;
    wire wire_13876;
    wire wire_13877;
    wire wire_13878;
    wire wire_13879;
    wire wire_13880;
    wire wire_13881;
    wire wire_13882;
    wire wire_13883;
    wire wire_13884;
    wire wire_13885;
    wire wire_13886;
    wire wire_13887;
    wire wire_13888;
    wire wire_13889;
    wire wire_13890;
    wire wire_13891;
    wire wire_13892;
    wire wire_13893;
    wire wire_13894;
    wire wire_13895;
    wire wire_13896;
    wire wire_13897;
    wire wire_13898;
    wire wire_13899;
    wire wire_13900;
    wire wire_13901;
    wire wire_13902;
    wire wire_13903;
    wire wire_13904;
    wire wire_13905;
    wire wire_13906;
    wire wire_13907;
    wire wire_13908;
    wire wire_13909;
    wire wire_13910;
    wire wire_13911;
    wire wire_13912;
    wire wire_13913;
    wire wire_13914;
    wire wire_13915;
    wire wire_13916;
    wire wire_13917;
    wire wire_13918;
    wire wire_13919;
    wire wire_13920;
    wire wire_13921;
    wire wire_13922;
    wire wire_13923;
    wire wire_13924;
    wire wire_13925;
    wire wire_13926;
    wire wire_13927;
    wire wire_13928;
    wire wire_13929;
    wire wire_13930;
    wire wire_13931;
    wire wire_13932;
    wire wire_13933;
    wire wire_13934;
    wire wire_13935;
    wire wire_13936;
    wire wire_13937;
    wire wire_13938;
    wire wire_13939;
    wire wire_13940;
    wire wire_13941;
    wire wire_13942;
    wire wire_13943;
    wire wire_13944;
    wire wire_13945;
    wire wire_13946;
    wire wire_13947;
    wire wire_13948;
    wire wire_13949;
    wire wire_13950;
    wire wire_13951;
    wire wire_13952;
    wire wire_13953;
    wire wire_13954;
    wire wire_13955;
    wire wire_13956;
    wire wire_13957;
    wire wire_13958;
    wire wire_13959;
    wire wire_13960;
    wire wire_13961;
    wire wire_13962;
    wire wire_13963;
    wire wire_13964;
    wire wire_13965;
    wire wire_13966;
    wire wire_13967;
    wire wire_13968;
    wire wire_13969;
    wire wire_13970;
    wire wire_13971;
    wire wire_13972;
    wire wire_13973;
    wire wire_13974;
    wire wire_13975;
    wire wire_13976;
    wire wire_13977;
    wire wire_13978;
    wire wire_13979;
    wire wire_13980;
    wire wire_13981;
    wire wire_13982;
    wire wire_13983;
    wire wire_13984;
    wire wire_13985;
    wire wire_13986;
    wire wire_13987;
    wire wire_13988;
    wire wire_13989;
    wire wire_13990;
    wire wire_13991;
    wire wire_13992;
    wire wire_13993;
    wire wire_13994;
    wire wire_13995;
    wire wire_13996;
    wire wire_13997;
    wire wire_13998;
    wire wire_13999;
    wire wire_14000;
    wire wire_14001;
    wire wire_14002;
    wire wire_14003;
    wire wire_14004;
    wire wire_14005;
    wire wire_14006;
    wire wire_14007;
    wire wire_14008;
    wire wire_14009;
    wire wire_14010;
    wire wire_14011;
    wire wire_14012;
    wire wire_14013;
    wire wire_14014;
    wire wire_14015;
    wire wire_14016;
    wire wire_14017;
    wire wire_14018;
    wire wire_14019;
    wire wire_14020;
    wire wire_14021;
    wire wire_14022;
    wire wire_14023;
    wire wire_14024;
    wire wire_14025;
    wire wire_14026;
    wire wire_14027;
    wire wire_14028;
    wire wire_14029;
    wire wire_14030;
    wire wire_14031;
    wire wire_14032;
    wire wire_14033;
    wire wire_14034;
    wire wire_14035;
    wire wire_14036;
    wire wire_14037;
    wire wire_14038;
    wire wire_14039;
    wire wire_14040;
    wire wire_14041;
    wire wire_14042;
    wire wire_14043;
    wire wire_14044;
    wire wire_14045;
    wire wire_14046;
    wire wire_14047;
    wire wire_14048;
    wire wire_14049;
    wire wire_14050;
    wire wire_14051;
    wire wire_14052;
    wire wire_14053;
    wire wire_14054;
    wire wire_14055;
    wire wire_14056;
    wire wire_14057;
    wire wire_14058;
    wire wire_14059;
    wire wire_14060;
    wire wire_14061;
    wire wire_14062;
    wire wire_14063;
    wire wire_14064;
    wire wire_14065;
    wire wire_14066;
    wire wire_14067;
    wire wire_14068;
    wire wire_14069;
    wire wire_14070;
    wire wire_14071;
    wire wire_14072;
    wire wire_14073;
    wire wire_14074;
    wire wire_14075;
    wire wire_14076;
    wire wire_14077;
    wire wire_14078;
    wire wire_14079;
    wire wire_14080;
    wire wire_14081;
    wire wire_14082;
    wire wire_14083;
    wire wire_14084;
    wire wire_14085;
    wire wire_14086;
    wire wire_14087;
    wire wire_14088;
    wire wire_14089;
    wire wire_14090;
    wire wire_14091;
    wire wire_14092;
    wire wire_14093;
    wire wire_14094;
    wire wire_14095;
    wire wire_14096;
    wire wire_14097;
    wire wire_14098;
    wire wire_14099;
    wire wire_14100;
    wire wire_14101;
    wire wire_14102;
    wire wire_14103;
    wire wire_14104;
    wire wire_14105;
    wire wire_14106;
    wire wire_14107;
    wire wire_14108;
    wire wire_14109;
    wire wire_14110;
    wire wire_14111;
    wire wire_14112;
    wire wire_14113;
    wire wire_14114;
    wire wire_14115;
    wire wire_14116;
    wire wire_14117;
    wire wire_14118;
    wire wire_14119;
    wire wire_14120;
    wire wire_14121;
    wire wire_14122;
    wire wire_14123;
    wire wire_14124;
    wire wire_14125;
    wire wire_14126;
    wire wire_14127;
    wire wire_14128;
    wire wire_14129;
    wire wire_14130;
    wire wire_14131;
    wire wire_14132;
    wire wire_14133;
    wire wire_14134;
    wire wire_14135;
    wire wire_14136;
    wire wire_14137;
    wire wire_14138;
    wire wire_14139;
    wire wire_14140;
    wire wire_14141;
    wire wire_14142;
    wire wire_14143;
    wire wire_14144;
    wire wire_14145;
    wire wire_14146;
    wire wire_14147;
    wire wire_14148;
    wire wire_14149;
    wire wire_14150;
    wire wire_14151;
    wire wire_14152;
    wire wire_14153;
    wire wire_14154;
    wire wire_14155;
    wire wire_14156;
    wire wire_14157;
    wire wire_14158;
    wire wire_14159;
    wire wire_14160;
    wire wire_14161;
    wire wire_14162;
    wire wire_14163;
    wire wire_14164;
    wire wire_14165;
    wire wire_14166;
    wire wire_14167;
    wire wire_14168;
    wire wire_14169;
    wire wire_14170;
    wire wire_14171;
    wire wire_14172;
    wire wire_14173;
    wire wire_14174;
    wire wire_14175;
    wire wire_14176;
    wire wire_14177;
    wire wire_14178;
    wire wire_14179;
    wire wire_14180;
    wire wire_14181;
    wire wire_14182;
    wire wire_14183;
    wire wire_14184;
    wire wire_14185;
    wire wire_14186;
    wire wire_14187;
    wire wire_14188;
    wire wire_14189;
    wire wire_14190;
    wire wire_14191;
    wire wire_14192;
    wire wire_14193;
    wire wire_14194;
    wire wire_14195;
    wire wire_14196;
    wire wire_14197;
    wire wire_14198;
    wire wire_14199;
    wire wire_14200;
    wire wire_14201;
    wire wire_14202;
    wire wire_14203;
    wire wire_14204;
    wire wire_14205;
    wire wire_14206;
    wire wire_14207;
    wire wire_14208;
    wire wire_14209;
    wire wire_14210;
    wire wire_14211;
    wire wire_14212;
    wire wire_14213;
    wire wire_14214;
    wire wire_14215;
    wire wire_14216;
    wire wire_14217;
    wire wire_14218;
    wire wire_14219;
    wire wire_14220;
    wire wire_14221;
    wire wire_14222;
    wire wire_14223;
    wire wire_14224;
    wire wire_14225;
    wire wire_14226;
    wire wire_14227;
    wire wire_14228;
    wire wire_14229;
    wire wire_14230;
    wire wire_14231;
    wire wire_14232;
    wire wire_14233;
    wire wire_14234;
    wire wire_14235;
    wire wire_14236;
    wire wire_14237;
    wire wire_14238;
    wire wire_14239;
    wire wire_14240;
    wire wire_14241;
    wire wire_14242;
    wire wire_14243;
    wire wire_14244;
    wire wire_14245;
    wire wire_14246;
    wire wire_14247;
    wire wire_14248;
    wire wire_14249;
    wire wire_14250;
    wire wire_14251;
    wire wire_14252;
    wire wire_14253;
    wire wire_14254;
    wire wire_14255;
    wire wire_14256;
    wire wire_14257;
    wire wire_14258;
    wire wire_14259;
    wire wire_14260;
    wire wire_14261;
    wire wire_14262;
    wire wire_14263;
    wire wire_14264;
    wire wire_14265;
    wire wire_14266;
    wire wire_14267;
    wire wire_14268;
    wire wire_14269;
    wire wire_14270;
    wire wire_14271;
    wire wire_14272;
    wire wire_14273;
    wire wire_14274;
    wire wire_14275;
    wire wire_14276;
    wire wire_14277;
    wire wire_14278;
    wire wire_14279;
    wire wire_14280;
    wire wire_14281;
    wire wire_14282;
    wire wire_14283;
    wire wire_14284;
    wire wire_14285;
    wire wire_14286;
    wire wire_14287;
    wire wire_14288;
    wire wire_14289;
    wire wire_14290;
    wire wire_14291;
    wire wire_14292;
    wire wire_14293;
    wire wire_14294;
    wire wire_14295;
    wire wire_14296;
    wire wire_14297;
    wire wire_14298;
    wire wire_14299;
    wire wire_14300;
    wire wire_14301;
    wire wire_14302;
    wire wire_14303;
    wire wire_14304;
    wire wire_14305;
    wire wire_14306;
    wire wire_14307;
    wire wire_14308;
    wire wire_14309;
    wire wire_14310;
    wire wire_14311;
    wire wire_14312;
    wire wire_14313;
    wire wire_14314;
    wire wire_14315;
    wire wire_14316;
    wire wire_14317;
    wire wire_14318;
    wire wire_14319;
    wire wire_14320;
    wire wire_14321;
    wire wire_14322;
    wire wire_14323;
    wire wire_14324;
    wire wire_14325;
    wire wire_14326;
    wire wire_14327;
    wire wire_14328;
    wire wire_14329;
    wire wire_14330;
    wire wire_14331;
    wire wire_14332;
    wire wire_14333;
    wire wire_14334;
    wire wire_14335;
    wire wire_14336;
    wire wire_14337;
    wire wire_14338;
    wire wire_14339;
    wire wire_14340;
    wire wire_14341;
    wire wire_14342;
    wire wire_14343;
    wire wire_14344;
    wire wire_14345;
    wire wire_14346;
    wire wire_14347;
    wire wire_14348;
    wire wire_14349;
    wire wire_14350;
    wire wire_14351;
    wire wire_14352;
    wire wire_14353;
    wire wire_14354;
    wire wire_14355;
    wire wire_14356;
    wire wire_14357;
    wire wire_14358;
    wire wire_14359;
    wire wire_14360;
    wire wire_14361;
    wire wire_14362;
    wire wire_14363;
    wire wire_14364;
    wire wire_14365;
    wire wire_14366;
    wire wire_14367;
    wire wire_14368;
    wire wire_14369;
    wire wire_14370;
    wire wire_14371;
    wire wire_14372;
    wire wire_14373;
    wire wire_14374;
    wire wire_14375;
    wire wire_14376;
    wire wire_14377;
    wire wire_14378;
    wire wire_14379;
    wire wire_14380;
    wire wire_14381;
    wire wire_14382;
    wire wire_14383;
    wire wire_14384;
    wire wire_14385;
    wire wire_14386;
    wire wire_14387;
    wire wire_14388;
    wire wire_14389;
    wire wire_14390;
    wire wire_14391;
    wire wire_14392;
    wire wire_14393;
    wire wire_14394;
    wire wire_14395;
    wire wire_14396;
    wire wire_14397;
    wire wire_14398;
    wire wire_14399;
    wire wire_14400;
    wire wire_14401;
    wire wire_14402;
    wire wire_14403;
    wire wire_14404;
    wire wire_14405;
    wire wire_14406;
    wire wire_14407;
    wire wire_14408;
    wire wire_14409;
    wire wire_14410;
    wire wire_14411;
    wire wire_14412;
    wire wire_14413;
    wire wire_14414;
    wire wire_14415;
    wire wire_14416;
    wire wire_14417;
    wire wire_14418;
    wire wire_14419;
    wire wire_14420;
    wire wire_14421;
    wire wire_14422;
    wire wire_14423;
    wire wire_14424;
    wire wire_14425;
    wire wire_14426;
    wire wire_14427;
    wire wire_14428;
    wire wire_14429;
    wire wire_14430;
    wire wire_14431;
    wire wire_14432;
    wire wire_14433;
    wire wire_14434;
    wire wire_14435;
    wire wire_14436;
    wire wire_14437;
    wire wire_14438;
    wire wire_14439;
    wire wire_14440;
    wire wire_14441;
    wire wire_14442;
    wire wire_14443;
    wire wire_14444;
    wire wire_14445;
    wire wire_14446;
    wire wire_14447;
    wire wire_14448;
    wire wire_14449;
    wire wire_14450;
    wire wire_14451;
    wire wire_14452;
    wire wire_14453;
    wire wire_14454;
    wire wire_14455;
    wire wire_14456;
    wire wire_14457;
    wire wire_14458;
    wire wire_14459;
    wire wire_14460;
    wire wire_14461;
    wire wire_14462;
    wire wire_14463;
    wire wire_14464;
    wire wire_14465;
    wire wire_14466;
    wire wire_14467;
    wire wire_14468;
    wire wire_14469;
    wire wire_14470;
    wire wire_14471;
    wire wire_14472;
    wire wire_14473;
    wire wire_14474;
    wire wire_14475;
    wire wire_14476;
    wire wire_14477;
    wire wire_14478;
    wire wire_14479;
    wire wire_14480;
    wire wire_14481;
    wire wire_14482;
    wire wire_14483;
    wire wire_14484;
    wire wire_14485;
    wire wire_14486;
    wire wire_14487;
    wire wire_14488;
    wire wire_14489;
    wire wire_14490;
    wire wire_14491;
    wire wire_14492;
    wire wire_14493;
    wire wire_14494;
    wire wire_14495;
    wire wire_14496;
    wire wire_14497;
    wire wire_14498;
    wire wire_14499;
    wire wire_14500;
    wire wire_14501;
    wire wire_14502;
    wire wire_14503;
    wire wire_14504;
    wire wire_14505;
    wire wire_14506;
    wire wire_14507;
    wire wire_14508;
    wire wire_14509;
    wire wire_14510;
    wire wire_14511;
    wire wire_14512;
    wire wire_14513;
    wire wire_14514;
    wire wire_14515;
    wire wire_14516;
    wire wire_14517;
    wire wire_14518;
    wire wire_14519;
    wire wire_14520;
    wire wire_14521;
    wire wire_14522;
    wire wire_14523;
    wire wire_14524;
    wire wire_14525;
    wire wire_14526;
    wire wire_14527;
    wire wire_14528;
    wire wire_14529;
    wire wire_14530;
    wire wire_14531;
    wire wire_14532;
    wire wire_14533;
    wire wire_14534;
    wire wire_14535;
    wire wire_14536;
    wire wire_14537;
    wire wire_14538;
    wire wire_14539;
    wire wire_14540;
    wire wire_14541;
    wire wire_14542;
    wire wire_14543;
    wire wire_14544;
    wire wire_14545;
    wire wire_14546;
    wire wire_14547;
    wire wire_14548;
    wire wire_14549;
    wire wire_14550;
    wire wire_14551;
    wire wire_14552;
    wire wire_14553;
    wire wire_14554;
    wire wire_14555;
    wire wire_14556;
    wire wire_14557;
    wire wire_14558;
    wire wire_14559;
    wire wire_14560;
    wire wire_14561;
    wire wire_14562;
    wire wire_14563;
    wire wire_14564;
    wire wire_14565;
    wire wire_14566;
    wire wire_14567;
    wire wire_14568;
    wire wire_14569;
    wire wire_14570;
    wire wire_14571;
    wire wire_14572;
    wire wire_14573;
    wire wire_14574;
    wire wire_14575;
    wire wire_14576;
    wire wire_14577;
    wire wire_14578;
    wire wire_14579;
    wire wire_14580;
    wire wire_14581;
    wire wire_14582;
    wire wire_14583;
    wire wire_14584;
    wire wire_14585;
    wire wire_14586;
    wire wire_14587;
    wire wire_14588;
    wire wire_14589;
    wire wire_14590;
    wire wire_14591;
    wire wire_14592;
    wire wire_14593;
    wire wire_14594;
    wire wire_14595;
    wire wire_14596;
    wire wire_14597;
    wire wire_14598;
    wire wire_14599;
    wire wire_14600;
    wire wire_14601;
    wire wire_14602;
    wire wire_14603;
    wire wire_14604;
    wire wire_14605;
    wire wire_14606;
    wire wire_14607;
    wire wire_14608;
    wire wire_14609;
    wire wire_14610;
    wire wire_14611;
    wire wire_14612;
    wire wire_14613;
    wire wire_14614;
    wire wire_14615;
    wire wire_14616;
    wire wire_14617;
    wire wire_14618;
    wire wire_14619;
    wire wire_14620;
    wire wire_14621;
    wire wire_14622;
    wire wire_14623;
    wire wire_14624;
    wire wire_14625;
    wire wire_14626;
    wire wire_14627;
    wire wire_14628;
    wire wire_14629;
    wire wire_14630;
    wire wire_14631;
    wire wire_14632;
    wire wire_14633;
    wire wire_14634;
    wire wire_14635;
    wire wire_14636;
    wire wire_14637;
    wire wire_14638;
    wire wire_14639;
    wire wire_14640;
    wire wire_14641;
    wire wire_14642;
    wire wire_14643;
    wire wire_14644;
    wire wire_14645;
    wire wire_14646;
    wire wire_14647;
    wire wire_14648;
    wire wire_14649;
    wire wire_14650;
    wire wire_14651;
    wire wire_14652;
    wire wire_14653;
    wire wire_14654;
    wire wire_14655;
    wire wire_14656;
    wire wire_14657;
    wire wire_14658;
    wire wire_14659;
    wire wire_14660;
    wire wire_14661;
    wire wire_14662;
    wire wire_14663;
    wire wire_14664;
    wire wire_14665;
    wire wire_14666;
    wire wire_14667;
    wire wire_14668;
    wire wire_14669;
    wire wire_14670;
    wire wire_14671;
    wire wire_14672;
    wire wire_14673;
    wire wire_14674;
    wire wire_14675;
    wire wire_14676;
    wire wire_14677;
    wire wire_14678;
    wire wire_14679;
    wire wire_14680;
    wire wire_14681;
    wire wire_14682;
    wire wire_14683;
    wire wire_14684;
    wire wire_14685;
    wire wire_14686;
    wire wire_14687;
    wire wire_14688;
    wire wire_14689;
    wire wire_14690;
    wire wire_14691;
    wire wire_14692;
    wire wire_14693;
    wire wire_14694;
    wire wire_14695;
    wire wire_14696;
    wire wire_14697;
    wire wire_14698;
    wire wire_14699;


    // FPGA IO TILES DECLARE
    wire [254:0] io_tile_1_0_chanxy_in;
    wire [74:0] io_tile_1_0_chanxy_out;
    wire [95:0] io_tile_1_0_ipin_in;
    wire [7:0] io_tile_1_0_opin_out;
    io_tile_sp_0 io_tile_1_0(
            .io_chanxy_in(io_tile_1_0_chanxy_in),
            .io_chanxy_out(io_tile_1_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[9:5]),
            .io_io_input(left_in[7:0]),
            .io_io_output(left_out[7:0]),
            .io_ipin_in(io_tile_1_0_ipin_in),
            .io_opin_out(io_tile_1_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_2_0_chanxy_in;
    wire [29:0] io_tile_2_0_chanxy_out;
    wire [95:0] io_tile_2_0_ipin_in;
    wire [7:0] io_tile_2_0_opin_out;
    io_tile_sp_1 io_tile_2_0(
            .io_chanxy_in(io_tile_2_0_chanxy_in),
            .io_chanxy_out(io_tile_2_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[36:32]),
            .io_io_input(left_in[15:8]),
            .io_io_output(left_out[15:8]),
            .io_ipin_in(io_tile_2_0_ipin_in),
            .io_opin_out(io_tile_2_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_3_0_chanxy_in;
    wire [29:0] io_tile_3_0_chanxy_out;
    wire [95:0] io_tile_3_0_ipin_in;
    wire [7:0] io_tile_3_0_opin_out;
    io_tile_sp_2 io_tile_3_0(
            .io_chanxy_in(io_tile_3_0_chanxy_in),
            .io_chanxy_out(io_tile_3_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[62:58]),
            .io_io_input(left_in[23:16]),
            .io_io_output(left_out[23:16]),
            .io_ipin_in(io_tile_3_0_ipin_in),
            .io_opin_out(io_tile_3_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_4_0_chanxy_in;
    wire [29:0] io_tile_4_0_chanxy_out;
    wire [95:0] io_tile_4_0_ipin_in;
    wire [7:0] io_tile_4_0_opin_out;
    io_tile_sp_3 io_tile_4_0(
            .io_chanxy_in(io_tile_4_0_chanxy_in),
            .io_chanxy_out(io_tile_4_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[88:84]),
            .io_io_input(left_in[31:24]),
            .io_io_output(left_out[31:24]),
            .io_ipin_in(io_tile_4_0_ipin_in),
            .io_opin_out(io_tile_4_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_5_0_chanxy_in;
    wire [29:0] io_tile_5_0_chanxy_out;
    wire [95:0] io_tile_5_0_ipin_in;
    wire [7:0] io_tile_5_0_opin_out;
    io_tile_sp_4 io_tile_5_0(
            .io_chanxy_in(io_tile_5_0_chanxy_in),
            .io_chanxy_out(io_tile_5_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[114:110]),
            .io_io_input(left_in[39:32]),
            .io_io_output(left_out[39:32]),
            .io_ipin_in(io_tile_5_0_ipin_in),
            .io_opin_out(io_tile_5_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_6_0_chanxy_in;
    wire [29:0] io_tile_6_0_chanxy_out;
    wire [95:0] io_tile_6_0_ipin_in;
    wire [7:0] io_tile_6_0_opin_out;
    io_tile_sp_5 io_tile_6_0(
            .io_chanxy_in(io_tile_6_0_chanxy_in),
            .io_chanxy_out(io_tile_6_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[140:136]),
            .io_io_input(left_in[47:40]),
            .io_io_output(left_out[47:40]),
            .io_ipin_in(io_tile_6_0_ipin_in),
            .io_opin_out(io_tile_6_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_7_0_chanxy_in;
    wire [29:0] io_tile_7_0_chanxy_out;
    wire [95:0] io_tile_7_0_ipin_in;
    wire [7:0] io_tile_7_0_opin_out;
    io_tile_sp_6 io_tile_7_0(
            .io_chanxy_in(io_tile_7_0_chanxy_in),
            .io_chanxy_out(io_tile_7_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[166:162]),
            .io_io_input(left_in[55:48]),
            .io_io_output(left_out[55:48]),
            .io_ipin_in(io_tile_7_0_ipin_in),
            .io_opin_out(io_tile_7_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_8_0_chanxy_in;
    wire [29:0] io_tile_8_0_chanxy_out;
    wire [95:0] io_tile_8_0_ipin_in;
    wire [7:0] io_tile_8_0_opin_out;
    io_tile_sp_7 io_tile_8_0(
            .io_chanxy_in(io_tile_8_0_chanxy_in),
            .io_chanxy_out(io_tile_8_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[192:188]),
            .io_io_input(left_in[63:56]),
            .io_io_output(left_out[63:56]),
            .io_ipin_in(io_tile_8_0_ipin_in),
            .io_opin_out(io_tile_8_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_9_0_chanxy_in;
    wire [29:0] io_tile_9_0_chanxy_out;
    wire [95:0] io_tile_9_0_ipin_in;
    wire [7:0] io_tile_9_0_opin_out;
    io_tile_sp_8 io_tile_9_0(
            .io_chanxy_in(io_tile_9_0_chanxy_in),
            .io_chanxy_out(io_tile_9_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[218:214]),
            .io_io_input(left_in[71:64]),
            .io_io_output(left_out[71:64]),
            .io_ipin_in(io_tile_9_0_ipin_in),
            .io_opin_out(io_tile_9_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [254:0] io_tile_10_0_chanxy_in;
    wire [74:0] io_tile_10_0_chanxy_out;
    wire [95:0] io_tile_10_0_ipin_in;
    wire [7:0] io_tile_10_0_opin_out;
    io_tile_sp_9 io_tile_10_0(
            .io_chanxy_in(io_tile_10_0_chanxy_in),
            .io_chanxy_out(io_tile_10_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[244:240]),
            .io_io_input(left_in[79:72]),
            .io_io_output(left_out[79:72]),
            .io_ipin_in(io_tile_10_0_ipin_in),
            .io_opin_out(io_tile_10_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_1_11_ipin_in;
    wire [7:0] io_tile_1_11_opin_out;
    io_tile_sp_10 io_tile_1_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[5:5]),
            .io_io_input(right_in[7:0]),
            .io_io_output(right_out[7:0]),
            .io_ipin_in(io_tile_1_11_ipin_in),
            .io_opin_out(io_tile_1_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_2_11_ipin_in;
    wire [7:0] io_tile_2_11_opin_out;
    io_tile_sp_11 io_tile_2_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[32:32]),
            .io_io_input(right_in[15:8]),
            .io_io_output(right_out[15:8]),
            .io_ipin_in(io_tile_2_11_ipin_in),
            .io_opin_out(io_tile_2_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_3_11_ipin_in;
    wire [7:0] io_tile_3_11_opin_out;
    io_tile_sp_12 io_tile_3_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[58:58]),
            .io_io_input(right_in[23:16]),
            .io_io_output(right_out[23:16]),
            .io_ipin_in(io_tile_3_11_ipin_in),
            .io_opin_out(io_tile_3_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_4_11_ipin_in;
    wire [7:0] io_tile_4_11_opin_out;
    io_tile_sp_13 io_tile_4_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[84:84]),
            .io_io_input(right_in[31:24]),
            .io_io_output(right_out[31:24]),
            .io_ipin_in(io_tile_4_11_ipin_in),
            .io_opin_out(io_tile_4_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_5_11_ipin_in;
    wire [7:0] io_tile_5_11_opin_out;
    io_tile_sp_14 io_tile_5_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[110:110]),
            .io_io_input(right_in[39:32]),
            .io_io_output(right_out[39:32]),
            .io_ipin_in(io_tile_5_11_ipin_in),
            .io_opin_out(io_tile_5_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_6_11_ipin_in;
    wire [7:0] io_tile_6_11_opin_out;
    io_tile_sp_15 io_tile_6_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[136:136]),
            .io_io_input(right_in[47:40]),
            .io_io_output(right_out[47:40]),
            .io_ipin_in(io_tile_6_11_ipin_in),
            .io_opin_out(io_tile_6_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_7_11_ipin_in;
    wire [7:0] io_tile_7_11_opin_out;
    io_tile_sp_16 io_tile_7_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[162:162]),
            .io_io_input(right_in[55:48]),
            .io_io_output(right_out[55:48]),
            .io_ipin_in(io_tile_7_11_ipin_in),
            .io_opin_out(io_tile_7_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_8_11_ipin_in;
    wire [7:0] io_tile_8_11_opin_out;
    io_tile_sp_17 io_tile_8_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[188:188]),
            .io_io_input(right_in[63:56]),
            .io_io_output(right_out[63:56]),
            .io_ipin_in(io_tile_8_11_ipin_in),
            .io_opin_out(io_tile_8_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_9_11_ipin_in;
    wire [7:0] io_tile_9_11_opin_out;
    io_tile_sp_18 io_tile_9_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[214:214]),
            .io_io_input(right_in[71:64]),
            .io_io_output(right_out[71:64]),
            .io_ipin_in(io_tile_9_11_ipin_in),
            .io_opin_out(io_tile_9_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_10_11_ipin_in;
    wire [7:0] io_tile_10_11_opin_out;
    io_tile_sp_19 io_tile_10_11(
            .io_configs_in(configs_in[383:352]),
            .io_configs_en(configs_en[240:240]),
            .io_io_input(right_in[79:72]),
            .io_io_output(right_out[79:72]),
            .io_ipin_in(io_tile_10_11_ipin_in),
            .io_opin_out(io_tile_10_11_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [254:0] io_tile_0_1_chanxy_in;
    wire [74:0] io_tile_0_1_chanxy_out;
    wire [95:0] io_tile_0_1_ipin_in;
    wire [7:0] io_tile_0_1_opin_out;
    io_tile_sp_20 io_tile_0_1(
            .io_chanxy_in(io_tile_0_1_chanxy_in),
            .io_chanxy_out(io_tile_0_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[7:0]),
            .io_io_output(bot_out[7:0]),
            .io_ipin_in(io_tile_0_1_ipin_in),
            .io_opin_out(io_tile_0_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_2_chanxy_in;
    wire [29:0] io_tile_0_2_chanxy_out;
    wire [95:0] io_tile_0_2_ipin_in;
    wire [7:0] io_tile_0_2_opin_out;
    io_tile_sp_21 io_tile_0_2(
            .io_chanxy_in(io_tile_0_2_chanxy_in),
            .io_chanxy_out(io_tile_0_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[15:8]),
            .io_io_output(bot_out[15:8]),
            .io_ipin_in(io_tile_0_2_ipin_in),
            .io_opin_out(io_tile_0_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_3_chanxy_in;
    wire [29:0] io_tile_0_3_chanxy_out;
    wire [95:0] io_tile_0_3_ipin_in;
    wire [7:0] io_tile_0_3_opin_out;
    io_tile_sp_22 io_tile_0_3(
            .io_chanxy_in(io_tile_0_3_chanxy_in),
            .io_chanxy_out(io_tile_0_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[23:16]),
            .io_io_output(bot_out[23:16]),
            .io_ipin_in(io_tile_0_3_ipin_in),
            .io_opin_out(io_tile_0_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_4_chanxy_in;
    wire [29:0] io_tile_0_4_chanxy_out;
    wire [95:0] io_tile_0_4_ipin_in;
    wire [7:0] io_tile_0_4_opin_out;
    io_tile_sp_23 io_tile_0_4(
            .io_chanxy_in(io_tile_0_4_chanxy_in),
            .io_chanxy_out(io_tile_0_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[31:24]),
            .io_io_output(bot_out[31:24]),
            .io_ipin_in(io_tile_0_4_ipin_in),
            .io_opin_out(io_tile_0_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_5_chanxy_in;
    wire [29:0] io_tile_0_5_chanxy_out;
    wire [95:0] io_tile_0_5_ipin_in;
    wire [7:0] io_tile_0_5_opin_out;
    io_tile_sp_24 io_tile_0_5(
            .io_chanxy_in(io_tile_0_5_chanxy_in),
            .io_chanxy_out(io_tile_0_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[39:32]),
            .io_io_output(bot_out[39:32]),
            .io_ipin_in(io_tile_0_5_ipin_in),
            .io_opin_out(io_tile_0_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_6_chanxy_in;
    wire [29:0] io_tile_0_6_chanxy_out;
    wire [95:0] io_tile_0_6_ipin_in;
    wire [7:0] io_tile_0_6_opin_out;
    io_tile_sp_25 io_tile_0_6(
            .io_chanxy_in(io_tile_0_6_chanxy_in),
            .io_chanxy_out(io_tile_0_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[47:40]),
            .io_io_output(bot_out[47:40]),
            .io_ipin_in(io_tile_0_6_ipin_in),
            .io_opin_out(io_tile_0_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_7_chanxy_in;
    wire [29:0] io_tile_0_7_chanxy_out;
    wire [95:0] io_tile_0_7_ipin_in;
    wire [7:0] io_tile_0_7_opin_out;
    io_tile_sp_26 io_tile_0_7(
            .io_chanxy_in(io_tile_0_7_chanxy_in),
            .io_chanxy_out(io_tile_0_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[55:48]),
            .io_io_output(bot_out[55:48]),
            .io_ipin_in(io_tile_0_7_ipin_in),
            .io_opin_out(io_tile_0_7_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_8_chanxy_in;
    wire [29:0] io_tile_0_8_chanxy_out;
    wire [95:0] io_tile_0_8_ipin_in;
    wire [7:0] io_tile_0_8_opin_out;
    io_tile_sp_27 io_tile_0_8(
            .io_chanxy_in(io_tile_0_8_chanxy_in),
            .io_chanxy_out(io_tile_0_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[63:56]),
            .io_io_output(bot_out[63:56]),
            .io_ipin_in(io_tile_0_8_ipin_in),
            .io_opin_out(io_tile_0_8_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [269:0] io_tile_0_9_chanxy_in;
    wire [29:0] io_tile_0_9_chanxy_out;
    wire [95:0] io_tile_0_9_ipin_in;
    wire [7:0] io_tile_0_9_opin_out;
    io_tile_sp_28 io_tile_0_9(
            .io_chanxy_in(io_tile_0_9_chanxy_in),
            .io_chanxy_out(io_tile_0_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[71:64]),
            .io_io_output(bot_out[71:64]),
            .io_ipin_in(io_tile_0_9_ipin_in),
            .io_opin_out(io_tile_0_9_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [254:0] io_tile_0_10_chanxy_in;
    wire [74:0] io_tile_0_10_chanxy_out;
    wire [95:0] io_tile_0_10_ipin_in;
    wire [7:0] io_tile_0_10_opin_out;
    io_tile_sp_29 io_tile_0_10(
            .io_chanxy_in(io_tile_0_10_chanxy_in),
            .io_chanxy_out(io_tile_0_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[4:0]),
            .io_io_input(bot_in[79:72]),
            .io_io_output(bot_out[79:72]),
            .io_ipin_in(io_tile_0_10_ipin_in),
            .io_opin_out(io_tile_0_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_1_ipin_in;
    wire [7:0] io_tile_11_1_opin_out;
    io_tile_sp_30 io_tile_11_1(
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[7:0]),
            .io_io_output(top_out[7:0]),
            .io_ipin_in(io_tile_11_1_ipin_in),
            .io_opin_out(io_tile_11_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_2_ipin_in;
    wire [7:0] io_tile_11_2_opin_out;
    io_tile_sp_31 io_tile_11_2(
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[15:8]),
            .io_io_output(top_out[15:8]),
            .io_ipin_in(io_tile_11_2_ipin_in),
            .io_opin_out(io_tile_11_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_3_ipin_in;
    wire [7:0] io_tile_11_3_opin_out;
    io_tile_sp_32 io_tile_11_3(
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[23:16]),
            .io_io_output(top_out[23:16]),
            .io_ipin_in(io_tile_11_3_ipin_in),
            .io_opin_out(io_tile_11_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_4_ipin_in;
    wire [7:0] io_tile_11_4_opin_out;
    io_tile_sp_33 io_tile_11_4(
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[31:24]),
            .io_io_output(top_out[31:24]),
            .io_ipin_in(io_tile_11_4_ipin_in),
            .io_opin_out(io_tile_11_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_5_ipin_in;
    wire [7:0] io_tile_11_5_opin_out;
    io_tile_sp_34 io_tile_11_5(
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[39:32]),
            .io_io_output(top_out[39:32]),
            .io_ipin_in(io_tile_11_5_ipin_in),
            .io_opin_out(io_tile_11_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_6_ipin_in;
    wire [7:0] io_tile_11_6_opin_out;
    io_tile_sp_35 io_tile_11_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[47:40]),
            .io_io_output(top_out[47:40]),
            .io_ipin_in(io_tile_11_6_ipin_in),
            .io_opin_out(io_tile_11_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_7_ipin_in;
    wire [7:0] io_tile_11_7_opin_out;
    io_tile_sp_36 io_tile_11_7(
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[55:48]),
            .io_io_output(top_out[55:48]),
            .io_ipin_in(io_tile_11_7_ipin_in),
            .io_opin_out(io_tile_11_7_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_8_ipin_in;
    wire [7:0] io_tile_11_8_opin_out;
    io_tile_sp_37 io_tile_11_8(
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[63:56]),
            .io_io_output(top_out[63:56]),
            .io_ipin_in(io_tile_11_8_ipin_in),
            .io_opin_out(io_tile_11_8_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_9_ipin_in;
    wire [7:0] io_tile_11_9_opin_out;
    io_tile_sp_38 io_tile_11_9(
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[71:64]),
            .io_io_output(top_out[71:64]),
            .io_ipin_in(io_tile_11_9_ipin_in),
            .io_opin_out(io_tile_11_9_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [95:0] io_tile_11_10_ipin_in;
    wire [7:0] io_tile_11_10_opin_out;
    io_tile_sp_39 io_tile_11_10(
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[266:266]),
            .io_io_input(top_in[79:72]),
            .io_io_output(top_out[79:72]),
            .io_ipin_in(io_tile_11_10_ipin_in),
            .io_opin_out(io_tile_11_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );



    // FPGA LUT TILES DECLARE
    wire [605:0] lut_tile_1_1_chanxy_in;
    wire [149:0] lut_tile_1_1_chanxy_out;
    wire [275:0] lut_tile_1_1_ipin_in;
    wire [7:0] lut_tile_1_1_opin_out;
    lut_tile_sp_0 lut_tile_1_1(
            .io_chanxy_in(lut_tile_1_1_chanxy_in),
            .io_chanxy_out(lut_tile_1_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[31:5]),
            .io_ipin_in(lut_tile_1_1_ipin_in),
            .io_opin_out(lut_tile_1_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_2_1_chanxy_in;
    wire [104:0] lut_tile_2_1_chanxy_out;
    wire [275:0] lut_tile_2_1_ipin_in;
    wire [7:0] lut_tile_2_1_opin_out;
    lut_tile_sp_1 lut_tile_2_1(
            .io_chanxy_in(lut_tile_2_1_chanxy_in),
            .io_chanxy_out(lut_tile_2_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[57:32]),
            .io_ipin_in(lut_tile_2_1_ipin_in),
            .io_opin_out(lut_tile_2_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_3_1_chanxy_in;
    wire [104:0] lut_tile_3_1_chanxy_out;
    wire [275:0] lut_tile_3_1_ipin_in;
    wire [7:0] lut_tile_3_1_opin_out;
    lut_tile_sp_2 lut_tile_3_1(
            .io_chanxy_in(lut_tile_3_1_chanxy_in),
            .io_chanxy_out(lut_tile_3_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[83:58]),
            .io_ipin_in(lut_tile_3_1_ipin_in),
            .io_opin_out(lut_tile_3_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_4_1_chanxy_in;
    wire [104:0] lut_tile_4_1_chanxy_out;
    wire [275:0] lut_tile_4_1_ipin_in;
    wire [7:0] lut_tile_4_1_opin_out;
    lut_tile_sp_3 lut_tile_4_1(
            .io_chanxy_in(lut_tile_4_1_chanxy_in),
            .io_chanxy_out(lut_tile_4_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[109:84]),
            .io_ipin_in(lut_tile_4_1_ipin_in),
            .io_opin_out(lut_tile_4_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_5_1_chanxy_in;
    wire [104:0] lut_tile_5_1_chanxy_out;
    wire [275:0] lut_tile_5_1_ipin_in;
    wire [7:0] lut_tile_5_1_opin_out;
    lut_tile_sp_4 lut_tile_5_1(
            .io_chanxy_in(lut_tile_5_1_chanxy_in),
            .io_chanxy_out(lut_tile_5_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[135:110]),
            .io_ipin_in(lut_tile_5_1_ipin_in),
            .io_opin_out(lut_tile_5_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_6_1_chanxy_in;
    wire [104:0] lut_tile_6_1_chanxy_out;
    wire [275:0] lut_tile_6_1_ipin_in;
    wire [7:0] lut_tile_6_1_opin_out;
    lut_tile_sp_5 lut_tile_6_1(
            .io_chanxy_in(lut_tile_6_1_chanxy_in),
            .io_chanxy_out(lut_tile_6_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[161:136]),
            .io_ipin_in(lut_tile_6_1_ipin_in),
            .io_opin_out(lut_tile_6_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_7_1_chanxy_in;
    wire [104:0] lut_tile_7_1_chanxy_out;
    wire [275:0] lut_tile_7_1_ipin_in;
    wire [7:0] lut_tile_7_1_opin_out;
    lut_tile_sp_6 lut_tile_7_1(
            .io_chanxy_in(lut_tile_7_1_chanxy_in),
            .io_chanxy_out(lut_tile_7_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[187:162]),
            .io_ipin_in(lut_tile_7_1_ipin_in),
            .io_opin_out(lut_tile_7_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_8_1_chanxy_in;
    wire [104:0] lut_tile_8_1_chanxy_out;
    wire [275:0] lut_tile_8_1_ipin_in;
    wire [7:0] lut_tile_8_1_opin_out;
    lut_tile_sp_7 lut_tile_8_1(
            .io_chanxy_in(lut_tile_8_1_chanxy_in),
            .io_chanxy_out(lut_tile_8_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[213:188]),
            .io_ipin_in(lut_tile_8_1_ipin_in),
            .io_opin_out(lut_tile_8_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_9_1_chanxy_in;
    wire [104:0] lut_tile_9_1_chanxy_out;
    wire [275:0] lut_tile_9_1_ipin_in;
    wire [7:0] lut_tile_9_1_opin_out;
    lut_tile_sp_8 lut_tile_9_1(
            .io_chanxy_in(lut_tile_9_1_chanxy_in),
            .io_chanxy_out(lut_tile_9_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[239:214]),
            .io_ipin_in(lut_tile_9_1_ipin_in),
            .io_opin_out(lut_tile_9_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [557:0] lut_tile_10_1_chanxy_in;
    wire [149:0] lut_tile_10_1_chanxy_out;
    wire [275:0] lut_tile_10_1_ipin_in;
    wire [7:0] lut_tile_10_1_opin_out;
    lut_tile_sp_9 lut_tile_10_1(
            .io_chanxy_in(lut_tile_10_1_chanxy_in),
            .io_chanxy_out(lut_tile_10_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_1_ipin_in),
            .io_opin_out(lut_tile_10_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [557:0] lut_tile_1_10_chanxy_in;
    wire [149:0] lut_tile_1_10_chanxy_out;
    wire [275:0] lut_tile_1_10_ipin_in;
    wire [7:0] lut_tile_1_10_opin_out;
    lut_tile_sp_10 lut_tile_1_10(
            .io_chanxy_in(lut_tile_1_10_chanxy_in),
            .io_chanxy_out(lut_tile_1_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_10_ipin_in),
            .io_opin_out(lut_tile_1_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_2_10_chanxy_in;
    wire [104:0] lut_tile_2_10_chanxy_out;
    wire [275:0] lut_tile_2_10_ipin_in;
    wire [7:0] lut_tile_2_10_opin_out;
    lut_tile_sp_11 lut_tile_2_10(
            .io_chanxy_in(lut_tile_2_10_chanxy_in),
            .io_chanxy_out(lut_tile_2_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[57:32]),
            .io_ipin_in(lut_tile_2_10_ipin_in),
            .io_opin_out(lut_tile_2_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_3_10_chanxy_in;
    wire [104:0] lut_tile_3_10_chanxy_out;
    wire [275:0] lut_tile_3_10_ipin_in;
    wire [7:0] lut_tile_3_10_opin_out;
    lut_tile_sp_12 lut_tile_3_10(
            .io_chanxy_in(lut_tile_3_10_chanxy_in),
            .io_chanxy_out(lut_tile_3_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[83:58]),
            .io_ipin_in(lut_tile_3_10_ipin_in),
            .io_opin_out(lut_tile_3_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_4_10_chanxy_in;
    wire [104:0] lut_tile_4_10_chanxy_out;
    wire [275:0] lut_tile_4_10_ipin_in;
    wire [7:0] lut_tile_4_10_opin_out;
    lut_tile_sp_13 lut_tile_4_10(
            .io_chanxy_in(lut_tile_4_10_chanxy_in),
            .io_chanxy_out(lut_tile_4_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[109:84]),
            .io_ipin_in(lut_tile_4_10_ipin_in),
            .io_opin_out(lut_tile_4_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_5_10_chanxy_in;
    wire [104:0] lut_tile_5_10_chanxy_out;
    wire [275:0] lut_tile_5_10_ipin_in;
    wire [7:0] lut_tile_5_10_opin_out;
    lut_tile_sp_14 lut_tile_5_10(
            .io_chanxy_in(lut_tile_5_10_chanxy_in),
            .io_chanxy_out(lut_tile_5_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[135:110]),
            .io_ipin_in(lut_tile_5_10_ipin_in),
            .io_opin_out(lut_tile_5_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_6_10_chanxy_in;
    wire [104:0] lut_tile_6_10_chanxy_out;
    wire [275:0] lut_tile_6_10_ipin_in;
    wire [7:0] lut_tile_6_10_opin_out;
    lut_tile_sp_15 lut_tile_6_10(
            .io_chanxy_in(lut_tile_6_10_chanxy_in),
            .io_chanxy_out(lut_tile_6_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[161:136]),
            .io_ipin_in(lut_tile_6_10_ipin_in),
            .io_opin_out(lut_tile_6_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_7_10_chanxy_in;
    wire [104:0] lut_tile_7_10_chanxy_out;
    wire [275:0] lut_tile_7_10_ipin_in;
    wire [7:0] lut_tile_7_10_opin_out;
    lut_tile_sp_16 lut_tile_7_10(
            .io_chanxy_in(lut_tile_7_10_chanxy_in),
            .io_chanxy_out(lut_tile_7_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[187:162]),
            .io_ipin_in(lut_tile_7_10_ipin_in),
            .io_opin_out(lut_tile_7_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_8_10_chanxy_in;
    wire [104:0] lut_tile_8_10_chanxy_out;
    wire [275:0] lut_tile_8_10_ipin_in;
    wire [7:0] lut_tile_8_10_opin_out;
    lut_tile_sp_17 lut_tile_8_10(
            .io_chanxy_in(lut_tile_8_10_chanxy_in),
            .io_chanxy_out(lut_tile_8_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[213:188]),
            .io_ipin_in(lut_tile_8_10_ipin_in),
            .io_opin_out(lut_tile_8_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_9_10_chanxy_in;
    wire [104:0] lut_tile_9_10_chanxy_out;
    wire [275:0] lut_tile_9_10_ipin_in;
    wire [7:0] lut_tile_9_10_opin_out;
    lut_tile_sp_18 lut_tile_9_10(
            .io_chanxy_in(lut_tile_9_10_chanxy_in),
            .io_chanxy_out(lut_tile_9_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[239:214]),
            .io_ipin_in(lut_tile_9_10_ipin_in),
            .io_opin_out(lut_tile_9_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [509:0] lut_tile_10_10_chanxy_in;
    wire [149:0] lut_tile_10_10_chanxy_out;
    wire [275:0] lut_tile_10_10_ipin_in;
    wire [7:0] lut_tile_10_10_opin_out;
    lut_tile_sp_19 lut_tile_10_10(
            .io_chanxy_in(lut_tile_10_10_chanxy_in),
            .io_chanxy_out(lut_tile_10_10_chanxy_out),
            .io_configs_in(configs_in[351:320]),
            .io_configs_en(configs_en[264:240]),
            .io_ipin_in(lut_tile_10_10_ipin_in),
            .io_opin_out(lut_tile_10_10_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_2_chanxy_in;
    wire [104:0] lut_tile_1_2_chanxy_out;
    wire [275:0] lut_tile_1_2_ipin_in;
    wire [7:0] lut_tile_1_2_opin_out;
    lut_tile_sp_20 lut_tile_1_2(
            .io_chanxy_in(lut_tile_1_2_chanxy_in),
            .io_chanxy_out(lut_tile_1_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_2_ipin_in),
            .io_opin_out(lut_tile_1_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_3_chanxy_in;
    wire [104:0] lut_tile_1_3_chanxy_out;
    wire [275:0] lut_tile_1_3_ipin_in;
    wire [7:0] lut_tile_1_3_opin_out;
    lut_tile_sp_21 lut_tile_1_3(
            .io_chanxy_in(lut_tile_1_3_chanxy_in),
            .io_chanxy_out(lut_tile_1_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_3_ipin_in),
            .io_opin_out(lut_tile_1_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_4_chanxy_in;
    wire [104:0] lut_tile_1_4_chanxy_out;
    wire [275:0] lut_tile_1_4_ipin_in;
    wire [7:0] lut_tile_1_4_opin_out;
    lut_tile_sp_22 lut_tile_1_4(
            .io_chanxy_in(lut_tile_1_4_chanxy_in),
            .io_chanxy_out(lut_tile_1_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_4_ipin_in),
            .io_opin_out(lut_tile_1_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_5_chanxy_in;
    wire [104:0] lut_tile_1_5_chanxy_out;
    wire [275:0] lut_tile_1_5_ipin_in;
    wire [7:0] lut_tile_1_5_opin_out;
    lut_tile_sp_23 lut_tile_1_5(
            .io_chanxy_in(lut_tile_1_5_chanxy_in),
            .io_chanxy_out(lut_tile_1_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_5_ipin_in),
            .io_opin_out(lut_tile_1_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_6_chanxy_in;
    wire [104:0] lut_tile_1_6_chanxy_out;
    wire [275:0] lut_tile_1_6_ipin_in;
    wire [7:0] lut_tile_1_6_opin_out;
    lut_tile_sp_24 lut_tile_1_6(
            .io_chanxy_in(lut_tile_1_6_chanxy_in),
            .io_chanxy_out(lut_tile_1_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_6_ipin_in),
            .io_opin_out(lut_tile_1_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_7_chanxy_in;
    wire [104:0] lut_tile_1_7_chanxy_out;
    wire [275:0] lut_tile_1_7_ipin_in;
    wire [7:0] lut_tile_1_7_opin_out;
    lut_tile_sp_25 lut_tile_1_7(
            .io_chanxy_in(lut_tile_1_7_chanxy_in),
            .io_chanxy_out(lut_tile_1_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_7_ipin_in),
            .io_opin_out(lut_tile_1_7_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_8_chanxy_in;
    wire [104:0] lut_tile_1_8_chanxy_out;
    wire [275:0] lut_tile_1_8_ipin_in;
    wire [7:0] lut_tile_1_8_opin_out;
    lut_tile_sp_26 lut_tile_1_8(
            .io_chanxy_in(lut_tile_1_8_chanxy_in),
            .io_chanxy_out(lut_tile_1_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_8_ipin_in),
            .io_opin_out(lut_tile_1_8_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [620:0] lut_tile_1_9_chanxy_in;
    wire [104:0] lut_tile_1_9_chanxy_out;
    wire [275:0] lut_tile_1_9_ipin_in;
    wire [7:0] lut_tile_1_9_opin_out;
    lut_tile_sp_27 lut_tile_1_9(
            .io_chanxy_in(lut_tile_1_9_chanxy_in),
            .io_chanxy_out(lut_tile_1_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[30:5]),
            .io_ipin_in(lut_tile_1_9_ipin_in),
            .io_opin_out(lut_tile_1_9_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_2_chanxy_in;
    wire [104:0] lut_tile_10_2_chanxy_out;
    wire [275:0] lut_tile_10_2_ipin_in;
    wire [7:0] lut_tile_10_2_opin_out;
    lut_tile_sp_28 lut_tile_10_2(
            .io_chanxy_in(lut_tile_10_2_chanxy_in),
            .io_chanxy_out(lut_tile_10_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_2_ipin_in),
            .io_opin_out(lut_tile_10_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_3_chanxy_in;
    wire [104:0] lut_tile_10_3_chanxy_out;
    wire [275:0] lut_tile_10_3_ipin_in;
    wire [7:0] lut_tile_10_3_opin_out;
    lut_tile_sp_29 lut_tile_10_3(
            .io_chanxy_in(lut_tile_10_3_chanxy_in),
            .io_chanxy_out(lut_tile_10_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_3_ipin_in),
            .io_opin_out(lut_tile_10_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_4_chanxy_in;
    wire [104:0] lut_tile_10_4_chanxy_out;
    wire [275:0] lut_tile_10_4_ipin_in;
    wire [7:0] lut_tile_10_4_opin_out;
    lut_tile_sp_30 lut_tile_10_4(
            .io_chanxy_in(lut_tile_10_4_chanxy_in),
            .io_chanxy_out(lut_tile_10_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_4_ipin_in),
            .io_opin_out(lut_tile_10_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_5_chanxy_in;
    wire [104:0] lut_tile_10_5_chanxy_out;
    wire [275:0] lut_tile_10_5_ipin_in;
    wire [7:0] lut_tile_10_5_opin_out;
    lut_tile_sp_31 lut_tile_10_5(
            .io_chanxy_in(lut_tile_10_5_chanxy_in),
            .io_chanxy_out(lut_tile_10_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_5_ipin_in),
            .io_opin_out(lut_tile_10_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_6_chanxy_in;
    wire [104:0] lut_tile_10_6_chanxy_out;
    wire [275:0] lut_tile_10_6_ipin_in;
    wire [7:0] lut_tile_10_6_opin_out;
    lut_tile_sp_32 lut_tile_10_6(
            .io_chanxy_in(lut_tile_10_6_chanxy_in),
            .io_chanxy_out(lut_tile_10_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_6_ipin_in),
            .io_opin_out(lut_tile_10_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_7_chanxy_in;
    wire [104:0] lut_tile_10_7_chanxy_out;
    wire [275:0] lut_tile_10_7_ipin_in;
    wire [7:0] lut_tile_10_7_opin_out;
    lut_tile_sp_33 lut_tile_10_7(
            .io_chanxy_in(lut_tile_10_7_chanxy_in),
            .io_chanxy_out(lut_tile_10_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_7_ipin_in),
            .io_opin_out(lut_tile_10_7_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_8_chanxy_in;
    wire [104:0] lut_tile_10_8_chanxy_out;
    wire [275:0] lut_tile_10_8_ipin_in;
    wire [7:0] lut_tile_10_8_opin_out;
    lut_tile_sp_34 lut_tile_10_8(
            .io_chanxy_in(lut_tile_10_8_chanxy_in),
            .io_chanxy_out(lut_tile_10_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_8_ipin_in),
            .io_opin_out(lut_tile_10_8_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [572:0] lut_tile_10_9_chanxy_in;
    wire [104:0] lut_tile_10_9_chanxy_out;
    wire [275:0] lut_tile_10_9_ipin_in;
    wire [7:0] lut_tile_10_9_opin_out;
    lut_tile_sp_35 lut_tile_10_9(
            .io_chanxy_in(lut_tile_10_9_chanxy_in),
            .io_chanxy_out(lut_tile_10_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[265:240]),
            .io_ipin_in(lut_tile_10_9_ipin_in),
            .io_opin_out(lut_tile_10_9_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_2_chanxy_in;
    wire [59:0] lut_tile_2_2_chanxy_out;
    wire [275:0] lut_tile_2_2_ipin_in;
    wire [7:0] lut_tile_2_2_opin_out;
    lut_tile lut_tile_2_2(
            .io_chanxy_in(lut_tile_2_2_chanxy_in),
            .io_chanxy_out(lut_tile_2_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_2_ipin_in),
            .io_opin_out(lut_tile_2_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_3_chanxy_in;
    wire [59:0] lut_tile_2_3_chanxy_out;
    wire [275:0] lut_tile_2_3_ipin_in;
    wire [7:0] lut_tile_2_3_opin_out;
    lut_tile lut_tile_2_3(
            .io_chanxy_in(lut_tile_2_3_chanxy_in),
            .io_chanxy_out(lut_tile_2_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_3_ipin_in),
            .io_opin_out(lut_tile_2_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_4_chanxy_in;
    wire [59:0] lut_tile_2_4_chanxy_out;
    wire [275:0] lut_tile_2_4_ipin_in;
    wire [7:0] lut_tile_2_4_opin_out;
    lut_tile lut_tile_2_4(
            .io_chanxy_in(lut_tile_2_4_chanxy_in),
            .io_chanxy_out(lut_tile_2_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_4_ipin_in),
            .io_opin_out(lut_tile_2_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_5_chanxy_in;
    wire [59:0] lut_tile_2_5_chanxy_out;
    wire [275:0] lut_tile_2_5_ipin_in;
    wire [7:0] lut_tile_2_5_opin_out;
    lut_tile lut_tile_2_5(
            .io_chanxy_in(lut_tile_2_5_chanxy_in),
            .io_chanxy_out(lut_tile_2_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_5_ipin_in),
            .io_opin_out(lut_tile_2_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_6_chanxy_in;
    wire [59:0] lut_tile_2_6_chanxy_out;
    wire [275:0] lut_tile_2_6_ipin_in;
    wire [7:0] lut_tile_2_6_opin_out;
    lut_tile lut_tile_2_6(
            .io_chanxy_in(lut_tile_2_6_chanxy_in),
            .io_chanxy_out(lut_tile_2_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_6_ipin_in),
            .io_opin_out(lut_tile_2_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_7_chanxy_in;
    wire [59:0] lut_tile_2_7_chanxy_out;
    wire [275:0] lut_tile_2_7_ipin_in;
    wire [7:0] lut_tile_2_7_opin_out;
    lut_tile lut_tile_2_7(
            .io_chanxy_in(lut_tile_2_7_chanxy_in),
            .io_chanxy_out(lut_tile_2_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_7_ipin_in),
            .io_opin_out(lut_tile_2_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_8_chanxy_in;
    wire [59:0] lut_tile_2_8_chanxy_out;
    wire [275:0] lut_tile_2_8_ipin_in;
    wire [7:0] lut_tile_2_8_opin_out;
    lut_tile lut_tile_2_8(
            .io_chanxy_in(lut_tile_2_8_chanxy_in),
            .io_chanxy_out(lut_tile_2_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_8_ipin_in),
            .io_opin_out(lut_tile_2_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_2_9_chanxy_in;
    wire [59:0] lut_tile_2_9_chanxy_out;
    wire [275:0] lut_tile_2_9_ipin_in;
    wire [7:0] lut_tile_2_9_opin_out;
    lut_tile lut_tile_2_9(
            .io_chanxy_in(lut_tile_2_9_chanxy_in),
            .io_chanxy_out(lut_tile_2_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[56:32]),
            .io_ipin_in(lut_tile_2_9_ipin_in),
            .io_opin_out(lut_tile_2_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_2_chanxy_in;
    wire [59:0] lut_tile_3_2_chanxy_out;
    wire [275:0] lut_tile_3_2_ipin_in;
    wire [7:0] lut_tile_3_2_opin_out;
    lut_tile lut_tile_3_2(
            .io_chanxy_in(lut_tile_3_2_chanxy_in),
            .io_chanxy_out(lut_tile_3_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_2_ipin_in),
            .io_opin_out(lut_tile_3_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_3_chanxy_in;
    wire [59:0] lut_tile_3_3_chanxy_out;
    wire [275:0] lut_tile_3_3_ipin_in;
    wire [7:0] lut_tile_3_3_opin_out;
    lut_tile lut_tile_3_3(
            .io_chanxy_in(lut_tile_3_3_chanxy_in),
            .io_chanxy_out(lut_tile_3_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_3_ipin_in),
            .io_opin_out(lut_tile_3_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_4_chanxy_in;
    wire [59:0] lut_tile_3_4_chanxy_out;
    wire [275:0] lut_tile_3_4_ipin_in;
    wire [7:0] lut_tile_3_4_opin_out;
    lut_tile lut_tile_3_4(
            .io_chanxy_in(lut_tile_3_4_chanxy_in),
            .io_chanxy_out(lut_tile_3_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_4_ipin_in),
            .io_opin_out(lut_tile_3_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_5_chanxy_in;
    wire [59:0] lut_tile_3_5_chanxy_out;
    wire [275:0] lut_tile_3_5_ipin_in;
    wire [7:0] lut_tile_3_5_opin_out;
    lut_tile lut_tile_3_5(
            .io_chanxy_in(lut_tile_3_5_chanxy_in),
            .io_chanxy_out(lut_tile_3_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_5_ipin_in),
            .io_opin_out(lut_tile_3_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_6_chanxy_in;
    wire [59:0] lut_tile_3_6_chanxy_out;
    wire [275:0] lut_tile_3_6_ipin_in;
    wire [7:0] lut_tile_3_6_opin_out;
    lut_tile lut_tile_3_6(
            .io_chanxy_in(lut_tile_3_6_chanxy_in),
            .io_chanxy_out(lut_tile_3_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_6_ipin_in),
            .io_opin_out(lut_tile_3_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_7_chanxy_in;
    wire [59:0] lut_tile_3_7_chanxy_out;
    wire [275:0] lut_tile_3_7_ipin_in;
    wire [7:0] lut_tile_3_7_opin_out;
    lut_tile lut_tile_3_7(
            .io_chanxy_in(lut_tile_3_7_chanxy_in),
            .io_chanxy_out(lut_tile_3_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_7_ipin_in),
            .io_opin_out(lut_tile_3_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_8_chanxy_in;
    wire [59:0] lut_tile_3_8_chanxy_out;
    wire [275:0] lut_tile_3_8_ipin_in;
    wire [7:0] lut_tile_3_8_opin_out;
    lut_tile lut_tile_3_8(
            .io_chanxy_in(lut_tile_3_8_chanxy_in),
            .io_chanxy_out(lut_tile_3_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_8_ipin_in),
            .io_opin_out(lut_tile_3_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_3_9_chanxy_in;
    wire [59:0] lut_tile_3_9_chanxy_out;
    wire [275:0] lut_tile_3_9_ipin_in;
    wire [7:0] lut_tile_3_9_opin_out;
    lut_tile lut_tile_3_9(
            .io_chanxy_in(lut_tile_3_9_chanxy_in),
            .io_chanxy_out(lut_tile_3_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[82:58]),
            .io_ipin_in(lut_tile_3_9_ipin_in),
            .io_opin_out(lut_tile_3_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_2_chanxy_in;
    wire [59:0] lut_tile_4_2_chanxy_out;
    wire [275:0] lut_tile_4_2_ipin_in;
    wire [7:0] lut_tile_4_2_opin_out;
    lut_tile lut_tile_4_2(
            .io_chanxy_in(lut_tile_4_2_chanxy_in),
            .io_chanxy_out(lut_tile_4_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_2_ipin_in),
            .io_opin_out(lut_tile_4_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_3_chanxy_in;
    wire [59:0] lut_tile_4_3_chanxy_out;
    wire [275:0] lut_tile_4_3_ipin_in;
    wire [7:0] lut_tile_4_3_opin_out;
    lut_tile lut_tile_4_3(
            .io_chanxy_in(lut_tile_4_3_chanxy_in),
            .io_chanxy_out(lut_tile_4_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_3_ipin_in),
            .io_opin_out(lut_tile_4_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_4_chanxy_in;
    wire [59:0] lut_tile_4_4_chanxy_out;
    wire [275:0] lut_tile_4_4_ipin_in;
    wire [7:0] lut_tile_4_4_opin_out;
    lut_tile lut_tile_4_4(
            .io_chanxy_in(lut_tile_4_4_chanxy_in),
            .io_chanxy_out(lut_tile_4_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_4_ipin_in),
            .io_opin_out(lut_tile_4_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_5_chanxy_in;
    wire [59:0] lut_tile_4_5_chanxy_out;
    wire [275:0] lut_tile_4_5_ipin_in;
    wire [7:0] lut_tile_4_5_opin_out;
    lut_tile lut_tile_4_5(
            .io_chanxy_in(lut_tile_4_5_chanxy_in),
            .io_chanxy_out(lut_tile_4_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_5_ipin_in),
            .io_opin_out(lut_tile_4_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_6_chanxy_in;
    wire [59:0] lut_tile_4_6_chanxy_out;
    wire [275:0] lut_tile_4_6_ipin_in;
    wire [7:0] lut_tile_4_6_opin_out;
    lut_tile lut_tile_4_6(
            .io_chanxy_in(lut_tile_4_6_chanxy_in),
            .io_chanxy_out(lut_tile_4_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_6_ipin_in),
            .io_opin_out(lut_tile_4_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_7_chanxy_in;
    wire [59:0] lut_tile_4_7_chanxy_out;
    wire [275:0] lut_tile_4_7_ipin_in;
    wire [7:0] lut_tile_4_7_opin_out;
    lut_tile lut_tile_4_7(
            .io_chanxy_in(lut_tile_4_7_chanxy_in),
            .io_chanxy_out(lut_tile_4_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_7_ipin_in),
            .io_opin_out(lut_tile_4_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_8_chanxy_in;
    wire [59:0] lut_tile_4_8_chanxy_out;
    wire [275:0] lut_tile_4_8_ipin_in;
    wire [7:0] lut_tile_4_8_opin_out;
    lut_tile lut_tile_4_8(
            .io_chanxy_in(lut_tile_4_8_chanxy_in),
            .io_chanxy_out(lut_tile_4_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_8_ipin_in),
            .io_opin_out(lut_tile_4_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_4_9_chanxy_in;
    wire [59:0] lut_tile_4_9_chanxy_out;
    wire [275:0] lut_tile_4_9_ipin_in;
    wire [7:0] lut_tile_4_9_opin_out;
    lut_tile lut_tile_4_9(
            .io_chanxy_in(lut_tile_4_9_chanxy_in),
            .io_chanxy_out(lut_tile_4_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[108:84]),
            .io_ipin_in(lut_tile_4_9_ipin_in),
            .io_opin_out(lut_tile_4_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_2_chanxy_in;
    wire [59:0] lut_tile_5_2_chanxy_out;
    wire [275:0] lut_tile_5_2_ipin_in;
    wire [7:0] lut_tile_5_2_opin_out;
    lut_tile lut_tile_5_2(
            .io_chanxy_in(lut_tile_5_2_chanxy_in),
            .io_chanxy_out(lut_tile_5_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_2_ipin_in),
            .io_opin_out(lut_tile_5_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_3_chanxy_in;
    wire [59:0] lut_tile_5_3_chanxy_out;
    wire [275:0] lut_tile_5_3_ipin_in;
    wire [7:0] lut_tile_5_3_opin_out;
    lut_tile lut_tile_5_3(
            .io_chanxy_in(lut_tile_5_3_chanxy_in),
            .io_chanxy_out(lut_tile_5_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_3_ipin_in),
            .io_opin_out(lut_tile_5_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_4_chanxy_in;
    wire [59:0] lut_tile_5_4_chanxy_out;
    wire [275:0] lut_tile_5_4_ipin_in;
    wire [7:0] lut_tile_5_4_opin_out;
    lut_tile lut_tile_5_4(
            .io_chanxy_in(lut_tile_5_4_chanxy_in),
            .io_chanxy_out(lut_tile_5_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_4_ipin_in),
            .io_opin_out(lut_tile_5_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_5_chanxy_in;
    wire [59:0] lut_tile_5_5_chanxy_out;
    wire [275:0] lut_tile_5_5_ipin_in;
    wire [7:0] lut_tile_5_5_opin_out;
    lut_tile lut_tile_5_5(
            .io_chanxy_in(lut_tile_5_5_chanxy_in),
            .io_chanxy_out(lut_tile_5_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_5_ipin_in),
            .io_opin_out(lut_tile_5_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_6_chanxy_in;
    wire [59:0] lut_tile_5_6_chanxy_out;
    wire [275:0] lut_tile_5_6_ipin_in;
    wire [7:0] lut_tile_5_6_opin_out;
    lut_tile lut_tile_5_6(
            .io_chanxy_in(lut_tile_5_6_chanxy_in),
            .io_chanxy_out(lut_tile_5_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_6_ipin_in),
            .io_opin_out(lut_tile_5_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_7_chanxy_in;
    wire [59:0] lut_tile_5_7_chanxy_out;
    wire [275:0] lut_tile_5_7_ipin_in;
    wire [7:0] lut_tile_5_7_opin_out;
    lut_tile lut_tile_5_7(
            .io_chanxy_in(lut_tile_5_7_chanxy_in),
            .io_chanxy_out(lut_tile_5_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_7_ipin_in),
            .io_opin_out(lut_tile_5_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_8_chanxy_in;
    wire [59:0] lut_tile_5_8_chanxy_out;
    wire [275:0] lut_tile_5_8_ipin_in;
    wire [7:0] lut_tile_5_8_opin_out;
    lut_tile lut_tile_5_8(
            .io_chanxy_in(lut_tile_5_8_chanxy_in),
            .io_chanxy_out(lut_tile_5_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_8_ipin_in),
            .io_opin_out(lut_tile_5_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_5_9_chanxy_in;
    wire [59:0] lut_tile_5_9_chanxy_out;
    wire [275:0] lut_tile_5_9_ipin_in;
    wire [7:0] lut_tile_5_9_opin_out;
    lut_tile lut_tile_5_9(
            .io_chanxy_in(lut_tile_5_9_chanxy_in),
            .io_chanxy_out(lut_tile_5_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[134:110]),
            .io_ipin_in(lut_tile_5_9_ipin_in),
            .io_opin_out(lut_tile_5_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_2_chanxy_in;
    wire [59:0] lut_tile_6_2_chanxy_out;
    wire [275:0] lut_tile_6_2_ipin_in;
    wire [7:0] lut_tile_6_2_opin_out;
    lut_tile lut_tile_6_2(
            .io_chanxy_in(lut_tile_6_2_chanxy_in),
            .io_chanxy_out(lut_tile_6_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_2_ipin_in),
            .io_opin_out(lut_tile_6_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_3_chanxy_in;
    wire [59:0] lut_tile_6_3_chanxy_out;
    wire [275:0] lut_tile_6_3_ipin_in;
    wire [7:0] lut_tile_6_3_opin_out;
    lut_tile lut_tile_6_3(
            .io_chanxy_in(lut_tile_6_3_chanxy_in),
            .io_chanxy_out(lut_tile_6_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_3_ipin_in),
            .io_opin_out(lut_tile_6_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_4_chanxy_in;
    wire [59:0] lut_tile_6_4_chanxy_out;
    wire [275:0] lut_tile_6_4_ipin_in;
    wire [7:0] lut_tile_6_4_opin_out;
    lut_tile lut_tile_6_4(
            .io_chanxy_in(lut_tile_6_4_chanxy_in),
            .io_chanxy_out(lut_tile_6_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_4_ipin_in),
            .io_opin_out(lut_tile_6_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_5_chanxy_in;
    wire [59:0] lut_tile_6_5_chanxy_out;
    wire [275:0] lut_tile_6_5_ipin_in;
    wire [7:0] lut_tile_6_5_opin_out;
    lut_tile lut_tile_6_5(
            .io_chanxy_in(lut_tile_6_5_chanxy_in),
            .io_chanxy_out(lut_tile_6_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_5_ipin_in),
            .io_opin_out(lut_tile_6_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_6_chanxy_in;
    wire [59:0] lut_tile_6_6_chanxy_out;
    wire [275:0] lut_tile_6_6_ipin_in;
    wire [7:0] lut_tile_6_6_opin_out;
    lut_tile lut_tile_6_6(
            .io_chanxy_in(lut_tile_6_6_chanxy_in),
            .io_chanxy_out(lut_tile_6_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_6_ipin_in),
            .io_opin_out(lut_tile_6_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_7_chanxy_in;
    wire [59:0] lut_tile_6_7_chanxy_out;
    wire [275:0] lut_tile_6_7_ipin_in;
    wire [7:0] lut_tile_6_7_opin_out;
    lut_tile lut_tile_6_7(
            .io_chanxy_in(lut_tile_6_7_chanxy_in),
            .io_chanxy_out(lut_tile_6_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_7_ipin_in),
            .io_opin_out(lut_tile_6_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_8_chanxy_in;
    wire [59:0] lut_tile_6_8_chanxy_out;
    wire [275:0] lut_tile_6_8_ipin_in;
    wire [7:0] lut_tile_6_8_opin_out;
    lut_tile lut_tile_6_8(
            .io_chanxy_in(lut_tile_6_8_chanxy_in),
            .io_chanxy_out(lut_tile_6_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_8_ipin_in),
            .io_opin_out(lut_tile_6_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_6_9_chanxy_in;
    wire [59:0] lut_tile_6_9_chanxy_out;
    wire [275:0] lut_tile_6_9_ipin_in;
    wire [7:0] lut_tile_6_9_opin_out;
    lut_tile lut_tile_6_9(
            .io_chanxy_in(lut_tile_6_9_chanxy_in),
            .io_chanxy_out(lut_tile_6_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[160:136]),
            .io_ipin_in(lut_tile_6_9_ipin_in),
            .io_opin_out(lut_tile_6_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_2_chanxy_in;
    wire [59:0] lut_tile_7_2_chanxy_out;
    wire [275:0] lut_tile_7_2_ipin_in;
    wire [7:0] lut_tile_7_2_opin_out;
    lut_tile lut_tile_7_2(
            .io_chanxy_in(lut_tile_7_2_chanxy_in),
            .io_chanxy_out(lut_tile_7_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_2_ipin_in),
            .io_opin_out(lut_tile_7_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_3_chanxy_in;
    wire [59:0] lut_tile_7_3_chanxy_out;
    wire [275:0] lut_tile_7_3_ipin_in;
    wire [7:0] lut_tile_7_3_opin_out;
    lut_tile lut_tile_7_3(
            .io_chanxy_in(lut_tile_7_3_chanxy_in),
            .io_chanxy_out(lut_tile_7_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_3_ipin_in),
            .io_opin_out(lut_tile_7_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_4_chanxy_in;
    wire [59:0] lut_tile_7_4_chanxy_out;
    wire [275:0] lut_tile_7_4_ipin_in;
    wire [7:0] lut_tile_7_4_opin_out;
    lut_tile lut_tile_7_4(
            .io_chanxy_in(lut_tile_7_4_chanxy_in),
            .io_chanxy_out(lut_tile_7_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_4_ipin_in),
            .io_opin_out(lut_tile_7_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_5_chanxy_in;
    wire [59:0] lut_tile_7_5_chanxy_out;
    wire [275:0] lut_tile_7_5_ipin_in;
    wire [7:0] lut_tile_7_5_opin_out;
    lut_tile lut_tile_7_5(
            .io_chanxy_in(lut_tile_7_5_chanxy_in),
            .io_chanxy_out(lut_tile_7_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_5_ipin_in),
            .io_opin_out(lut_tile_7_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_6_chanxy_in;
    wire [59:0] lut_tile_7_6_chanxy_out;
    wire [275:0] lut_tile_7_6_ipin_in;
    wire [7:0] lut_tile_7_6_opin_out;
    lut_tile lut_tile_7_6(
            .io_chanxy_in(lut_tile_7_6_chanxy_in),
            .io_chanxy_out(lut_tile_7_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_6_ipin_in),
            .io_opin_out(lut_tile_7_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_7_chanxy_in;
    wire [59:0] lut_tile_7_7_chanxy_out;
    wire [275:0] lut_tile_7_7_ipin_in;
    wire [7:0] lut_tile_7_7_opin_out;
    lut_tile lut_tile_7_7(
            .io_chanxy_in(lut_tile_7_7_chanxy_in),
            .io_chanxy_out(lut_tile_7_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_7_ipin_in),
            .io_opin_out(lut_tile_7_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_8_chanxy_in;
    wire [59:0] lut_tile_7_8_chanxy_out;
    wire [275:0] lut_tile_7_8_ipin_in;
    wire [7:0] lut_tile_7_8_opin_out;
    lut_tile lut_tile_7_8(
            .io_chanxy_in(lut_tile_7_8_chanxy_in),
            .io_chanxy_out(lut_tile_7_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_8_ipin_in),
            .io_opin_out(lut_tile_7_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_7_9_chanxy_in;
    wire [59:0] lut_tile_7_9_chanxy_out;
    wire [275:0] lut_tile_7_9_ipin_in;
    wire [7:0] lut_tile_7_9_opin_out;
    lut_tile lut_tile_7_9(
            .io_chanxy_in(lut_tile_7_9_chanxy_in),
            .io_chanxy_out(lut_tile_7_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[186:162]),
            .io_ipin_in(lut_tile_7_9_ipin_in),
            .io_opin_out(lut_tile_7_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_2_chanxy_in;
    wire [59:0] lut_tile_8_2_chanxy_out;
    wire [275:0] lut_tile_8_2_ipin_in;
    wire [7:0] lut_tile_8_2_opin_out;
    lut_tile lut_tile_8_2(
            .io_chanxy_in(lut_tile_8_2_chanxy_in),
            .io_chanxy_out(lut_tile_8_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_2_ipin_in),
            .io_opin_out(lut_tile_8_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_3_chanxy_in;
    wire [59:0] lut_tile_8_3_chanxy_out;
    wire [275:0] lut_tile_8_3_ipin_in;
    wire [7:0] lut_tile_8_3_opin_out;
    lut_tile lut_tile_8_3(
            .io_chanxy_in(lut_tile_8_3_chanxy_in),
            .io_chanxy_out(lut_tile_8_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_3_ipin_in),
            .io_opin_out(lut_tile_8_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_4_chanxy_in;
    wire [59:0] lut_tile_8_4_chanxy_out;
    wire [275:0] lut_tile_8_4_ipin_in;
    wire [7:0] lut_tile_8_4_opin_out;
    lut_tile lut_tile_8_4(
            .io_chanxy_in(lut_tile_8_4_chanxy_in),
            .io_chanxy_out(lut_tile_8_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_4_ipin_in),
            .io_opin_out(lut_tile_8_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_5_chanxy_in;
    wire [59:0] lut_tile_8_5_chanxy_out;
    wire [275:0] lut_tile_8_5_ipin_in;
    wire [7:0] lut_tile_8_5_opin_out;
    lut_tile lut_tile_8_5(
            .io_chanxy_in(lut_tile_8_5_chanxy_in),
            .io_chanxy_out(lut_tile_8_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_5_ipin_in),
            .io_opin_out(lut_tile_8_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_6_chanxy_in;
    wire [59:0] lut_tile_8_6_chanxy_out;
    wire [275:0] lut_tile_8_6_ipin_in;
    wire [7:0] lut_tile_8_6_opin_out;
    lut_tile lut_tile_8_6(
            .io_chanxy_in(lut_tile_8_6_chanxy_in),
            .io_chanxy_out(lut_tile_8_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_6_ipin_in),
            .io_opin_out(lut_tile_8_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_7_chanxy_in;
    wire [59:0] lut_tile_8_7_chanxy_out;
    wire [275:0] lut_tile_8_7_ipin_in;
    wire [7:0] lut_tile_8_7_opin_out;
    lut_tile lut_tile_8_7(
            .io_chanxy_in(lut_tile_8_7_chanxy_in),
            .io_chanxy_out(lut_tile_8_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_7_ipin_in),
            .io_opin_out(lut_tile_8_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_8_chanxy_in;
    wire [59:0] lut_tile_8_8_chanxy_out;
    wire [275:0] lut_tile_8_8_ipin_in;
    wire [7:0] lut_tile_8_8_opin_out;
    lut_tile lut_tile_8_8(
            .io_chanxy_in(lut_tile_8_8_chanxy_in),
            .io_chanxy_out(lut_tile_8_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_8_ipin_in),
            .io_opin_out(lut_tile_8_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_8_9_chanxy_in;
    wire [59:0] lut_tile_8_9_chanxy_out;
    wire [275:0] lut_tile_8_9_ipin_in;
    wire [7:0] lut_tile_8_9_opin_out;
    lut_tile lut_tile_8_9(
            .io_chanxy_in(lut_tile_8_9_chanxy_in),
            .io_chanxy_out(lut_tile_8_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[212:188]),
            .io_ipin_in(lut_tile_8_9_ipin_in),
            .io_opin_out(lut_tile_8_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_2_chanxy_in;
    wire [59:0] lut_tile_9_2_chanxy_out;
    wire [275:0] lut_tile_9_2_ipin_in;
    wire [7:0] lut_tile_9_2_opin_out;
    lut_tile lut_tile_9_2(
            .io_chanxy_in(lut_tile_9_2_chanxy_in),
            .io_chanxy_out(lut_tile_9_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_2_ipin_in),
            .io_opin_out(lut_tile_9_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_3_chanxy_in;
    wire [59:0] lut_tile_9_3_chanxy_out;
    wire [275:0] lut_tile_9_3_ipin_in;
    wire [7:0] lut_tile_9_3_opin_out;
    lut_tile lut_tile_9_3(
            .io_chanxy_in(lut_tile_9_3_chanxy_in),
            .io_chanxy_out(lut_tile_9_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_3_ipin_in),
            .io_opin_out(lut_tile_9_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_4_chanxy_in;
    wire [59:0] lut_tile_9_4_chanxy_out;
    wire [275:0] lut_tile_9_4_ipin_in;
    wire [7:0] lut_tile_9_4_opin_out;
    lut_tile lut_tile_9_4(
            .io_chanxy_in(lut_tile_9_4_chanxy_in),
            .io_chanxy_out(lut_tile_9_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_4_ipin_in),
            .io_opin_out(lut_tile_9_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_5_chanxy_in;
    wire [59:0] lut_tile_9_5_chanxy_out;
    wire [275:0] lut_tile_9_5_ipin_in;
    wire [7:0] lut_tile_9_5_opin_out;
    lut_tile lut_tile_9_5(
            .io_chanxy_in(lut_tile_9_5_chanxy_in),
            .io_chanxy_out(lut_tile_9_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_5_ipin_in),
            .io_opin_out(lut_tile_9_5_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_6_chanxy_in;
    wire [59:0] lut_tile_9_6_chanxy_out;
    wire [275:0] lut_tile_9_6_ipin_in;
    wire [7:0] lut_tile_9_6_opin_out;
    lut_tile lut_tile_9_6(
            .io_chanxy_in(lut_tile_9_6_chanxy_in),
            .io_chanxy_out(lut_tile_9_6_chanxy_out),
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_6_ipin_in),
            .io_opin_out(lut_tile_9_6_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_7_chanxy_in;
    wire [59:0] lut_tile_9_7_chanxy_out;
    wire [275:0] lut_tile_9_7_ipin_in;
    wire [7:0] lut_tile_9_7_opin_out;
    lut_tile lut_tile_9_7(
            .io_chanxy_in(lut_tile_9_7_chanxy_in),
            .io_chanxy_out(lut_tile_9_7_chanxy_out),
            .io_configs_in(configs_in[255:224]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_7_ipin_in),
            .io_opin_out(lut_tile_9_7_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_8_chanxy_in;
    wire [59:0] lut_tile_9_8_chanxy_out;
    wire [275:0] lut_tile_9_8_ipin_in;
    wire [7:0] lut_tile_9_8_opin_out;
    lut_tile lut_tile_9_8(
            .io_chanxy_in(lut_tile_9_8_chanxy_in),
            .io_chanxy_out(lut_tile_9_8_chanxy_out),
            .io_configs_in(configs_in[287:256]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_8_ipin_in),
            .io_opin_out(lut_tile_9_8_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [635:0] lut_tile_9_9_chanxy_in;
    wire [59:0] lut_tile_9_9_chanxy_out;
    wire [275:0] lut_tile_9_9_ipin_in;
    wire [7:0] lut_tile_9_9_opin_out;
    lut_tile lut_tile_9_9(
            .io_chanxy_in(lut_tile_9_9_chanxy_in),
            .io_chanxy_out(lut_tile_9_9_chanxy_out),
            .io_configs_in(configs_in[319:288]),
            .io_configs_en(configs_en[238:214]),
            .io_ipin_in(lut_tile_9_9_ipin_in),
            .io_opin_out(lut_tile_9_9_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );



    // LUT TILE IPIN
    assign lut_tile_1_1_ipin_in = {wire_6239, wire_6238, wire_6219, wire_6218, wire_6199, wire_6198, wire_6179, wire_6178, wire_6159, wire_6158, wire_6139, wire_6138, wire_10917, wire_10916, wire_10897, wire_10896, wire_10877, wire_10876, wire_10857, wire_10856, wire_10837, wire_10836, wire_10817, wire_10816, wire_6625, wire_6624, wire_6613, wire_6612, wire_6585, wire_6584, wire_6573, wire_6572, wire_6545, wire_6544, wire_6533, wire_6532, wire_10527, wire_10526, wire_10507, wire_10506, wire_10487, wire_10486, wire_10467, wire_10466, wire_10447, wire_10446, wire_10427, wire_10426, wire_6235, wire_6234, wire_6215, wire_6214, wire_6195, wire_6194, wire_6175, wire_6174, wire_6155, wire_6154, wire_6135, wire_6134, wire_10913, wire_10912, wire_10893, wire_10892, wire_10873, wire_10872, wire_10853, wire_10852, wire_10833, wire_10832, wire_10813, wire_10812, wire_6629, wire_6628, wire_6601, wire_6600, wire_6589, wire_6588, wire_6561, wire_6560, wire_6549, wire_6548, wire_6521, wire_6520, wire_10523, wire_10522, wire_10503, wire_10502, wire_10483, wire_10482, wire_10463, wire_10462, wire_10443, wire_10442, wire_10423, wire_10422, wire_6233, wire_6232, wire_6213, wire_6212, wire_6193, wire_6192, wire_6173, wire_6172, wire_6153, wire_6152, wire_6133, wire_6132, wire_10909, wire_10908, wire_10889, wire_10888, wire_10869, wire_10868, wire_10849, wire_10848, wire_10829, wire_10828, wire_10809, wire_10808, wire_6619, wire_6618, wire_6599, wire_6598, wire_6579, wire_6578, wire_6559, wire_6558, wire_6539, wire_6538, wire_6519, wire_6518, wire_10519, wire_10518, wire_10499, wire_10498, wire_10479, wire_10478, wire_10459, wire_10458, wire_10439, wire_10438, wire_10419, wire_10418, wire_6229, wire_6228, wire_6209, wire_6208, wire_6189, wire_6188, wire_6169, wire_6168, wire_6149, wire_6148, wire_6129, wire_6128, wire_10905, wire_10904, wire_10885, wire_10884, wire_10865, wire_10864, wire_10845, wire_10844, wire_10825, wire_10824, wire_10805, wire_10804, wire_6615, wire_6614, wire_6595, wire_6594, wire_6575, wire_6574, wire_6555, wire_6554, wire_6535, wire_6534, wire_6515, wire_6514, wire_10517, wire_10516, wire_10497, wire_10496, wire_10477, wire_10476, wire_10457, wire_10456, wire_10437, wire_10436, wire_10417, wire_10416, wire_6225, wire_6224, wire_6205, wire_6204, wire_6185, wire_6184, wire_6165, wire_6164, wire_6145, wire_6144, wire_6125, wire_6124, wire_10911, wire_10910, wire_10883, wire_10882, wire_10871, wire_10870, wire_10843, wire_10842, wire_10831, wire_10830, wire_10803, wire_10802, wire_6611, wire_6610, wire_6591, wire_6590, wire_6571, wire_6570, wire_6551, wire_6550, wire_6531, wire_6530, wire_6511, wire_6510, wire_10513, wire_10512, wire_10493, wire_10492, wire_10473, wire_10472, wire_10453, wire_10452, wire_10433, wire_10432, wire_10413, wire_10412, wire_6221, wire_6220, wire_6201, wire_6200, wire_6181, wire_6180, wire_6161, wire_6160, wire_6141, wire_6140, wire_6121, wire_6120, wire_10899, wire_10898, wire_10887, wire_10886, wire_10859, wire_10858, wire_10847, wire_10846, wire_10819, wire_10818, wire_10807, wire_10806, wire_6609, wire_6608, wire_6597, wire_6596, wire_6569, wire_6568, wire_6557, wire_6556, wire_6529, wire_6528, wire_6517, wire_6516};
    // IPIN TOTAL: 276
    assign lut_tile_2_1_ipin_in = {wire_6627, wire_6626, wire_6607, wire_6606, wire_6587, wire_6586, wire_6567, wire_6566, wire_6547, wire_6546, wire_6527, wire_6526, wire_10915, wire_10914, wire_10903, wire_10902, wire_10875, wire_10874, wire_10863, wire_10862, wire_10835, wire_10834, wire_10823, wire_10822, wire_7013, wire_7012, wire_7001, wire_7000, wire_6973, wire_6972, wire_6961, wire_6960, wire_6933, wire_6932, wire_6921, wire_6920, wire_10559, wire_10558, wire_10549, wire_10548, wire_10539, wire_10538, wire_10513, wire_10512, wire_10473, wire_10472, wire_10433, wire_10432, wire_6623, wire_6622, wire_6603, wire_6602, wire_6583, wire_6582, wire_6563, wire_6562, wire_6543, wire_6542, wire_6523, wire_6522, wire_10919, wire_10918, wire_10891, wire_10890, wire_10879, wire_10878, wire_10851, wire_10850, wire_10839, wire_10838, wire_10811, wire_10810, wire_7017, wire_7016, wire_6989, wire_6988, wire_6977, wire_6976, wire_6949, wire_6948, wire_6937, wire_6936, wire_6909, wire_6908, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_10529, wire_10528, wire_10489, wire_10488, wire_10449, wire_10448, wire_6629, wire_6628, wire_6601, wire_6600, wire_6589, wire_6588, wire_6561, wire_6560, wire_6549, wire_6548, wire_6521, wire_6520, wire_10907, wire_10906, wire_10895, wire_10894, wire_10867, wire_10866, wire_10855, wire_10854, wire_10827, wire_10826, wire_10815, wire_10814, wire_7007, wire_7006, wire_6995, wire_6994, wire_6967, wire_6966, wire_6955, wire_6954, wire_6927, wire_6926, wire_6915, wire_6914, wire_10557, wire_10556, wire_10547, wire_10546, wire_10537, wire_10536, wire_10505, wire_10504, wire_10465, wire_10464, wire_10425, wire_10424, wire_6617, wire_6616, wire_6605, wire_6604, wire_6577, wire_6576, wire_6565, wire_6564, wire_6537, wire_6536, wire_6525, wire_6524, wire_10911, wire_10910, wire_10883, wire_10882, wire_10871, wire_10870, wire_10843, wire_10842, wire_10831, wire_10830, wire_10803, wire_10802, wire_7011, wire_7010, wire_6983, wire_6982, wire_6971, wire_6970, wire_6943, wire_6942, wire_6931, wire_6930, wire_6903, wire_6902, wire_10515, wire_10514, wire_10495, wire_10494, wire_10475, wire_10474, wire_10455, wire_10454, wire_10435, wire_10434, wire_10415, wire_10414, wire_6621, wire_6620, wire_6593, wire_6592, wire_6581, wire_6580, wire_6553, wire_6552, wire_6541, wire_6540, wire_6513, wire_6512, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_6999, wire_6998, wire_6987, wire_6986, wire_6959, wire_6958, wire_6947, wire_6946, wire_6919, wire_6918, wire_6907, wire_6906, wire_10511, wire_10510, wire_10491, wire_10490, wire_10471, wire_10470, wire_10451, wire_10450, wire_10431, wire_10430, wire_10411, wire_10410, wire_6609, wire_6608, wire_6597, wire_6596, wire_6569, wire_6568, wire_6557, wire_6556, wire_6529, wire_6528, wire_6517, wire_6516, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10897, wire_10896, wire_10857, wire_10856, wire_10817, wire_10816, wire_6997, wire_6996, wire_6985, wire_6984, wire_6957, wire_6956, wire_6945, wire_6944, wire_6917, wire_6916, wire_6905, wire_6904};
    // IPIN TOTAL: 276
    assign lut_tile_3_1_ipin_in = {wire_7015, wire_7014, wire_7003, wire_7002, wire_6975, wire_6974, wire_6963, wire_6962, wire_6935, wire_6934, wire_6923, wire_6922, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10913, wire_10912, wire_10873, wire_10872, wire_10833, wire_10832, wire_7409, wire_7408, wire_7389, wire_7388, wire_7369, wire_7368, wire_7349, wire_7348, wire_7329, wire_7328, wire_7309, wire_7308, wire_10585, wire_10584, wire_10575, wire_10574, wire_10565, wire_10564, wire_10523, wire_10522, wire_10483, wire_10482, wire_10443, wire_10442, wire_7019, wire_7018, wire_6991, wire_6990, wire_6979, wire_6978, wire_6951, wire_6950, wire_6939, wire_6938, wire_6911, wire_6910, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10889, wire_10888, wire_10849, wire_10848, wire_10809, wire_10808, wire_7405, wire_7404, wire_7385, wire_7384, wire_7365, wire_7364, wire_7345, wire_7344, wire_7325, wire_7324, wire_7305, wire_7304, wire_10589, wire_10588, wire_10579, wire_10578, wire_10569, wire_10568, wire_10499, wire_10498, wire_10459, wire_10458, wire_10419, wire_10418, wire_7017, wire_7016, wire_6989, wire_6988, wire_6977, wire_6976, wire_6949, wire_6948, wire_6937, wire_6936, wire_6909, wire_6908, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10905, wire_10904, wire_10865, wire_10864, wire_10825, wire_10824, wire_7395, wire_7394, wire_7383, wire_7382, wire_7355, wire_7354, wire_7343, wire_7342, wire_7315, wire_7314, wire_7303, wire_7302, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_10515, wire_10514, wire_10475, wire_10474, wire_10435, wire_10434, wire_7005, wire_7004, wire_6993, wire_6992, wire_6965, wire_6964, wire_6953, wire_6952, wire_6925, wire_6924, wire_6913, wire_6912, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_7399, wire_7398, wire_7371, wire_7370, wire_7359, wire_7358, wire_7331, wire_7330, wire_7319, wire_7318, wire_7291, wire_7290, wire_10551, wire_10550, wire_10541, wire_10540, wire_10531, wire_10530, wire_10521, wire_10520, wire_10481, wire_10480, wire_10441, wire_10440, wire_7009, wire_7008, wire_6981, wire_6980, wire_6969, wire_6968, wire_6941, wire_6940, wire_6929, wire_6928, wire_6901, wire_6900, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10907, wire_10906, wire_10867, wire_10866, wire_10827, wire_10826, wire_7387, wire_7386, wire_7375, wire_7374, wire_7347, wire_7346, wire_7335, wire_7334, wire_7307, wire_7306, wire_7295, wire_7294, wire_10555, wire_10554, wire_10545, wire_10544, wire_10535, wire_10534, wire_10497, wire_10496, wire_10457, wire_10456, wire_10417, wire_10416, wire_6997, wire_6996, wire_6985, wire_6984, wire_6957, wire_6956, wire_6945, wire_6944, wire_6917, wire_6916, wire_6905, wire_6904, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_7393, wire_7392, wire_7373, wire_7372, wire_7353, wire_7352, wire_7333, wire_7332, wire_7313, wire_7312, wire_7293, wire_7292};
    // IPIN TOTAL: 276
    assign lut_tile_4_1_ipin_in = {wire_7403, wire_7402, wire_7391, wire_7390, wire_7363, wire_7362, wire_7351, wire_7350, wire_7323, wire_7322, wire_7311, wire_7310, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10899, wire_10898, wire_10859, wire_10858, wire_10819, wire_10818, wire_7797, wire_7796, wire_7777, wire_7776, wire_7757, wire_7756, wire_7737, wire_7736, wire_7717, wire_7716, wire_7697, wire_7696, wire_10619, wire_10618, wire_10609, wire_10608, wire_10599, wire_10598, wire_10555, wire_10554, wire_10545, wire_10544, wire_10535, wire_10534, wire_7407, wire_7406, wire_7379, wire_7378, wire_7367, wire_7366, wire_7339, wire_7338, wire_7327, wire_7326, wire_7299, wire_7298, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10915, wire_10914, wire_10875, wire_10874, wire_10835, wire_10834, wire_7793, wire_7792, wire_7773, wire_7772, wire_7753, wire_7752, wire_7733, wire_7732, wire_7713, wire_7712, wire_7693, wire_7692, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_10559, wire_10558, wire_10549, wire_10548, wire_10539, wire_10538, wire_7405, wire_7404, wire_7385, wire_7384, wire_7365, wire_7364, wire_7345, wire_7344, wire_7325, wire_7324, wire_7305, wire_7304, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10891, wire_10890, wire_10851, wire_10850, wire_10811, wire_10810, wire_7791, wire_7790, wire_7771, wire_7770, wire_7751, wire_7750, wire_7731, wire_7730, wire_7711, wire_7710, wire_7691, wire_7690, wire_10617, wire_10616, wire_10607, wire_10606, wire_10597, wire_10596, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_7401, wire_7400, wire_7381, wire_7380, wire_7361, wire_7360, wire_7341, wire_7340, wire_7321, wire_7320, wire_7301, wire_7300, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10907, wire_10906, wire_10867, wire_10866, wire_10827, wire_10826, wire_7787, wire_7786, wire_7767, wire_7766, wire_7747, wire_7746, wire_7727, wire_7726, wire_7707, wire_7706, wire_7687, wire_7686, wire_10587, wire_10586, wire_10577, wire_10576, wire_10567, wire_10566, wire_10491, wire_10490, wire_10451, wire_10450, wire_10411, wire_10410, wire_7397, wire_7396, wire_7377, wire_7376, wire_7357, wire_7356, wire_7337, wire_7336, wire_7317, wire_7316, wire_7297, wire_7296, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_7783, wire_7782, wire_7763, wire_7762, wire_7743, wire_7742, wire_7723, wire_7722, wire_7703, wire_7702, wire_7683, wire_7682, wire_10581, wire_10580, wire_10571, wire_10570, wire_10561, wire_10560, wire_10507, wire_10506, wire_10467, wire_10466, wire_10427, wire_10426, wire_7393, wire_7392, wire_7373, wire_7372, wire_7353, wire_7352, wire_7333, wire_7332, wire_7313, wire_7312, wire_7293, wire_7292, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_7781, wire_7780, wire_7761, wire_7760, wire_7741, wire_7740, wire_7721, wire_7720, wire_7701, wire_7700, wire_7681, wire_7680};
    // IPIN TOTAL: 276
    assign lut_tile_5_1_ipin_in = {wire_7799, wire_7798, wire_7779, wire_7778, wire_7759, wire_7758, wire_7739, wire_7738, wire_7719, wire_7718, wire_7699, wire_7698, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_8185, wire_8184, wire_8173, wire_8172, wire_8145, wire_8144, wire_8133, wire_8132, wire_8105, wire_8104, wire_8093, wire_8092, wire_10645, wire_10644, wire_10635, wire_10634, wire_10625, wire_10624, wire_10589, wire_10588, wire_10579, wire_10578, wire_10569, wire_10568, wire_7795, wire_7794, wire_7775, wire_7774, wire_7755, wire_7754, wire_7735, wire_7734, wire_7715, wire_7714, wire_7695, wire_7694, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_8189, wire_8188, wire_8161, wire_8160, wire_8149, wire_8148, wire_8121, wire_8120, wire_8109, wire_8108, wire_8081, wire_8080, wire_10649, wire_10648, wire_10639, wire_10638, wire_10629, wire_10628, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_7793, wire_7792, wire_7773, wire_7772, wire_7753, wire_7752, wire_7733, wire_7732, wire_7713, wire_7712, wire_7693, wire_7692, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_8179, wire_8178, wire_8159, wire_8158, wire_8139, wire_8138, wire_8119, wire_8118, wire_8099, wire_8098, wire_8079, wire_8078, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_10587, wire_10586, wire_10577, wire_10576, wire_10567, wire_10566, wire_7789, wire_7788, wire_7769, wire_7768, wire_7749, wire_7748, wire_7729, wire_7728, wire_7709, wire_7708, wire_7689, wire_7688, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_8175, wire_8174, wire_8155, wire_8154, wire_8135, wire_8134, wire_8115, wire_8114, wire_8095, wire_8094, wire_8075, wire_8074, wire_10611, wire_10610, wire_10601, wire_10600, wire_10591, wire_10590, wire_10557, wire_10556, wire_10547, wire_10546, wire_10537, wire_10536, wire_7785, wire_7784, wire_7765, wire_7764, wire_7745, wire_7744, wire_7725, wire_7724, wire_7705, wire_7704, wire_7685, wire_7684, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_8171, wire_8170, wire_8151, wire_8150, wire_8131, wire_8130, wire_8111, wire_8110, wire_8091, wire_8090, wire_8071, wire_8070, wire_10615, wire_10614, wire_10605, wire_10604, wire_10595, wire_10594, wire_10551, wire_10550, wire_10541, wire_10540, wire_10531, wire_10530, wire_7781, wire_7780, wire_7761, wire_7760, wire_7741, wire_7740, wire_7721, wire_7720, wire_7701, wire_7700, wire_7681, wire_7680, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_8169, wire_8168, wire_8157, wire_8156, wire_8129, wire_8128, wire_8117, wire_8116, wire_8089, wire_8088, wire_8077, wire_8076};
    // IPIN TOTAL: 276
    assign lut_tile_6_1_ipin_in = {wire_8187, wire_8186, wire_8167, wire_8166, wire_8147, wire_8146, wire_8127, wire_8126, wire_8107, wire_8106, wire_8087, wire_8086, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_8573, wire_8572, wire_8561, wire_8560, wire_8533, wire_8532, wire_8521, wire_8520, wire_8493, wire_8492, wire_8481, wire_8480, wire_10679, wire_10678, wire_10669, wire_10668, wire_10659, wire_10658, wire_10615, wire_10614, wire_10605, wire_10604, wire_10595, wire_10594, wire_8183, wire_8182, wire_8163, wire_8162, wire_8143, wire_8142, wire_8123, wire_8122, wire_8103, wire_8102, wire_8083, wire_8082, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_8577, wire_8576, wire_8549, wire_8548, wire_8537, wire_8536, wire_8509, wire_8508, wire_8497, wire_8496, wire_8469, wire_8468, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_10619, wire_10618, wire_10609, wire_10608, wire_10599, wire_10598, wire_8189, wire_8188, wire_8161, wire_8160, wire_8149, wire_8148, wire_8121, wire_8120, wire_8109, wire_8108, wire_8081, wire_8080, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_8567, wire_8566, wire_8555, wire_8554, wire_8527, wire_8526, wire_8515, wire_8514, wire_8487, wire_8486, wire_8475, wire_8474, wire_10677, wire_10676, wire_10667, wire_10666, wire_10657, wire_10656, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_8177, wire_8176, wire_8165, wire_8164, wire_8137, wire_8136, wire_8125, wire_8124, wire_8097, wire_8096, wire_8085, wire_8084, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_8571, wire_8570, wire_8543, wire_8542, wire_8531, wire_8530, wire_8503, wire_8502, wire_8491, wire_8490, wire_8463, wire_8462, wire_10647, wire_10646, wire_10637, wire_10636, wire_10627, wire_10626, wire_10581, wire_10580, wire_10571, wire_10570, wire_10561, wire_10560, wire_8181, wire_8180, wire_8153, wire_8152, wire_8141, wire_8140, wire_8113, wire_8112, wire_8101, wire_8100, wire_8073, wire_8072, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_8559, wire_8558, wire_8547, wire_8546, wire_8519, wire_8518, wire_8507, wire_8506, wire_8479, wire_8478, wire_8467, wire_8466, wire_10641, wire_10640, wire_10631, wire_10630, wire_10621, wire_10620, wire_10585, wire_10584, wire_10575, wire_10574, wire_10565, wire_10564, wire_8169, wire_8168, wire_8157, wire_8156, wire_8129, wire_8128, wire_8117, wire_8116, wire_8089, wire_8088, wire_8077, wire_8076, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_8557, wire_8556, wire_8545, wire_8544, wire_8517, wire_8516, wire_8505, wire_8504, wire_8477, wire_8476, wire_8465, wire_8464};
    // IPIN TOTAL: 276
    assign lut_tile_7_1_ipin_in = {wire_8575, wire_8574, wire_8563, wire_8562, wire_8535, wire_8534, wire_8523, wire_8522, wire_8495, wire_8494, wire_8483, wire_8482, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_8969, wire_8968, wire_8949, wire_8948, wire_8929, wire_8928, wire_8909, wire_8908, wire_8889, wire_8888, wire_8869, wire_8868, wire_10705, wire_10704, wire_10695, wire_10694, wire_10685, wire_10684, wire_10649, wire_10648, wire_10639, wire_10638, wire_10629, wire_10628, wire_8579, wire_8578, wire_8551, wire_8550, wire_8539, wire_8538, wire_8511, wire_8510, wire_8499, wire_8498, wire_8471, wire_8470, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_8965, wire_8964, wire_8945, wire_8944, wire_8925, wire_8924, wire_8905, wire_8904, wire_8885, wire_8884, wire_8865, wire_8864, wire_10709, wire_10708, wire_10699, wire_10698, wire_10689, wire_10688, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_8577, wire_8576, wire_8549, wire_8548, wire_8537, wire_8536, wire_8509, wire_8508, wire_8497, wire_8496, wire_8469, wire_8468, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_8955, wire_8954, wire_8943, wire_8942, wire_8915, wire_8914, wire_8903, wire_8902, wire_8875, wire_8874, wire_8863, wire_8862, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_10647, wire_10646, wire_10637, wire_10636, wire_10627, wire_10626, wire_8565, wire_8564, wire_8553, wire_8552, wire_8525, wire_8524, wire_8513, wire_8512, wire_8485, wire_8484, wire_8473, wire_8472, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_8959, wire_8958, wire_8931, wire_8930, wire_8919, wire_8918, wire_8891, wire_8890, wire_8879, wire_8878, wire_8851, wire_8850, wire_10671, wire_10670, wire_10661, wire_10660, wire_10651, wire_10650, wire_10617, wire_10616, wire_10607, wire_10606, wire_10597, wire_10596, wire_8569, wire_8568, wire_8541, wire_8540, wire_8529, wire_8528, wire_8501, wire_8500, wire_8489, wire_8488, wire_8461, wire_8460, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_8947, wire_8946, wire_8935, wire_8934, wire_8907, wire_8906, wire_8895, wire_8894, wire_8867, wire_8866, wire_8855, wire_8854, wire_10675, wire_10674, wire_10665, wire_10664, wire_10655, wire_10654, wire_10611, wire_10610, wire_10601, wire_10600, wire_10591, wire_10590, wire_8557, wire_8556, wire_8545, wire_8544, wire_8517, wire_8516, wire_8505, wire_8504, wire_8477, wire_8476, wire_8465, wire_8464, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_8953, wire_8952, wire_8933, wire_8932, wire_8913, wire_8912, wire_8893, wire_8892, wire_8873, wire_8872, wire_8853, wire_8852};
    // IPIN TOTAL: 276
    assign lut_tile_8_1_ipin_in = {wire_8963, wire_8962, wire_8951, wire_8950, wire_8923, wire_8922, wire_8911, wire_8910, wire_8883, wire_8882, wire_8871, wire_8870, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_9357, wire_9356, wire_9337, wire_9336, wire_9317, wire_9316, wire_9297, wire_9296, wire_9277, wire_9276, wire_9257, wire_9256, wire_10739, wire_10738, wire_10729, wire_10728, wire_10719, wire_10718, wire_10675, wire_10674, wire_10665, wire_10664, wire_10655, wire_10654, wire_8967, wire_8966, wire_8939, wire_8938, wire_8927, wire_8926, wire_8899, wire_8898, wire_8887, wire_8886, wire_8859, wire_8858, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_9353, wire_9352, wire_9333, wire_9332, wire_9313, wire_9312, wire_9293, wire_9292, wire_9273, wire_9272, wire_9253, wire_9252, wire_10733, wire_10732, wire_10723, wire_10722, wire_10713, wire_10712, wire_10679, wire_10678, wire_10669, wire_10668, wire_10659, wire_10658, wire_8965, wire_8964, wire_8945, wire_8944, wire_8925, wire_8924, wire_8905, wire_8904, wire_8885, wire_8884, wire_8865, wire_8864, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_9351, wire_9350, wire_9331, wire_9330, wire_9311, wire_9310, wire_9291, wire_9290, wire_9271, wire_9270, wire_9251, wire_9250, wire_10737, wire_10736, wire_10727, wire_10726, wire_10717, wire_10716, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_8961, wire_8960, wire_8941, wire_8940, wire_8921, wire_8920, wire_8901, wire_8900, wire_8881, wire_8880, wire_8861, wire_8860, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_9347, wire_9346, wire_9327, wire_9326, wire_9307, wire_9306, wire_9287, wire_9286, wire_9267, wire_9266, wire_9247, wire_9246, wire_10707, wire_10706, wire_10697, wire_10696, wire_10687, wire_10686, wire_10641, wire_10640, wire_10631, wire_10630, wire_10621, wire_10620, wire_8957, wire_8956, wire_8937, wire_8936, wire_8917, wire_8916, wire_8897, wire_8896, wire_8877, wire_8876, wire_8857, wire_8856, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_9343, wire_9342, wire_9323, wire_9322, wire_9303, wire_9302, wire_9283, wire_9282, wire_9263, wire_9262, wire_9243, wire_9242, wire_10701, wire_10700, wire_10691, wire_10690, wire_10681, wire_10680, wire_10645, wire_10644, wire_10635, wire_10634, wire_10625, wire_10624, wire_8953, wire_8952, wire_8933, wire_8932, wire_8913, wire_8912, wire_8893, wire_8892, wire_8873, wire_8872, wire_8853, wire_8852, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_9341, wire_9340, wire_9321, wire_9320, wire_9301, wire_9300, wire_9281, wire_9280, wire_9261, wire_9260, wire_9241, wire_9240};
    // IPIN TOTAL: 276
    assign lut_tile_9_1_ipin_in = {wire_9359, wire_9358, wire_9339, wire_9338, wire_9319, wire_9318, wire_9299, wire_9298, wire_9279, wire_9278, wire_9259, wire_9258, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_9745, wire_9744, wire_9733, wire_9732, wire_9705, wire_9704, wire_9693, wire_9692, wire_9665, wire_9664, wire_9653, wire_9652, wire_10765, wire_10764, wire_10755, wire_10754, wire_10745, wire_10744, wire_10709, wire_10708, wire_10699, wire_10698, wire_10689, wire_10688, wire_9355, wire_9354, wire_9335, wire_9334, wire_9315, wire_9314, wire_9295, wire_9294, wire_9275, wire_9274, wire_9255, wire_9254, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_9749, wire_9748, wire_9721, wire_9720, wire_9709, wire_9708, wire_9681, wire_9680, wire_9669, wire_9668, wire_9641, wire_9640, wire_10769, wire_10768, wire_10759, wire_10758, wire_10749, wire_10748, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_9353, wire_9352, wire_9333, wire_9332, wire_9313, wire_9312, wire_9293, wire_9292, wire_9273, wire_9272, wire_9253, wire_9252, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_9739, wire_9738, wire_9719, wire_9718, wire_9699, wire_9698, wire_9679, wire_9678, wire_9659, wire_9658, wire_9639, wire_9638, wire_10763, wire_10762, wire_10753, wire_10752, wire_10743, wire_10742, wire_10707, wire_10706, wire_10697, wire_10696, wire_10687, wire_10686, wire_9349, wire_9348, wire_9329, wire_9328, wire_9309, wire_9308, wire_9289, wire_9288, wire_9269, wire_9268, wire_9249, wire_9248, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_9735, wire_9734, wire_9715, wire_9714, wire_9695, wire_9694, wire_9675, wire_9674, wire_9655, wire_9654, wire_9635, wire_9634, wire_10731, wire_10730, wire_10721, wire_10720, wire_10711, wire_10710, wire_10677, wire_10676, wire_10667, wire_10666, wire_10657, wire_10656, wire_9345, wire_9344, wire_9325, wire_9324, wire_9305, wire_9304, wire_9285, wire_9284, wire_9265, wire_9264, wire_9245, wire_9244, wire_11151, wire_11150, wire_11141, wire_11140, wire_11131, wire_11130, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_9731, wire_9730, wire_9711, wire_9710, wire_9691, wire_9690, wire_9671, wire_9670, wire_9651, wire_9650, wire_9631, wire_9630, wire_10735, wire_10734, wire_10725, wire_10724, wire_10715, wire_10714, wire_10671, wire_10670, wire_10661, wire_10660, wire_10651, wire_10650, wire_9341, wire_9340, wire_9321, wire_9320, wire_9301, wire_9300, wire_9281, wire_9280, wire_9261, wire_9260, wire_9241, wire_9240, wire_11155, wire_11154, wire_11145, wire_11144, wire_11135, wire_11134, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_9729, wire_9728, wire_9717, wire_9716, wire_9689, wire_9688, wire_9677, wire_9676, wire_9649, wire_9648, wire_9637, wire_9636};
    // IPIN TOTAL: 276
    assign lut_tile_10_1_ipin_in = {wire_9747, wire_9746, wire_9727, wire_9726, wire_9707, wire_9706, wire_9687, wire_9686, wire_9667, wire_9666, wire_9647, wire_9646, wire_11159, wire_11158, wire_11149, wire_11148, wire_11139, wire_11138, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_10133, wire_10132, wire_10121, wire_10120, wire_10093, wire_10092, wire_10081, wire_10080, wire_10053, wire_10052, wire_10041, wire_10040, wire_10799, wire_10798, wire_10789, wire_10788, wire_10779, wire_10778, wire_10735, wire_10734, wire_10725, wire_10724, wire_10715, wire_10714, wire_9743, wire_9742, wire_9723, wire_9722, wire_9703, wire_9702, wire_9683, wire_9682, wire_9663, wire_9662, wire_9643, wire_9642, wire_11153, wire_11152, wire_11143, wire_11142, wire_11133, wire_11132, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_10137, wire_10136, wire_10109, wire_10108, wire_10097, wire_10096, wire_10069, wire_10068, wire_10057, wire_10056, wire_10029, wire_10028, wire_10793, wire_10792, wire_10783, wire_10782, wire_10773, wire_10772, wire_10739, wire_10738, wire_10729, wire_10728, wire_10719, wire_10718, wire_9749, wire_9748, wire_9721, wire_9720, wire_9709, wire_9708, wire_9681, wire_9680, wire_9669, wire_9668, wire_9641, wire_9640, wire_11157, wire_11156, wire_11147, wire_11146, wire_11137, wire_11136, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_10127, wire_10126, wire_10115, wire_10114, wire_10087, wire_10086, wire_10075, wire_10074, wire_10047, wire_10046, wire_10035, wire_10034, wire_10797, wire_10796, wire_10787, wire_10786, wire_10777, wire_10776, wire_10733, wire_10732, wire_10723, wire_10722, wire_10713, wire_10712, wire_9737, wire_9736, wire_9725, wire_9724, wire_9697, wire_9696, wire_9685, wire_9684, wire_9657, wire_9656, wire_9645, wire_9644, wire_11151, wire_11150, wire_11141, wire_11140, wire_11131, wire_11130, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_10131, wire_10130, wire_10103, wire_10102, wire_10091, wire_10090, wire_10063, wire_10062, wire_10051, wire_10050, wire_10023, wire_10022, wire_10767, wire_10766, wire_10757, wire_10756, wire_10747, wire_10746, wire_10701, wire_10700, wire_10691, wire_10690, wire_10681, wire_10680, wire_9741, wire_9740, wire_9713, wire_9712, wire_9701, wire_9700, wire_9673, wire_9672, wire_9661, wire_9660, wire_9633, wire_9632, wire_11187, wire_11186, wire_11177, wire_11176, wire_11167, wire_11166, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_10119, wire_10118, wire_10107, wire_10106, wire_10079, wire_10078, wire_10067, wire_10066, wire_10039, wire_10038, wire_10027, wire_10026, wire_10761, wire_10760, wire_10751, wire_10750, wire_10741, wire_10740, wire_10705, wire_10704, wire_10695, wire_10694, wire_10685, wire_10684, wire_9729, wire_9728, wire_9717, wire_9716, wire_9689, wire_9688, wire_9677, wire_9676, wire_9649, wire_9648, wire_9637, wire_9636, wire_11181, wire_11180, wire_11171, wire_11170, wire_11161, wire_11160, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_10117, wire_10116, wire_10105, wire_10104, wire_10077, wire_10076, wire_10065, wire_10064, wire_10037, wire_10036, wire_10025, wire_10024};
    // IPIN TOTAL: 276
    assign lut_tile_1_2_ipin_in = {wire_6237, wire_6236, wire_6217, wire_6216, wire_6197, wire_6196, wire_6177, wire_6176, wire_6157, wire_6156, wire_6137, wire_6136, wire_11305, wire_11304, wire_11293, wire_11292, wire_11265, wire_11264, wire_11253, wire_11252, wire_11225, wire_11224, wire_11213, wire_11212, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6623, wire_6622, wire_6583, wire_6582, wire_6543, wire_6542, wire_10915, wire_10914, wire_10903, wire_10902, wire_10875, wire_10874, wire_10863, wire_10862, wire_10835, wire_10834, wire_10823, wire_10822, wire_6233, wire_6232, wire_6213, wire_6212, wire_6193, wire_6192, wire_6173, wire_6172, wire_6153, wire_6152, wire_6133, wire_6132, wire_11309, wire_11308, wire_11281, wire_11280, wire_11269, wire_11268, wire_11241, wire_11240, wire_11229, wire_11228, wire_11201, wire_11200, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6599, wire_6598, wire_6559, wire_6558, wire_6519, wire_6518, wire_10919, wire_10918, wire_10891, wire_10890, wire_10879, wire_10878, wire_10851, wire_10850, wire_10839, wire_10838, wire_10811, wire_10810, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_6239, wire_6238, wire_6199, wire_6198, wire_6159, wire_6158, wire_11297, wire_11296, wire_11285, wire_11284, wire_11257, wire_11256, wire_11245, wire_11244, wire_11217, wire_11216, wire_11205, wire_11204, wire_6617, wire_6616, wire_6605, wire_6604, wire_6577, wire_6576, wire_6565, wire_6564, wire_6537, wire_6536, wire_6525, wire_6524, wire_10907, wire_10906, wire_10895, wire_10894, wire_10867, wire_10866, wire_10855, wire_10854, wire_10827, wire_10826, wire_10815, wire_10814, wire_6267, wire_6266, wire_6257, wire_6256, wire_6247, wire_6246, wire_6215, wire_6214, wire_6175, wire_6174, wire_6135, wire_6134, wire_11301, wire_11300, wire_11273, wire_11272, wire_11261, wire_11260, wire_11233, wire_11232, wire_11221, wire_11220, wire_11193, wire_11192, wire_6621, wire_6620, wire_6593, wire_6592, wire_6581, wire_6580, wire_6553, wire_6552, wire_6541, wire_6540, wire_6513, wire_6512, wire_10905, wire_10904, wire_10885, wire_10884, wire_10865, wire_10864, wire_10845, wire_10844, wire_10825, wire_10824, wire_10805, wire_10804, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240, wire_6231, wire_6230, wire_6191, wire_6190, wire_6151, wire_6150, wire_11299, wire_11298, wire_11271, wire_11270, wire_11259, wire_11258, wire_11231, wire_11230, wire_11219, wire_11218, wire_11191, wire_11190, wire_6609, wire_6608, wire_6597, wire_6596, wire_6569, wire_6568, wire_6557, wire_6556, wire_6529, wire_6528, wire_6517, wire_6516, wire_10901, wire_10900, wire_10881, wire_10880, wire_10861, wire_10860, wire_10841, wire_10840, wire_10821, wire_10820, wire_10801, wire_10800, wire_6265, wire_6264, wire_6255, wire_6254, wire_6245, wire_6244, wire_6207, wire_6206, wire_6167, wire_6166, wire_6127, wire_6126, wire_11287, wire_11286, wire_11275, wire_11274, wire_11247, wire_11246, wire_11235, wire_11234, wire_11207, wire_11206, wire_11195, wire_11194, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6607, wire_6606, wire_6567, wire_6566, wire_6527, wire_6526};
    // IPIN TOTAL: 276
    assign lut_tile_2_2_ipin_in = {wire_6625, wire_6624, wire_6613, wire_6612, wire_6585, wire_6584, wire_6573, wire_6572, wire_6545, wire_6544, wire_6533, wire_6532, wire_11303, wire_11302, wire_11291, wire_11290, wire_11263, wire_11262, wire_11251, wire_11250, wire_11223, wire_11222, wire_11211, wire_11210, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6999, wire_6998, wire_6959, wire_6958, wire_6919, wire_6918, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10913, wire_10912, wire_10873, wire_10872, wire_10833, wire_10832, wire_6629, wire_6628, wire_6601, wire_6600, wire_6589, wire_6588, wire_6561, wire_6560, wire_6549, wire_6548, wire_6521, wire_6520, wire_11307, wire_11306, wire_11279, wire_11278, wire_11267, wire_11266, wire_11239, wire_11238, wire_11227, wire_11226, wire_11199, wire_11198, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10889, wire_10888, wire_10849, wire_10848, wire_10809, wire_10808, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6599, wire_6598, wire_6559, wire_6558, wire_6519, wire_6518, wire_11295, wire_11294, wire_11283, wire_11282, wire_11255, wire_11254, wire_11243, wire_11242, wire_11215, wire_11214, wire_11203, wire_11202, wire_7005, wire_7004, wire_6993, wire_6992, wire_6965, wire_6964, wire_6953, wire_6952, wire_6925, wire_6924, wire_6913, wire_6912, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10905, wire_10904, wire_10865, wire_10864, wire_10825, wire_10824, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6615, wire_6614, wire_6575, wire_6574, wire_6535, wire_6534, wire_11299, wire_11298, wire_11271, wire_11270, wire_11259, wire_11258, wire_11231, wire_11230, wire_11219, wire_11218, wire_11191, wire_11190, wire_7009, wire_7008, wire_6981, wire_6980, wire_6969, wire_6968, wire_6941, wire_6940, wire_6929, wire_6928, wire_6901, wire_6900, wire_10911, wire_10910, wire_10883, wire_10882, wire_10871, wire_10870, wire_10843, wire_10842, wire_10831, wire_10830, wire_10803, wire_10802, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6591, wire_6590, wire_6551, wire_6550, wire_6511, wire_6510, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11297, wire_11296, wire_11257, wire_11256, wire_11217, wire_11216, wire_6997, wire_6996, wire_6985, wire_6984, wire_6957, wire_6956, wire_6945, wire_6944, wire_6917, wire_6916, wire_6905, wire_6904, wire_10899, wire_10898, wire_10887, wire_10886, wire_10859, wire_10858, wire_10847, wire_10846, wire_10819, wire_10818, wire_10807, wire_10806, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6607, wire_6606, wire_6567, wire_6566, wire_6527, wire_6526, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11273, wire_11272, wire_11233, wire_11232, wire_11193, wire_11192, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6983, wire_6982, wire_6943, wire_6942, wire_6903, wire_6902};
    // IPIN TOTAL: 276
    assign lut_tile_3_2_ipin_in = {wire_7013, wire_7012, wire_7001, wire_7000, wire_6973, wire_6972, wire_6961, wire_6960, wire_6933, wire_6932, wire_6921, wire_6920, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11289, wire_11288, wire_11249, wire_11248, wire_11209, wire_11208, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7407, wire_7406, wire_7367, wire_7366, wire_7327, wire_7326, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10899, wire_10898, wire_10859, wire_10858, wire_10819, wire_10818, wire_7017, wire_7016, wire_6989, wire_6988, wire_6977, wire_6976, wire_6949, wire_6948, wire_6937, wire_6936, wire_6909, wire_6908, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11305, wire_11304, wire_11265, wire_11264, wire_11225, wire_11224, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7383, wire_7382, wire_7343, wire_7342, wire_7303, wire_7302, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10915, wire_10914, wire_10875, wire_10874, wire_10835, wire_10834, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11281, wire_11280, wire_11241, wire_11240, wire_11201, wire_11200, wire_7401, wire_7400, wire_7381, wire_7380, wire_7361, wire_7360, wire_7341, wire_7340, wire_7321, wire_7320, wire_7301, wire_7300, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10891, wire_10890, wire_10851, wire_10850, wire_10811, wire_10810, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6991, wire_6990, wire_6951, wire_6950, wire_6911, wire_6910, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11297, wire_11296, wire_11257, wire_11256, wire_11217, wire_11216, wire_7397, wire_7396, wire_7377, wire_7376, wire_7357, wire_7356, wire_7337, wire_7336, wire_7317, wire_7316, wire_7297, wire_7296, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_7007, wire_7006, wire_6967, wire_6966, wire_6927, wire_6926, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_7393, wire_7392, wire_7373, wire_7372, wire_7353, wire_7352, wire_7333, wire_7332, wire_7313, wire_7312, wire_7293, wire_7292, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10897, wire_10896, wire_10857, wire_10856, wire_10817, wire_10816, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6983, wire_6982, wire_6943, wire_6942, wire_6903, wire_6902, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11291, wire_11290, wire_11251, wire_11250, wire_11211, wire_11210, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7391, wire_7390, wire_7351, wire_7350, wire_7311, wire_7310};
    // IPIN TOTAL: 276
    assign lut_tile_4_2_ipin_in = {wire_7409, wire_7408, wire_7389, wire_7388, wire_7369, wire_7368, wire_7349, wire_7348, wire_7329, wire_7328, wire_7309, wire_7308, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11307, wire_11306, wire_11267, wire_11266, wire_11227, wire_11226, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7783, wire_7782, wire_7743, wire_7742, wire_7703, wire_7702, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_7405, wire_7404, wire_7385, wire_7384, wire_7365, wire_7364, wire_7345, wire_7344, wire_7325, wire_7324, wire_7305, wire_7304, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11283, wire_11282, wire_11243, wire_11242, wire_11203, wire_11202, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7383, wire_7382, wire_7343, wire_7342, wire_7303, wire_7302, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11299, wire_11298, wire_11259, wire_11258, wire_11219, wire_11218, wire_7789, wire_7788, wire_7769, wire_7768, wire_7749, wire_7748, wire_7729, wire_7728, wire_7709, wire_7708, wire_7689, wire_7688, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7399, wire_7398, wire_7359, wire_7358, wire_7319, wire_7318, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_7785, wire_7784, wire_7765, wire_7764, wire_7745, wire_7744, wire_7725, wire_7724, wire_7705, wire_7704, wire_7685, wire_7684, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10907, wire_10906, wire_10867, wire_10866, wire_10827, wire_10826, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7375, wire_7374, wire_7335, wire_7334, wire_7295, wire_7294, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_7781, wire_7780, wire_7761, wire_7760, wire_7741, wire_7740, wire_7721, wire_7720, wire_7701, wire_7700, wire_7681, wire_7680, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7391, wire_7390, wire_7351, wire_7350, wire_7311, wire_7310, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7767, wire_7766, wire_7727, wire_7726, wire_7687, wire_7686};
    // IPIN TOTAL: 276
    assign lut_tile_5_2_ipin_in = {wire_7797, wire_7796, wire_7777, wire_7776, wire_7757, wire_7756, wire_7737, wire_7736, wire_7717, wire_7716, wire_7697, wire_7696, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8183, wire_8182, wire_8143, wire_8142, wire_8103, wire_8102, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_7793, wire_7792, wire_7773, wire_7772, wire_7753, wire_7752, wire_7733, wire_7732, wire_7713, wire_7712, wire_7693, wire_7692, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8159, wire_8158, wire_8119, wire_8118, wire_8079, wire_8078, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_8177, wire_8176, wire_8165, wire_8164, wire_8137, wire_8136, wire_8125, wire_8124, wire_8097, wire_8096, wire_8085, wire_8084, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7775, wire_7774, wire_7735, wire_7734, wire_7695, wire_7694, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_8181, wire_8180, wire_8153, wire_8152, wire_8141, wire_8140, wire_8113, wire_8112, wire_8101, wire_8100, wire_8073, wire_8072, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7791, wire_7790, wire_7751, wire_7750, wire_7711, wire_7710, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_8169, wire_8168, wire_8157, wire_8156, wire_8129, wire_8128, wire_8117, wire_8116, wire_8089, wire_8088, wire_8077, wire_8076, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7767, wire_7766, wire_7727, wire_7726, wire_7687, wire_7686, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8167, wire_8166, wire_8127, wire_8126, wire_8087, wire_8086};
    // IPIN TOTAL: 276
    assign lut_tile_6_2_ipin_in = {wire_8185, wire_8184, wire_8173, wire_8172, wire_8145, wire_8144, wire_8133, wire_8132, wire_8105, wire_8104, wire_8093, wire_8092, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8559, wire_8558, wire_8519, wire_8518, wire_8479, wire_8478, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_8189, wire_8188, wire_8161, wire_8160, wire_8149, wire_8148, wire_8121, wire_8120, wire_8109, wire_8108, wire_8081, wire_8080, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8159, wire_8158, wire_8119, wire_8118, wire_8079, wire_8078, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_8565, wire_8564, wire_8553, wire_8552, wire_8525, wire_8524, wire_8513, wire_8512, wire_8485, wire_8484, wire_8473, wire_8472, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8175, wire_8174, wire_8135, wire_8134, wire_8095, wire_8094, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_8569, wire_8568, wire_8541, wire_8540, wire_8529, wire_8528, wire_8501, wire_8500, wire_8489, wire_8488, wire_8461, wire_8460, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8151, wire_8150, wire_8111, wire_8110, wire_8071, wire_8070, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_8557, wire_8556, wire_8545, wire_8544, wire_8517, wire_8516, wire_8505, wire_8504, wire_8477, wire_8476, wire_8465, wire_8464, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8167, wire_8166, wire_8127, wire_8126, wire_8087, wire_8086, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8543, wire_8542, wire_8503, wire_8502, wire_8463, wire_8462};
    // IPIN TOTAL: 276
    assign lut_tile_7_2_ipin_in = {wire_8573, wire_8572, wire_8561, wire_8560, wire_8533, wire_8532, wire_8521, wire_8520, wire_8493, wire_8492, wire_8481, wire_8480, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8967, wire_8966, wire_8927, wire_8926, wire_8887, wire_8886, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_8577, wire_8576, wire_8549, wire_8548, wire_8537, wire_8536, wire_8509, wire_8508, wire_8497, wire_8496, wire_8469, wire_8468, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8943, wire_8942, wire_8903, wire_8902, wire_8863, wire_8862, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_8961, wire_8960, wire_8941, wire_8940, wire_8921, wire_8920, wire_8901, wire_8900, wire_8881, wire_8880, wire_8861, wire_8860, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8551, wire_8550, wire_8511, wire_8510, wire_8471, wire_8470, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_8957, wire_8956, wire_8937, wire_8936, wire_8917, wire_8916, wire_8897, wire_8896, wire_8877, wire_8876, wire_8857, wire_8856, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8567, wire_8566, wire_8527, wire_8526, wire_8487, wire_8486, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_8953, wire_8952, wire_8933, wire_8932, wire_8913, wire_8912, wire_8893, wire_8892, wire_8873, wire_8872, wire_8853, wire_8852, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8543, wire_8542, wire_8503, wire_8502, wire_8463, wire_8462, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8951, wire_8950, wire_8911, wire_8910, wire_8871, wire_8870};
    // IPIN TOTAL: 276
    assign lut_tile_8_2_ipin_in = {wire_8969, wire_8968, wire_8949, wire_8948, wire_8929, wire_8928, wire_8909, wire_8908, wire_8889, wire_8888, wire_8869, wire_8868, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9343, wire_9342, wire_9303, wire_9302, wire_9263, wire_9262, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_8965, wire_8964, wire_8945, wire_8944, wire_8925, wire_8924, wire_8905, wire_8904, wire_8885, wire_8884, wire_8865, wire_8864, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8943, wire_8942, wire_8903, wire_8902, wire_8863, wire_8862, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_9349, wire_9348, wire_9329, wire_9328, wire_9309, wire_9308, wire_9289, wire_9288, wire_9269, wire_9268, wire_9249, wire_9248, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8959, wire_8958, wire_8919, wire_8918, wire_8879, wire_8878, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_9345, wire_9344, wire_9325, wire_9324, wire_9305, wire_9304, wire_9285, wire_9284, wire_9265, wire_9264, wire_9245, wire_9244, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8935, wire_8934, wire_8895, wire_8894, wire_8855, wire_8854, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_9341, wire_9340, wire_9321, wire_9320, wire_9301, wire_9300, wire_9281, wire_9280, wire_9261, wire_9260, wire_9241, wire_9240, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8951, wire_8950, wire_8911, wire_8910, wire_8871, wire_8870, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9327, wire_9326, wire_9287, wire_9286, wire_9247, wire_9246};
    // IPIN TOTAL: 276
    assign lut_tile_9_2_ipin_in = {wire_9357, wire_9356, wire_9337, wire_9336, wire_9317, wire_9316, wire_9297, wire_9296, wire_9277, wire_9276, wire_9257, wire_9256, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9743, wire_9742, wire_9703, wire_9702, wire_9663, wire_9662, wire_11159, wire_11158, wire_11149, wire_11148, wire_11139, wire_11138, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_9353, wire_9352, wire_9333, wire_9332, wire_9313, wire_9312, wire_9293, wire_9292, wire_9273, wire_9272, wire_9253, wire_9252, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9719, wire_9718, wire_9679, wire_9678, wire_9639, wire_9638, wire_11153, wire_11152, wire_11143, wire_11142, wire_11133, wire_11132, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_9737, wire_9736, wire_9725, wire_9724, wire_9697, wire_9696, wire_9685, wire_9684, wire_9657, wire_9656, wire_9645, wire_9644, wire_11157, wire_11156, wire_11147, wire_11146, wire_11137, wire_11136, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9335, wire_9334, wire_9295, wire_9294, wire_9255, wire_9254, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_9741, wire_9740, wire_9713, wire_9712, wire_9701, wire_9700, wire_9673, wire_9672, wire_9661, wire_9660, wire_9633, wire_9632, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9351, wire_9350, wire_9311, wire_9310, wire_9271, wire_9270, wire_11547, wire_11546, wire_11537, wire_11536, wire_11527, wire_11526, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_9729, wire_9728, wire_9717, wire_9716, wire_9689, wire_9688, wire_9677, wire_9676, wire_9649, wire_9648, wire_9637, wire_9636, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9327, wire_9326, wire_9287, wire_9286, wire_9247, wire_9246, wire_11541, wire_11540, wire_11531, wire_11530, wire_11521, wire_11520, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9727, wire_9726, wire_9687, wire_9686, wire_9647, wire_9646};
    // IPIN TOTAL: 276
    assign lut_tile_10_2_ipin_in = {wire_9745, wire_9744, wire_9733, wire_9732, wire_9705, wire_9704, wire_9693, wire_9692, wire_9665, wire_9664, wire_9653, wire_9652, wire_11545, wire_11544, wire_11535, wire_11534, wire_11525, wire_11524, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_10169, wire_10168, wire_10159, wire_10158, wire_10149, wire_10148, wire_10119, wire_10118, wire_10079, wire_10078, wire_10039, wire_10038, wire_11185, wire_11184, wire_11175, wire_11174, wire_11165, wire_11164, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_9749, wire_9748, wire_9721, wire_9720, wire_9709, wire_9708, wire_9681, wire_9680, wire_9669, wire_9668, wire_9641, wire_9640, wire_11549, wire_11548, wire_11539, wire_11538, wire_11529, wire_11528, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_10163, wire_10162, wire_10153, wire_10152, wire_10143, wire_10142, wire_10135, wire_10134, wire_10095, wire_10094, wire_10055, wire_10054, wire_11189, wire_11188, wire_11179, wire_11178, wire_11169, wire_11168, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9719, wire_9718, wire_9679, wire_9678, wire_9639, wire_9638, wire_11543, wire_11542, wire_11533, wire_11532, wire_11523, wire_11522, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_10125, wire_10124, wire_10113, wire_10112, wire_10085, wire_10084, wire_10073, wire_10072, wire_10045, wire_10044, wire_10033, wire_10032, wire_11183, wire_11182, wire_11173, wire_11172, wire_11163, wire_11162, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9735, wire_9734, wire_9695, wire_9694, wire_9655, wire_9654, wire_11547, wire_11546, wire_11537, wire_11536, wire_11527, wire_11526, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_10129, wire_10128, wire_10101, wire_10100, wire_10089, wire_10088, wire_10061, wire_10060, wire_10049, wire_10048, wire_10021, wire_10020, wire_11151, wire_11150, wire_11141, wire_11140, wire_11131, wire_11130, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9711, wire_9710, wire_9671, wire_9670, wire_9631, wire_9630, wire_11571, wire_11570, wire_11561, wire_11560, wire_11551, wire_11550, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_10117, wire_10116, wire_10105, wire_10104, wire_10077, wire_10076, wire_10065, wire_10064, wire_10037, wire_10036, wire_10025, wire_10024, wire_11155, wire_11154, wire_11145, wire_11144, wire_11135, wire_11134, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9727, wire_9726, wire_9687, wire_9686, wire_9647, wire_9646, wire_11575, wire_11574, wire_11565, wire_11564, wire_11555, wire_11554, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10103, wire_10102, wire_10063, wire_10062, wire_10023, wire_10022};
    // IPIN TOTAL: 276
    assign lut_tile_1_3_ipin_in = {wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_6223, wire_6222, wire_6183, wire_6182, wire_6143, wire_6142, wire_11693, wire_11692, wire_11681, wire_11680, wire_11653, wire_11652, wire_11641, wire_11640, wire_11613, wire_11612, wire_11601, wire_11600, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6609, wire_6608, wire_6569, wire_6568, wire_6529, wire_6528, wire_11303, wire_11302, wire_11291, wire_11290, wire_11263, wire_11262, wire_11251, wire_11250, wire_11223, wire_11222, wire_11211, wire_11210, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_6239, wire_6238, wire_6199, wire_6198, wire_6159, wire_6158, wire_11697, wire_11696, wire_11669, wire_11668, wire_11657, wire_11656, wire_11629, wire_11628, wire_11617, wire_11616, wire_11589, wire_11588, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_11307, wire_11306, wire_11279, wire_11278, wire_11267, wire_11266, wire_11239, wire_11238, wire_11227, wire_11226, wire_11199, wire_11198, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_6209, wire_6208, wire_6169, wire_6168, wire_6129, wire_6128, wire_11685, wire_11684, wire_11673, wire_11672, wire_11645, wire_11644, wire_11633, wire_11632, wire_11605, wire_11604, wire_11593, wire_11592, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6615, wire_6614, wire_6575, wire_6574, wire_6535, wire_6534, wire_11295, wire_11294, wire_11283, wire_11282, wire_11255, wire_11254, wire_11243, wire_11242, wire_11215, wire_11214, wire_11203, wire_11202, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_6225, wire_6224, wire_6185, wire_6184, wire_6145, wire_6144, wire_11689, wire_11688, wire_11661, wire_11660, wire_11649, wire_11648, wire_11621, wire_11620, wire_11609, wire_11608, wire_11581, wire_11580, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6591, wire_6590, wire_6551, wire_6550, wire_6511, wire_6510, wire_11301, wire_11300, wire_11273, wire_11272, wire_11261, wire_11260, wire_11233, wire_11232, wire_11221, wire_11220, wire_11193, wire_11192, wire_6297, wire_6296, wire_6287, wire_6286, wire_6277, wire_6276, wire_6201, wire_6200, wire_6161, wire_6160, wire_6121, wire_6120, wire_11687, wire_11686, wire_11667, wire_11666, wire_11647, wire_11646, wire_11627, wire_11626, wire_11607, wire_11606, wire_11587, wire_11586, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6607, wire_6606, wire_6567, wire_6566, wire_6527, wire_6526, wire_11289, wire_11288, wire_11277, wire_11276, wire_11249, wire_11248, wire_11237, wire_11236, wire_11209, wire_11208, wire_11197, wire_11196, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_6217, wire_6216, wire_6177, wire_6176, wire_6137, wire_6136, wire_11683, wire_11682, wire_11663, wire_11662, wire_11643, wire_11642, wire_11623, wire_11622, wire_11603, wire_11602, wire_11583, wire_11582, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512};
    // IPIN TOTAL: 276
    assign lut_tile_2_3_ipin_in = {wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6623, wire_6622, wire_6583, wire_6582, wire_6543, wire_6542, wire_11699, wire_11698, wire_11679, wire_11678, wire_11659, wire_11658, wire_11639, wire_11638, wire_11619, wire_11618, wire_11599, wire_11598, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11289, wire_11288, wire_11249, wire_11248, wire_11209, wire_11208, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6599, wire_6598, wire_6559, wire_6558, wire_6519, wire_6518, wire_11695, wire_11694, wire_11675, wire_11674, wire_11655, wire_11654, wire_11635, wire_11634, wire_11615, wire_11614, wire_11595, wire_11594, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_6993, wire_6992, wire_6953, wire_6952, wire_6913, wire_6912, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11305, wire_11304, wire_11265, wire_11264, wire_11225, wire_11224, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_11691, wire_11690, wire_11671, wire_11670, wire_11651, wire_11650, wire_11631, wire_11630, wire_11611, wire_11610, wire_11591, wire_11590, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6991, wire_6990, wire_6951, wire_6950, wire_6911, wire_6910, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11281, wire_11280, wire_11241, wire_11240, wire_11201, wire_11200, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6601, wire_6600, wire_6561, wire_6560, wire_6521, wire_6520, wire_11687, wire_11686, wire_11667, wire_11666, wire_11647, wire_11646, wire_11627, wire_11626, wire_11607, wire_11606, wire_11587, wire_11586, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_7007, wire_7006, wire_6967, wire_6966, wire_6927, wire_6926, wire_11299, wire_11298, wire_11271, wire_11270, wire_11259, wire_11258, wire_11231, wire_11230, wire_11219, wire_11218, wire_11191, wire_11190, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6617, wire_6616, wire_6577, wire_6576, wire_6537, wire_6536, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6983, wire_6982, wire_6943, wire_6942, wire_6903, wire_6902, wire_11287, wire_11286, wire_11275, wire_11274, wire_11247, wire_11246, wire_11235, wire_11234, wire_11207, wire_11206, wire_11195, wire_11194, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11681, wire_11680, wire_11641, wire_11640, wire_11601, wire_11600, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_7001, wire_7000, wire_6961, wire_6960, wire_6921, wire_6920};
    // IPIN TOTAL: 276
    assign lut_tile_3_3_ipin_in = {wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6999, wire_6998, wire_6959, wire_6958, wire_6919, wire_6918, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11697, wire_11696, wire_11657, wire_11656, wire_11617, wire_11616, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7393, wire_7392, wire_7353, wire_7352, wire_7313, wire_7312, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11307, wire_11306, wire_11267, wire_11266, wire_11227, wire_11226, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11673, wire_11672, wire_11633, wire_11632, wire_11593, wire_11592, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11283, wire_11282, wire_11243, wire_11242, wire_11203, wire_11202, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_6993, wire_6992, wire_6953, wire_6952, wire_6913, wire_6912, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11689, wire_11688, wire_11649, wire_11648, wire_11609, wire_11608, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7399, wire_7398, wire_7359, wire_7358, wire_7319, wire_7318, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11299, wire_11298, wire_11259, wire_11258, wire_11219, wire_11218, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_7009, wire_7008, wire_6969, wire_6968, wire_6929, wire_6928, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7375, wire_7374, wire_7335, wire_7334, wire_7295, wire_7294, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11297, wire_11296, wire_11257, wire_11256, wire_11217, wire_11216, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6985, wire_6984, wire_6945, wire_6944, wire_6905, wire_6904, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7391, wire_7390, wire_7351, wire_7350, wire_7311, wire_7310, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11273, wire_11272, wire_11233, wire_11232, wire_11193, wire_11192, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_7001, wire_7000, wire_6961, wire_6960, wire_6921, wire_6920, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11667, wire_11666, wire_11627, wire_11626, wire_11587, wire_11586, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296};
    // IPIN TOTAL: 276
    assign lut_tile_4_3_ipin_in = {wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7407, wire_7406, wire_7367, wire_7366, wire_7327, wire_7326, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11683, wire_11682, wire_11643, wire_11642, wire_11603, wire_11602, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7793, wire_7792, wire_7753, wire_7752, wire_7713, wire_7712, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7383, wire_7382, wire_7343, wire_7342, wire_7303, wire_7302, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11699, wire_11698, wire_11659, wire_11658, wire_11619, wire_11618, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11675, wire_11674, wire_11635, wire_11634, wire_11595, wire_11594, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7775, wire_7774, wire_7735, wire_7734, wire_7695, wire_7694, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7385, wire_7384, wire_7345, wire_7344, wire_7305, wire_7304, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7791, wire_7790, wire_7751, wire_7750, wire_7711, wire_7710, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7401, wire_7400, wire_7361, wire_7360, wire_7321, wire_7320, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7767, wire_7766, wire_7727, wire_7726, wire_7687, wire_7686, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11291, wire_11290, wire_11251, wire_11250, wire_11211, wire_11210, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7777, wire_7776, wire_7737, wire_7736, wire_7697, wire_7696};
    // IPIN TOTAL: 276
    assign lut_tile_5_3_ipin_in = {wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7783, wire_7782, wire_7743, wire_7742, wire_7703, wire_7702, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8169, wire_8168, wire_8129, wire_8128, wire_8089, wire_8088, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8175, wire_8174, wire_8135, wire_8134, wire_8095, wire_8094, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7785, wire_7784, wire_7745, wire_7744, wire_7705, wire_7704, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8151, wire_8150, wire_8111, wire_8110, wire_8071, wire_8070, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7761, wire_7760, wire_7721, wire_7720, wire_7681, wire_7680, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8167, wire_8166, wire_8127, wire_8126, wire_8087, wire_8086, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7777, wire_7776, wire_7737, wire_7736, wire_7697, wire_7696, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072};
    // IPIN TOTAL: 276
    assign lut_tile_6_3_ipin_in = {wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8183, wire_8182, wire_8143, wire_8142, wire_8103, wire_8102, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8159, wire_8158, wire_8119, wire_8118, wire_8079, wire_8078, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8553, wire_8552, wire_8513, wire_8512, wire_8473, wire_8472, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8551, wire_8550, wire_8511, wire_8510, wire_8471, wire_8470, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8161, wire_8160, wire_8121, wire_8120, wire_8081, wire_8080, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8567, wire_8566, wire_8527, wire_8526, wire_8487, wire_8486, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8177, wire_8176, wire_8137, wire_8136, wire_8097, wire_8096, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8543, wire_8542, wire_8503, wire_8502, wire_8463, wire_8462, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8561, wire_8560, wire_8521, wire_8520, wire_8481, wire_8480};
    // IPIN TOTAL: 276
    assign lut_tile_7_3_ipin_in = {wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8559, wire_8558, wire_8519, wire_8518, wire_8479, wire_8478, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8953, wire_8952, wire_8913, wire_8912, wire_8873, wire_8872, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8553, wire_8552, wire_8513, wire_8512, wire_8473, wire_8472, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8959, wire_8958, wire_8919, wire_8918, wire_8879, wire_8878, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8569, wire_8568, wire_8529, wire_8528, wire_8489, wire_8488, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8935, wire_8934, wire_8895, wire_8894, wire_8855, wire_8854, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8545, wire_8544, wire_8505, wire_8504, wire_8465, wire_8464, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8951, wire_8950, wire_8911, wire_8910, wire_8871, wire_8870, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8561, wire_8560, wire_8521, wire_8520, wire_8481, wire_8480, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856};
    // IPIN TOTAL: 276
    assign lut_tile_8_3_ipin_in = {wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8967, wire_8966, wire_8927, wire_8926, wire_8887, wire_8886, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9353, wire_9352, wire_9313, wire_9312, wire_9273, wire_9272, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8943, wire_8942, wire_8903, wire_8902, wire_8863, wire_8862, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9335, wire_9334, wire_9295, wire_9294, wire_9255, wire_9254, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8945, wire_8944, wire_8905, wire_8904, wire_8865, wire_8864, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9351, wire_9350, wire_9311, wire_9310, wire_9271, wire_9270, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8961, wire_8960, wire_8921, wire_8920, wire_8881, wire_8880, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9327, wire_9326, wire_9287, wire_9286, wire_9247, wire_9246, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9337, wire_9336, wire_9297, wire_9296, wire_9257, wire_9256};
    // IPIN TOTAL: 276
    assign lut_tile_9_3_ipin_in = {wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9343, wire_9342, wire_9303, wire_9302, wire_9263, wire_9262, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9729, wire_9728, wire_9689, wire_9688, wire_9649, wire_9648, wire_11545, wire_11544, wire_11535, wire_11534, wire_11525, wire_11524, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_11549, wire_11548, wire_11539, wire_11538, wire_11529, wire_11528, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9735, wire_9734, wire_9695, wire_9694, wire_9655, wire_9654, wire_11543, wire_11542, wire_11533, wire_11532, wire_11523, wire_11522, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9345, wire_9344, wire_9305, wire_9304, wire_9265, wire_9264, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9711, wire_9710, wire_9671, wire_9670, wire_9631, wire_9630, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9321, wire_9320, wire_9281, wire_9280, wire_9241, wire_9240, wire_11931, wire_11930, wire_11921, wire_11920, wire_11911, wire_11910, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9727, wire_9726, wire_9687, wire_9686, wire_9647, wire_9646, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9337, wire_9336, wire_9297, wire_9296, wire_9257, wire_9256, wire_11935, wire_11934, wire_11925, wire_11924, wire_11915, wire_11914, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632};
    // IPIN TOTAL: 276
    assign lut_tile_10_3_ipin_in = {wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9743, wire_9742, wire_9703, wire_9702, wire_9663, wire_9662, wire_11939, wire_11938, wire_11929, wire_11928, wire_11919, wire_11918, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174, wire_10137, wire_10136, wire_10097, wire_10096, wire_10057, wire_10056, wire_11579, wire_11578, wire_11569, wire_11568, wire_11559, wire_11558, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9719, wire_9718, wire_9679, wire_9678, wire_9639, wire_9638, wire_11933, wire_11932, wire_11923, wire_11922, wire_11913, wire_11912, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_10199, wire_10198, wire_10189, wire_10188, wire_10179, wire_10178, wire_10113, wire_10112, wire_10073, wire_10072, wire_10033, wire_10032, wire_11573, wire_11572, wire_11563, wire_11562, wire_11553, wire_11552, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_11937, wire_11936, wire_11927, wire_11926, wire_11917, wire_11916, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_10167, wire_10166, wire_10157, wire_10156, wire_10147, wire_10146, wire_10111, wire_10110, wire_10071, wire_10070, wire_10031, wire_10030, wire_11577, wire_11576, wire_11567, wire_11566, wire_11557, wire_11556, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9721, wire_9720, wire_9681, wire_9680, wire_9641, wire_9640, wire_11931, wire_11930, wire_11921, wire_11920, wire_11911, wire_11910, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140, wire_10127, wire_10126, wire_10087, wire_10086, wire_10047, wire_10046, wire_11547, wire_11546, wire_11537, wire_11536, wire_11527, wire_11526, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9737, wire_9736, wire_9697, wire_9696, wire_9657, wire_9656, wire_11967, wire_11966, wire_11957, wire_11956, wire_11947, wire_11946, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10103, wire_10102, wire_10063, wire_10062, wire_10023, wire_10022, wire_11541, wire_11540, wire_11531, wire_11530, wire_11521, wire_11520, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632, wire_11961, wire_11960, wire_11951, wire_11950, wire_11941, wire_11940, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_10121, wire_10120, wire_10081, wire_10080, wire_10041, wire_10040};
    // IPIN TOTAL: 276
    assign lut_tile_1_4_ipin_in = {wire_6295, wire_6294, wire_6285, wire_6284, wire_6275, wire_6274, wire_6233, wire_6232, wire_6193, wire_6192, wire_6153, wire_6152, wire_12089, wire_12088, wire_12069, wire_12068, wire_12049, wire_12048, wire_12029, wire_12028, wire_12009, wire_12008, wire_11989, wire_11988, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_11699, wire_11698, wire_11679, wire_11678, wire_11659, wire_11658, wire_11639, wire_11638, wire_11619, wire_11618, wire_11599, wire_11598, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_6209, wire_6208, wire_6169, wire_6168, wire_6129, wire_6128, wire_12085, wire_12084, wire_12065, wire_12064, wire_12045, wire_12044, wire_12025, wire_12024, wire_12005, wire_12004, wire_11985, wire_11984, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_11695, wire_11694, wire_11675, wire_11674, wire_11655, wire_11654, wire_11635, wire_11634, wire_11615, wire_11614, wire_11595, wire_11594, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_12081, wire_12080, wire_12061, wire_12060, wire_12041, wire_12040, wire_12021, wire_12020, wire_12001, wire_12000, wire_11981, wire_11980, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6601, wire_6600, wire_6561, wire_6560, wire_6521, wire_6520, wire_11691, wire_11690, wire_11671, wire_11670, wire_11651, wire_11650, wire_11631, wire_11630, wire_11611, wire_11610, wire_11591, wire_11590, wire_6327, wire_6326, wire_6317, wire_6316, wire_6307, wire_6306, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_12077, wire_12076, wire_12057, wire_12056, wire_12037, wire_12036, wire_12017, wire_12016, wire_11997, wire_11996, wire_11977, wire_11976, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6617, wire_6616, wire_6577, wire_6576, wire_6537, wire_6536, wire_11689, wire_11688, wire_11661, wire_11660, wire_11649, wire_11648, wire_11621, wire_11620, wire_11609, wire_11608, wire_11581, wire_11580, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300, wire_6267, wire_6266, wire_6257, wire_6256, wire_6247, wire_6246, wire_12075, wire_12074, wire_12055, wire_12054, wire_12035, wire_12034, wire_12015, wire_12014, wire_11995, wire_11994, wire_11975, wire_11974, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512, wire_11677, wire_11676, wire_11665, wire_11664, wire_11637, wire_11636, wire_11625, wire_11624, wire_11597, wire_11596, wire_11585, wire_11584, wire_6325, wire_6324, wire_6315, wire_6314, wire_6305, wire_6304, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240, wire_12071, wire_12070, wire_12051, wire_12050, wire_12031, wire_12030, wire_12011, wire_12010, wire_11991, wire_11990, wire_11971, wire_11970, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634};
    // IPIN TOTAL: 276
    assign lut_tile_2_4_ipin_in = {wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6609, wire_6608, wire_6569, wire_6568, wire_6529, wire_6528, wire_12087, wire_12086, wire_12067, wire_12066, wire_12047, wire_12046, wire_12027, wire_12026, wire_12007, wire_12006, wire_11987, wire_11986, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11697, wire_11696, wire_11657, wire_11656, wire_11617, wire_11616, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_12083, wire_12082, wire_12063, wire_12062, wire_12043, wire_12042, wire_12023, wire_12022, wire_12003, wire_12002, wire_11983, wire_11982, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11673, wire_11672, wire_11633, wire_11632, wire_11593, wire_11592, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_12079, wire_12078, wire_12059, wire_12058, wire_12039, wire_12038, wire_12019, wire_12018, wire_11999, wire_11998, wire_11979, wire_11978, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_7009, wire_7008, wire_6969, wire_6968, wire_6929, wire_6928, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11689, wire_11688, wire_11649, wire_11648, wire_11609, wire_11608, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_12075, wire_12074, wire_12055, wire_12054, wire_12035, wire_12034, wire_12015, wire_12014, wire_11995, wire_11994, wire_11975, wire_11974, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6985, wire_6984, wire_6945, wire_6944, wire_6905, wire_6904, wire_11687, wire_11686, wire_11667, wire_11666, wire_11647, wire_11646, wire_11627, wire_11626, wire_11607, wire_11606, wire_11587, wire_11586, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12081, wire_12080, wire_12041, wire_12040, wire_12001, wire_12000, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_7001, wire_7000, wire_6961, wire_6960, wire_6921, wire_6920, wire_11683, wire_11682, wire_11663, wire_11662, wire_11643, wire_11642, wire_11623, wire_11622, wire_11603, wire_11602, wire_11583, wire_11582, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12057, wire_12056, wire_12017, wire_12016, wire_11977, wire_11976, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020};
    // IPIN TOTAL: 276
    assign lut_tile_3_4_ipin_in = {wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_12073, wire_12072, wire_12033, wire_12032, wire_11993, wire_11992, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11683, wire_11682, wire_11643, wire_11642, wire_11603, wire_11602, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_6993, wire_6992, wire_6953, wire_6952, wire_6913, wire_6912, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12089, wire_12088, wire_12049, wire_12048, wire_12009, wire_12008, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11699, wire_11698, wire_11659, wire_11658, wire_11619, wire_11618, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12065, wire_12064, wire_12025, wire_12024, wire_11985, wire_11984, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7385, wire_7384, wire_7345, wire_7344, wire_7305, wire_7304, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11675, wire_11674, wire_11635, wire_11634, wire_11595, wire_11594, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12081, wire_12080, wire_12041, wire_12040, wire_12001, wire_12000, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7401, wire_7400, wire_7361, wire_7360, wire_7321, wire_7320, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11681, wire_11680, wire_11641, wire_11640, wire_11601, wire_11600, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12067, wire_12066, wire_12027, wire_12026, wire_11987, wire_11986, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414};
    // IPIN TOTAL: 276
    assign lut_tile_4_4_ipin_in = {wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7393, wire_7392, wire_7353, wire_7352, wire_7313, wire_7312, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12083, wire_12082, wire_12043, wire_12042, wire_12003, wire_12002, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12059, wire_12058, wire_12019, wire_12018, wire_11979, wire_11978, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12075, wire_12074, wire_12035, wire_12034, wire_11995, wire_11994, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7785, wire_7784, wire_7745, wire_7744, wire_7705, wire_7704, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7761, wire_7760, wire_7721, wire_7720, wire_7681, wire_7680, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7777, wire_7776, wire_7737, wire_7736, wire_7697, wire_7696, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11667, wire_11666, wire_11627, wire_11626, wire_11587, wire_11586, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800};
    // IPIN TOTAL: 276
    assign lut_tile_5_4_ipin_in = {wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7793, wire_7792, wire_7753, wire_7752, wire_7713, wire_7712, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8161, wire_8160, wire_8121, wire_8120, wire_8081, wire_8080, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8177, wire_8176, wire_8137, wire_8136, wire_8097, wire_8096, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194};
    // IPIN TOTAL: 276
    assign lut_tile_6_4_ipin_in = {wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8169, wire_8168, wire_8129, wire_8128, wire_8089, wire_8088, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8569, wire_8568, wire_8529, wire_8528, wire_8489, wire_8488, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8545, wire_8544, wire_8505, wire_8504, wire_8465, wire_8464, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8561, wire_8560, wire_8521, wire_8520, wire_8481, wire_8480, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580};
    // IPIN TOTAL: 276
    assign lut_tile_7_4_ipin_in = {wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8553, wire_8552, wire_8513, wire_8512, wire_8473, wire_8472, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8945, wire_8944, wire_8905, wire_8904, wire_8865, wire_8864, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8961, wire_8960, wire_8921, wire_8920, wire_8881, wire_8880, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974};
    // IPIN TOTAL: 276
    assign lut_tile_8_4_ipin_in = {wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8953, wire_8952, wire_8913, wire_8912, wire_8873, wire_8872, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9345, wire_9344, wire_9305, wire_9304, wire_9265, wire_9264, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9321, wire_9320, wire_9281, wire_9280, wire_9241, wire_9240, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9337, wire_9336, wire_9297, wire_9296, wire_9257, wire_9256, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360};
    // IPIN TOTAL: 276
    assign lut_tile_9_4_ipin_in = {wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9353, wire_9352, wire_9313, wire_9312, wire_9273, wire_9272, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_11939, wire_11938, wire_11929, wire_11928, wire_11919, wire_11918, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_11933, wire_11932, wire_11923, wire_11922, wire_11913, wire_11912, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9721, wire_9720, wire_9681, wire_9680, wire_9641, wire_9640, wire_11937, wire_11936, wire_11927, wire_11926, wire_11917, wire_11916, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9737, wire_9736, wire_9697, wire_9696, wire_9657, wire_9656, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_12327, wire_12326, wire_12317, wire_12316, wire_12307, wire_12306, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_12321, wire_12320, wire_12311, wire_12310, wire_12301, wire_12300, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754};
    // IPIN TOTAL: 276
    assign lut_tile_10_4_ipin_in = {wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9729, wire_9728, wire_9689, wire_9688, wire_9649, wire_9648, wire_12325, wire_12324, wire_12315, wire_12314, wire_12305, wire_12304, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_10229, wire_10228, wire_10219, wire_10218, wire_10209, wire_10208, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_11965, wire_11964, wire_11955, wire_11954, wire_11945, wire_11944, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_12329, wire_12328, wire_12319, wire_12318, wire_12309, wire_12308, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_10223, wire_10222, wire_10213, wire_10212, wire_10203, wire_10202, wire_10169, wire_10168, wire_10159, wire_10158, wire_10149, wire_10148, wire_11969, wire_11968, wire_11959, wire_11958, wire_11949, wire_11948, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_12323, wire_12322, wire_12313, wire_12312, wire_12303, wire_12302, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_10193, wire_10192, wire_10183, wire_10182, wire_10173, wire_10172, wire_10129, wire_10128, wire_10089, wire_10088, wire_10049, wire_10048, wire_11963, wire_11962, wire_11953, wire_11952, wire_11943, wire_11942, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_12327, wire_12326, wire_12317, wire_12316, wire_12307, wire_12306, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_10197, wire_10196, wire_10187, wire_10186, wire_10177, wire_10176, wire_10105, wire_10104, wire_10065, wire_10064, wire_10025, wire_10024, wire_11931, wire_11930, wire_11921, wire_11920, wire_11911, wire_11910, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_12351, wire_12350, wire_12341, wire_12340, wire_12331, wire_12330, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_10121, wire_10120, wire_10081, wire_10080, wire_10041, wire_10040, wire_11935, wire_11934, wire_11925, wire_11924, wire_11915, wire_11914, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_12355, wire_12354, wire_12345, wire_12344, wire_12335, wire_12334, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140};
    // IPIN TOTAL: 276
    assign lut_tile_1_5_ipin_in = {wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_6265, wire_6264, wire_6255, wire_6254, wire_6245, wire_6244, wire_12477, wire_12476, wire_12457, wire_12456, wire_12437, wire_12436, wire_12417, wire_12416, wire_12397, wire_12396, wire_12377, wire_12376, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_12087, wire_12086, wire_12067, wire_12066, wire_12047, wire_12046, wire_12027, wire_12026, wire_12007, wire_12006, wire_11987, wire_11986, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_12473, wire_12472, wire_12453, wire_12452, wire_12433, wire_12432, wire_12413, wire_12412, wire_12393, wire_12392, wire_12373, wire_12372, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_12083, wire_12082, wire_12063, wire_12062, wire_12043, wire_12042, wire_12023, wire_12022, wire_12003, wire_12002, wire_11983, wire_11982, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_12469, wire_12468, wire_12449, wire_12448, wire_12429, wire_12428, wire_12409, wire_12408, wire_12389, wire_12388, wire_12369, wire_12368, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_12079, wire_12078, wire_12059, wire_12058, wire_12039, wire_12038, wire_12019, wire_12018, wire_11999, wire_11998, wire_11979, wire_11978, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_6297, wire_6296, wire_6287, wire_6286, wire_6277, wire_6276, wire_12465, wire_12464, wire_12445, wire_12444, wire_12425, wire_12424, wire_12405, wire_12404, wire_12385, wire_12384, wire_12365, wire_12364, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_12077, wire_12076, wire_12057, wire_12056, wire_12037, wire_12036, wire_12017, wire_12016, wire_11997, wire_11996, wire_11977, wire_11976, wire_6357, wire_6356, wire_6347, wire_6346, wire_6337, wire_6336, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_12471, wire_12470, wire_12443, wire_12442, wire_12431, wire_12430, wire_12403, wire_12402, wire_12391, wire_12390, wire_12363, wire_12362, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_12073, wire_12072, wire_12053, wire_12052, wire_12033, wire_12032, wire_12013, wire_12012, wire_11993, wire_11992, wire_11973, wire_11972, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_6295, wire_6294, wire_6285, wire_6284, wire_6275, wire_6274, wire_12459, wire_12458, wire_12447, wire_12446, wire_12419, wire_12418, wire_12407, wire_12406, wire_12379, wire_12378, wire_12367, wire_12366, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660};
    // IPIN TOTAL: 276
    assign lut_tile_2_5_ipin_in = {wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_12475, wire_12474, wire_12463, wire_12462, wire_12435, wire_12434, wire_12423, wire_12422, wire_12395, wire_12394, wire_12383, wire_12382, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_12073, wire_12072, wire_12033, wire_12032, wire_11993, wire_11992, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_12479, wire_12478, wire_12451, wire_12450, wire_12439, wire_12438, wire_12411, wire_12410, wire_12399, wire_12398, wire_12371, wire_12370, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12089, wire_12088, wire_12049, wire_12048, wire_12009, wire_12008, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_12467, wire_12466, wire_12455, wire_12454, wire_12427, wire_12426, wire_12415, wire_12414, wire_12387, wire_12386, wire_12375, wire_12374, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12065, wire_12064, wire_12025, wire_12024, wire_11985, wire_11984, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_12471, wire_12470, wire_12443, wire_12442, wire_12431, wire_12430, wire_12403, wire_12402, wire_12391, wire_12390, wire_12363, wire_12362, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_12075, wire_12074, wire_12055, wire_12054, wire_12035, wire_12034, wire_12015, wire_12014, wire_11995, wire_11994, wire_11975, wire_11974, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_12071, wire_12070, wire_12051, wire_12050, wire_12031, wire_12030, wire_12011, wire_12010, wire_11991, wire_11990, wire_11971, wire_11970, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12457, wire_12456, wire_12417, wire_12416, wire_12377, wire_12376, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054};
    // IPIN TOTAL: 276
    assign lut_tile_3_5_ipin_in = {wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12473, wire_12472, wire_12433, wire_12432, wire_12393, wire_12392, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12083, wire_12082, wire_12043, wire_12042, wire_12003, wire_12002, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12449, wire_12448, wire_12409, wire_12408, wire_12369, wire_12368, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12059, wire_12058, wire_12019, wire_12018, wire_11979, wire_11978, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12465, wire_12464, wire_12425, wire_12424, wire_12385, wire_12384, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12075, wire_12074, wire_12035, wire_12034, wire_11995, wire_11994, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12081, wire_12080, wire_12041, wire_12040, wire_12001, wire_12000, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12467, wire_12466, wire_12427, wire_12426, wire_12387, wire_12386, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12057, wire_12056, wire_12017, wire_12016, wire_11977, wire_11976, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440};
    // IPIN TOTAL: 276
    assign lut_tile_4_5_ipin_in = {wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12459, wire_12458, wire_12419, wire_12418, wire_12379, wire_12378, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12475, wire_12474, wire_12435, wire_12434, wire_12395, wire_12394, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12451, wire_12450, wire_12411, wire_12410, wire_12371, wire_12370, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12467, wire_12466, wire_12427, wire_12426, wire_12387, wire_12386, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12067, wire_12066, wire_12027, wire_12026, wire_11987, wire_11986, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834};
    // IPIN TOTAL: 276
    assign lut_tile_5_5_ipin_in = {wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220};
    // IPIN TOTAL: 276
    assign lut_tile_6_5_ipin_in = {wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614};
    // IPIN TOTAL: 276
    assign lut_tile_7_5_ipin_in = {wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000};
    // IPIN TOTAL: 276
    assign lut_tile_8_5_ipin_in = {wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394};
    // IPIN TOTAL: 276
    assign lut_tile_9_5_ipin_in = {wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_12325, wire_12324, wire_12315, wire_12314, wire_12305, wire_12304, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_12329, wire_12328, wire_12319, wire_12318, wire_12309, wire_12308, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_12323, wire_12322, wire_12313, wire_12312, wire_12303, wire_12302, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_12711, wire_12710, wire_12701, wire_12700, wire_12691, wire_12690, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_12715, wire_12714, wire_12705, wire_12704, wire_12695, wire_12694, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780};
    // IPIN TOTAL: 276
    assign lut_tile_10_5_ipin_in = {wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_12719, wire_12718, wire_12709, wire_12708, wire_12699, wire_12698, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234, wire_10199, wire_10198, wire_10189, wire_10188, wire_10179, wire_10178, wire_12359, wire_12358, wire_12349, wire_12348, wire_12339, wire_12338, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_12713, wire_12712, wire_12703, wire_12702, wire_12693, wire_12692, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_10259, wire_10258, wire_10249, wire_10248, wire_10239, wire_10238, wire_10193, wire_10192, wire_10183, wire_10182, wire_10173, wire_10172, wire_12353, wire_12352, wire_12343, wire_12342, wire_12333, wire_12332, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_12717, wire_12716, wire_12707, wire_12706, wire_12697, wire_12696, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_10227, wire_10226, wire_10217, wire_10216, wire_10207, wire_10206, wire_10163, wire_10162, wire_10153, wire_10152, wire_10143, wire_10142, wire_12357, wire_12356, wire_12347, wire_12346, wire_12337, wire_12336, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_12711, wire_12710, wire_12701, wire_12700, wire_12691, wire_12690, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200, wire_10167, wire_10166, wire_10157, wire_10156, wire_10147, wire_10146, wire_12327, wire_12326, wire_12317, wire_12316, wire_12307, wire_12306, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_12747, wire_12746, wire_12737, wire_12736, wire_12727, wire_12726, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140, wire_12321, wire_12320, wire_12311, wire_12310, wire_12301, wire_12300, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_12741, wire_12740, wire_12731, wire_12730, wire_12721, wire_12720, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174};
    // IPIN TOTAL: 276
    assign lut_tile_1_6_ipin_in = {wire_6355, wire_6354, wire_6345, wire_6344, wire_6335, wire_6334, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_12865, wire_12864, wire_12853, wire_12852, wire_12825, wire_12824, wire_12813, wire_12812, wire_12785, wire_12784, wire_12773, wire_12772, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_12475, wire_12474, wire_12463, wire_12462, wire_12435, wire_12434, wire_12423, wire_12422, wire_12395, wire_12394, wire_12383, wire_12382, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_12869, wire_12868, wire_12841, wire_12840, wire_12829, wire_12828, wire_12801, wire_12800, wire_12789, wire_12788, wire_12761, wire_12760, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_12479, wire_12478, wire_12451, wire_12450, wire_12439, wire_12438, wire_12411, wire_12410, wire_12399, wire_12398, wire_12371, wire_12370, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_12857, wire_12856, wire_12845, wire_12844, wire_12817, wire_12816, wire_12805, wire_12804, wire_12777, wire_12776, wire_12765, wire_12764, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_12467, wire_12466, wire_12455, wire_12454, wire_12427, wire_12426, wire_12415, wire_12414, wire_12387, wire_12386, wire_12375, wire_12374, wire_6387, wire_6386, wire_6377, wire_6376, wire_6367, wire_6366, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_12861, wire_12860, wire_12833, wire_12832, wire_12821, wire_12820, wire_12793, wire_12792, wire_12781, wire_12780, wire_12753, wire_12752, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_12465, wire_12464, wire_12445, wire_12444, wire_12425, wire_12424, wire_12405, wire_12404, wire_12385, wire_12384, wire_12365, wire_12364, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360, wire_6327, wire_6326, wire_6317, wire_6316, wire_6307, wire_6306, wire_12859, wire_12858, wire_12831, wire_12830, wire_12819, wire_12818, wire_12791, wire_12790, wire_12779, wire_12778, wire_12751, wire_12750, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_12461, wire_12460, wire_12441, wire_12440, wire_12421, wire_12420, wire_12401, wire_12400, wire_12381, wire_12380, wire_12361, wire_12360, wire_6385, wire_6384, wire_6375, wire_6374, wire_6365, wire_6364, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300, wire_12847, wire_12846, wire_12835, wire_12834, wire_12807, wire_12806, wire_12795, wire_12794, wire_12767, wire_12766, wire_12755, wire_12754, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694};
    // IPIN TOTAL: 276
    assign lut_tile_2_6_ipin_in = {wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_12863, wire_12862, wire_12851, wire_12850, wire_12823, wire_12822, wire_12811, wire_12810, wire_12783, wire_12782, wire_12771, wire_12770, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12473, wire_12472, wire_12433, wire_12432, wire_12393, wire_12392, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_12867, wire_12866, wire_12839, wire_12838, wire_12827, wire_12826, wire_12799, wire_12798, wire_12787, wire_12786, wire_12759, wire_12758, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12449, wire_12448, wire_12409, wire_12408, wire_12369, wire_12368, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_12855, wire_12854, wire_12843, wire_12842, wire_12815, wire_12814, wire_12803, wire_12802, wire_12775, wire_12774, wire_12763, wire_12762, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12465, wire_12464, wire_12425, wire_12424, wire_12385, wire_12384, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_12859, wire_12858, wire_12831, wire_12830, wire_12819, wire_12818, wire_12791, wire_12790, wire_12779, wire_12778, wire_12751, wire_12750, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_12471, wire_12470, wire_12443, wire_12442, wire_12431, wire_12430, wire_12403, wire_12402, wire_12391, wire_12390, wire_12363, wire_12362, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12857, wire_12856, wire_12817, wire_12816, wire_12777, wire_12776, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_12459, wire_12458, wire_12447, wire_12446, wire_12419, wire_12418, wire_12407, wire_12406, wire_12379, wire_12378, wire_12367, wire_12366, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12833, wire_12832, wire_12793, wire_12792, wire_12753, wire_12752, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080};
    // IPIN TOTAL: 276
    assign lut_tile_3_6_ipin_in = {wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12849, wire_12848, wire_12809, wire_12808, wire_12769, wire_12768, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12459, wire_12458, wire_12419, wire_12418, wire_12379, wire_12378, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12865, wire_12864, wire_12825, wire_12824, wire_12785, wire_12784, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12475, wire_12474, wire_12435, wire_12434, wire_12395, wire_12394, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12841, wire_12840, wire_12801, wire_12800, wire_12761, wire_12760, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12451, wire_12450, wire_12411, wire_12410, wire_12371, wire_12370, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12857, wire_12856, wire_12817, wire_12816, wire_12777, wire_12776, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12457, wire_12456, wire_12417, wire_12416, wire_12377, wire_12376, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12851, wire_12850, wire_12811, wire_12810, wire_12771, wire_12770, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474};
    // IPIN TOTAL: 276
    assign lut_tile_4_6_ipin_in = {wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12867, wire_12866, wire_12827, wire_12826, wire_12787, wire_12786, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12843, wire_12842, wire_12803, wire_12802, wire_12763, wire_12762, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12859, wire_12858, wire_12819, wire_12818, wire_12779, wire_12778, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12467, wire_12466, wire_12427, wire_12426, wire_12387, wire_12386, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860};
    // IPIN TOTAL: 276
    assign lut_tile_5_6_ipin_in = {wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254};
    // IPIN TOTAL: 276
    assign lut_tile_6_6_ipin_in = {wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640};
    // IPIN TOTAL: 276
    assign lut_tile_7_6_ipin_in = {wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034};
    // IPIN TOTAL: 276
    assign lut_tile_8_6_ipin_in = {wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420};
    // IPIN TOTAL: 276
    assign lut_tile_9_6_ipin_in = {wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_12719, wire_12718, wire_12709, wire_12708, wire_12699, wire_12698, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_12713, wire_12712, wire_12703, wire_12702, wire_12693, wire_12692, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_12717, wire_12716, wire_12707, wire_12706, wire_12697, wire_12696, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_13107, wire_13106, wire_13097, wire_13096, wire_13087, wire_13086, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_13101, wire_13100, wire_13091, wire_13090, wire_13081, wire_13080, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814};
    // IPIN TOTAL: 276
    assign lut_tile_10_6_ipin_in = {wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_13105, wire_13104, wire_13095, wire_13094, wire_13085, wire_13084, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_10289, wire_10288, wire_10279, wire_10278, wire_10269, wire_10268, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_12745, wire_12744, wire_12735, wire_12734, wire_12725, wire_12724, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_13109, wire_13108, wire_13099, wire_13098, wire_13089, wire_13088, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_10283, wire_10282, wire_10273, wire_10272, wire_10263, wire_10262, wire_10229, wire_10228, wire_10219, wire_10218, wire_10209, wire_10208, wire_12749, wire_12748, wire_12739, wire_12738, wire_12729, wire_12728, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_13103, wire_13102, wire_13093, wire_13092, wire_13083, wire_13082, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_10253, wire_10252, wire_10243, wire_10242, wire_10233, wire_10232, wire_10197, wire_10196, wire_10187, wire_10186, wire_10177, wire_10176, wire_12743, wire_12742, wire_12733, wire_12732, wire_12723, wire_12722, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_13107, wire_13106, wire_13097, wire_13096, wire_13087, wire_13086, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_10257, wire_10256, wire_10247, wire_10246, wire_10237, wire_10236, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_12711, wire_12710, wire_12701, wire_12700, wire_12691, wire_12690, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_13131, wire_13130, wire_13121, wire_13120, wire_13111, wire_13110, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174, wire_12715, wire_12714, wire_12705, wire_12704, wire_12695, wire_12694, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_13135, wire_13134, wire_13125, wire_13124, wire_13115, wire_13114, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200};
    // IPIN TOTAL: 276
    assign lut_tile_1_7_ipin_in = {wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_6325, wire_6324, wire_6315, wire_6314, wire_6305, wire_6304, wire_13253, wire_13252, wire_13241, wire_13240, wire_13213, wire_13212, wire_13201, wire_13200, wire_13173, wire_13172, wire_13161, wire_13160, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_12863, wire_12862, wire_12851, wire_12850, wire_12823, wire_12822, wire_12811, wire_12810, wire_12783, wire_12782, wire_12771, wire_12770, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_13257, wire_13256, wire_13229, wire_13228, wire_13217, wire_13216, wire_13189, wire_13188, wire_13177, wire_13176, wire_13149, wire_13148, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_12867, wire_12866, wire_12839, wire_12838, wire_12827, wire_12826, wire_12799, wire_12798, wire_12787, wire_12786, wire_12759, wire_12758, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_13245, wire_13244, wire_13233, wire_13232, wire_13205, wire_13204, wire_13193, wire_13192, wire_13165, wire_13164, wire_13153, wire_13152, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_12855, wire_12854, wire_12843, wire_12842, wire_12815, wire_12814, wire_12803, wire_12802, wire_12775, wire_12774, wire_12763, wire_12762, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_6357, wire_6356, wire_6347, wire_6346, wire_6337, wire_6336, wire_13249, wire_13248, wire_13221, wire_13220, wire_13209, wire_13208, wire_13181, wire_13180, wire_13169, wire_13168, wire_13141, wire_13140, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_12861, wire_12860, wire_12833, wire_12832, wire_12821, wire_12820, wire_12793, wire_12792, wire_12781, wire_12780, wire_12753, wire_12752, wire_6417, wire_6416, wire_6407, wire_6406, wire_6397, wire_6396, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_13247, wire_13246, wire_13227, wire_13226, wire_13207, wire_13206, wire_13187, wire_13186, wire_13167, wire_13166, wire_13147, wire_13146, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_12849, wire_12848, wire_12837, wire_12836, wire_12809, wire_12808, wire_12797, wire_12796, wire_12769, wire_12768, wire_12757, wire_12756, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_6355, wire_6354, wire_6345, wire_6344, wire_6335, wire_6334, wire_13243, wire_13242, wire_13223, wire_13222, wire_13203, wire_13202, wire_13183, wire_13182, wire_13163, wire_13162, wire_13143, wire_13142, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720};
    // IPIN TOTAL: 276
    assign lut_tile_2_7_ipin_in = {wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_13259, wire_13258, wire_13239, wire_13238, wire_13219, wire_13218, wire_13199, wire_13198, wire_13179, wire_13178, wire_13159, wire_13158, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12849, wire_12848, wire_12809, wire_12808, wire_12769, wire_12768, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_13255, wire_13254, wire_13235, wire_13234, wire_13215, wire_13214, wire_13195, wire_13194, wire_13175, wire_13174, wire_13155, wire_13154, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12865, wire_12864, wire_12825, wire_12824, wire_12785, wire_12784, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_13251, wire_13250, wire_13231, wire_13230, wire_13211, wire_13210, wire_13191, wire_13190, wire_13171, wire_13170, wire_13151, wire_13150, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12841, wire_12840, wire_12801, wire_12800, wire_12761, wire_12760, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_13247, wire_13246, wire_13227, wire_13226, wire_13207, wire_13206, wire_13187, wire_13186, wire_13167, wire_13166, wire_13147, wire_13146, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_12859, wire_12858, wire_12831, wire_12830, wire_12819, wire_12818, wire_12791, wire_12790, wire_12779, wire_12778, wire_12751, wire_12750, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_12847, wire_12846, wire_12835, wire_12834, wire_12807, wire_12806, wire_12795, wire_12794, wire_12767, wire_12766, wire_12755, wire_12754, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13241, wire_13240, wire_13201, wire_13200, wire_13161, wire_13160, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114};
    // IPIN TOTAL: 276
    assign lut_tile_3_7_ipin_in = {wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13257, wire_13256, wire_13217, wire_13216, wire_13177, wire_13176, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12867, wire_12866, wire_12827, wire_12826, wire_12787, wire_12786, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13233, wire_13232, wire_13193, wire_13192, wire_13153, wire_13152, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12843, wire_12842, wire_12803, wire_12802, wire_12763, wire_12762, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13249, wire_13248, wire_13209, wire_13208, wire_13169, wire_13168, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12859, wire_12858, wire_12819, wire_12818, wire_12779, wire_12778, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12857, wire_12856, wire_12817, wire_12816, wire_12777, wire_12776, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12833, wire_12832, wire_12793, wire_12792, wire_12753, wire_12752, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13227, wire_13226, wire_13187, wire_13186, wire_13147, wire_13146, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500};
    // IPIN TOTAL: 276
    assign lut_tile_4_7_ipin_in = {wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13243, wire_13242, wire_13203, wire_13202, wire_13163, wire_13162, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13259, wire_13258, wire_13219, wire_13218, wire_13179, wire_13178, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13235, wire_13234, wire_13195, wire_13194, wire_13155, wire_13154, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12851, wire_12850, wire_12811, wire_12810, wire_12771, wire_12770, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894};
    // IPIN TOTAL: 276
    assign lut_tile_5_7_ipin_in = {wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280};
    // IPIN TOTAL: 276
    assign lut_tile_6_7_ipin_in = {wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674};
    // IPIN TOTAL: 276
    assign lut_tile_7_7_ipin_in = {wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060};
    // IPIN TOTAL: 276
    assign lut_tile_8_7_ipin_in = {wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454};
    // IPIN TOTAL: 276
    assign lut_tile_9_7_ipin_in = {wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_13105, wire_13104, wire_13095, wire_13094, wire_13085, wire_13084, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_13109, wire_13108, wire_13099, wire_13098, wire_13089, wire_13088, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_13103, wire_13102, wire_13093, wire_13092, wire_13083, wire_13082, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_13491, wire_13490, wire_13481, wire_13480, wire_13471, wire_13470, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_13495, wire_13494, wire_13485, wire_13484, wire_13475, wire_13474, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840};
    // IPIN TOTAL: 276
    assign lut_tile_10_7_ipin_in = {wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_13499, wire_13498, wire_13489, wire_13488, wire_13479, wire_13478, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294, wire_10259, wire_10258, wire_10249, wire_10248, wire_10239, wire_10238, wire_13139, wire_13138, wire_13129, wire_13128, wire_13119, wire_13118, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_13493, wire_13492, wire_13483, wire_13482, wire_13473, wire_13472, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_10319, wire_10318, wire_10309, wire_10308, wire_10299, wire_10298, wire_10253, wire_10252, wire_10243, wire_10242, wire_10233, wire_10232, wire_13133, wire_13132, wire_13123, wire_13122, wire_13113, wire_13112, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_13497, wire_13496, wire_13487, wire_13486, wire_13477, wire_13476, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_10287, wire_10286, wire_10277, wire_10276, wire_10267, wire_10266, wire_10223, wire_10222, wire_10213, wire_10212, wire_10203, wire_10202, wire_13137, wire_13136, wire_13127, wire_13126, wire_13117, wire_13116, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_13491, wire_13490, wire_13481, wire_13480, wire_13471, wire_13470, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260, wire_10227, wire_10226, wire_10217, wire_10216, wire_10207, wire_10206, wire_13107, wire_13106, wire_13097, wire_13096, wire_13087, wire_13086, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_13527, wire_13526, wire_13517, wire_13516, wire_13507, wire_13506, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200, wire_13101, wire_13100, wire_13091, wire_13090, wire_13081, wire_13080, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_13521, wire_13520, wire_13511, wire_13510, wire_13501, wire_13500, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234};
    // IPIN TOTAL: 276
    assign lut_tile_1_8_ipin_in = {wire_6415, wire_6414, wire_6405, wire_6404, wire_6395, wire_6394, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_13649, wire_13648, wire_13629, wire_13628, wire_13609, wire_13608, wire_13589, wire_13588, wire_13569, wire_13568, wire_13549, wire_13548, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_13259, wire_13258, wire_13239, wire_13238, wire_13219, wire_13218, wire_13199, wire_13198, wire_13179, wire_13178, wire_13159, wire_13158, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_13645, wire_13644, wire_13625, wire_13624, wire_13605, wire_13604, wire_13585, wire_13584, wire_13565, wire_13564, wire_13545, wire_13544, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_13255, wire_13254, wire_13235, wire_13234, wire_13215, wire_13214, wire_13195, wire_13194, wire_13175, wire_13174, wire_13155, wire_13154, wire_6443, wire_6442, wire_6433, wire_6432, wire_6423, wire_6422, wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_13641, wire_13640, wire_13621, wire_13620, wire_13601, wire_13600, wire_13581, wire_13580, wire_13561, wire_13560, wire_13541, wire_13540, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_13251, wire_13250, wire_13231, wire_13230, wire_13211, wire_13210, wire_13191, wire_13190, wire_13171, wire_13170, wire_13151, wire_13150, wire_6447, wire_6446, wire_6437, wire_6436, wire_6427, wire_6426, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_13637, wire_13636, wire_13617, wire_13616, wire_13597, wire_13596, wire_13577, wire_13576, wire_13557, wire_13556, wire_13537, wire_13536, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_13249, wire_13248, wire_13221, wire_13220, wire_13209, wire_13208, wire_13181, wire_13180, wire_13169, wire_13168, wire_13141, wire_13140, wire_6441, wire_6440, wire_6431, wire_6430, wire_6421, wire_6420, wire_6387, wire_6386, wire_6377, wire_6376, wire_6367, wire_6366, wire_13635, wire_13634, wire_13615, wire_13614, wire_13595, wire_13594, wire_13575, wire_13574, wire_13555, wire_13554, wire_13535, wire_13534, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_13237, wire_13236, wire_13225, wire_13224, wire_13197, wire_13196, wire_13185, wire_13184, wire_13157, wire_13156, wire_13145, wire_13144, wire_6445, wire_6444, wire_6435, wire_6434, wire_6425, wire_6424, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360, wire_13631, wire_13630, wire_13611, wire_13610, wire_13591, wire_13590, wire_13571, wire_13570, wire_13551, wire_13550, wire_13531, wire_13530, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754};
    // IPIN TOTAL: 276
    assign lut_tile_2_8_ipin_in = {wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_13647, wire_13646, wire_13627, wire_13626, wire_13607, wire_13606, wire_13587, wire_13586, wire_13567, wire_13566, wire_13547, wire_13546, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13257, wire_13256, wire_13217, wire_13216, wire_13177, wire_13176, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_13643, wire_13642, wire_13623, wire_13622, wire_13603, wire_13602, wire_13583, wire_13582, wire_13563, wire_13562, wire_13543, wire_13542, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13233, wire_13232, wire_13193, wire_13192, wire_13153, wire_13152, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_13639, wire_13638, wire_13619, wire_13618, wire_13599, wire_13598, wire_13579, wire_13578, wire_13559, wire_13558, wire_13539, wire_13538, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13249, wire_13248, wire_13209, wire_13208, wire_13169, wire_13168, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_13635, wire_13634, wire_13615, wire_13614, wire_13595, wire_13594, wire_13575, wire_13574, wire_13555, wire_13554, wire_13535, wire_13534, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_13247, wire_13246, wire_13227, wire_13226, wire_13207, wire_13206, wire_13187, wire_13186, wire_13167, wire_13166, wire_13147, wire_13146, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13641, wire_13640, wire_13601, wire_13600, wire_13561, wire_13560, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_13243, wire_13242, wire_13223, wire_13222, wire_13203, wire_13202, wire_13183, wire_13182, wire_13163, wire_13162, wire_13143, wire_13142, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13617, wire_13616, wire_13577, wire_13576, wire_13537, wire_13536, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140};
    // IPIN TOTAL: 276
    assign lut_tile_3_8_ipin_in = {wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13633, wire_13632, wire_13593, wire_13592, wire_13553, wire_13552, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13243, wire_13242, wire_13203, wire_13202, wire_13163, wire_13162, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13649, wire_13648, wire_13609, wire_13608, wire_13569, wire_13568, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13259, wire_13258, wire_13219, wire_13218, wire_13179, wire_13178, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13625, wire_13624, wire_13585, wire_13584, wire_13545, wire_13544, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13235, wire_13234, wire_13195, wire_13194, wire_13155, wire_13154, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13641, wire_13640, wire_13601, wire_13600, wire_13561, wire_13560, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13241, wire_13240, wire_13201, wire_13200, wire_13161, wire_13160, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13627, wire_13626, wire_13587, wire_13586, wire_13547, wire_13546, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534};
    // IPIN TOTAL: 276
    assign lut_tile_4_8_ipin_in = {wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13643, wire_13642, wire_13603, wire_13602, wire_13563, wire_13562, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13619, wire_13618, wire_13579, wire_13578, wire_13539, wire_13538, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13635, wire_13634, wire_13595, wire_13594, wire_13555, wire_13554, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13227, wire_13226, wire_13187, wire_13186, wire_13147, wire_13146, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920};
    // IPIN TOTAL: 276
    assign lut_tile_5_8_ipin_in = {wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314};
    // IPIN TOTAL: 276
    assign lut_tile_6_8_ipin_in = {wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700};
    // IPIN TOTAL: 276
    assign lut_tile_7_8_ipin_in = {wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094};
    // IPIN TOTAL: 276
    assign lut_tile_8_8_ipin_in = {wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480};
    // IPIN TOTAL: 276
    assign lut_tile_9_8_ipin_in = {wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_13499, wire_13498, wire_13489, wire_13488, wire_13479, wire_13478, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_13493, wire_13492, wire_13483, wire_13482, wire_13473, wire_13472, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_13497, wire_13496, wire_13487, wire_13486, wire_13477, wire_13476, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_13887, wire_13886, wire_13877, wire_13876, wire_13867, wire_13866, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_13881, wire_13880, wire_13871, wire_13870, wire_13861, wire_13860, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874};
    // IPIN TOTAL: 276
    assign lut_tile_10_8_ipin_in = {wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_13885, wire_13884, wire_13875, wire_13874, wire_13865, wire_13864, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_10349, wire_10348, wire_10339, wire_10338, wire_10329, wire_10328, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_13525, wire_13524, wire_13515, wire_13514, wire_13505, wire_13504, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_13889, wire_13888, wire_13879, wire_13878, wire_13869, wire_13868, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_10343, wire_10342, wire_10333, wire_10332, wire_10323, wire_10322, wire_10289, wire_10288, wire_10279, wire_10278, wire_10269, wire_10268, wire_13529, wire_13528, wire_13519, wire_13518, wire_13509, wire_13508, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_13883, wire_13882, wire_13873, wire_13872, wire_13863, wire_13862, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_10313, wire_10312, wire_10303, wire_10302, wire_10293, wire_10292, wire_10257, wire_10256, wire_10247, wire_10246, wire_10237, wire_10236, wire_13523, wire_13522, wire_13513, wire_13512, wire_13503, wire_13502, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_13887, wire_13886, wire_13877, wire_13876, wire_13867, wire_13866, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_10317, wire_10316, wire_10307, wire_10306, wire_10297, wire_10296, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_13491, wire_13490, wire_13481, wire_13480, wire_13471, wire_13470, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_13911, wire_13910, wire_13901, wire_13900, wire_13891, wire_13890, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234, wire_13495, wire_13494, wire_13485, wire_13484, wire_13475, wire_13474, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_13915, wire_13914, wire_13905, wire_13904, wire_13895, wire_13894, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260};
    // IPIN TOTAL: 276
    assign lut_tile_1_9_ipin_in = {wire_6449, wire_6448, wire_6439, wire_6438, wire_6429, wire_6428, wire_6385, wire_6384, wire_6375, wire_6374, wire_6365, wire_6364, wire_14037, wire_14036, wire_14017, wire_14016, wire_13997, wire_13996, wire_13977, wire_13976, wire_13957, wire_13956, wire_13937, wire_13936, wire_6869, wire_6868, wire_6859, wire_6858, wire_6849, wire_6848, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_13647, wire_13646, wire_13627, wire_13626, wire_13607, wire_13606, wire_13587, wire_13586, wire_13567, wire_13566, wire_13547, wire_13546, wire_6443, wire_6442, wire_6433, wire_6432, wire_6423, wire_6422, wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_14033, wire_14032, wire_14013, wire_14012, wire_13993, wire_13992, wire_13973, wire_13972, wire_13953, wire_13952, wire_13933, wire_13932, wire_6863, wire_6862, wire_6853, wire_6852, wire_6843, wire_6842, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_13643, wire_13642, wire_13623, wire_13622, wire_13603, wire_13602, wire_13583, wire_13582, wire_13563, wire_13562, wire_13543, wire_13542, wire_6479, wire_6478, wire_6469, wire_6468, wire_6459, wire_6458, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_14029, wire_14028, wire_14009, wire_14008, wire_13989, wire_13988, wire_13969, wire_13968, wire_13949, wire_13948, wire_13929, wire_13928, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_13639, wire_13638, wire_13619, wire_13618, wire_13599, wire_13598, wire_13579, wire_13578, wire_13559, wire_13558, wire_13539, wire_13538, wire_6473, wire_6472, wire_6463, wire_6462, wire_6453, wire_6452, wire_6417, wire_6416, wire_6407, wire_6406, wire_6397, wire_6396, wire_14025, wire_14024, wire_14005, wire_14004, wire_13985, wire_13984, wire_13965, wire_13964, wire_13945, wire_13944, wire_13925, wire_13924, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_13637, wire_13636, wire_13617, wire_13616, wire_13597, wire_13596, wire_13577, wire_13576, wire_13557, wire_13556, wire_13537, wire_13536, wire_6477, wire_6476, wire_6467, wire_6466, wire_6457, wire_6456, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_14031, wire_14030, wire_14003, wire_14002, wire_13991, wire_13990, wire_13963, wire_13962, wire_13951, wire_13950, wire_13923, wire_13922, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_13633, wire_13632, wire_13613, wire_13612, wire_13593, wire_13592, wire_13573, wire_13572, wire_13553, wire_13552, wire_13533, wire_13532, wire_6471, wire_6470, wire_6461, wire_6460, wire_6451, wire_6450, wire_6415, wire_6414, wire_6405, wire_6404, wire_6395, wire_6394, wire_14019, wire_14018, wire_14007, wire_14006, wire_13979, wire_13978, wire_13967, wire_13966, wire_13939, wire_13938, wire_13927, wire_13926, wire_6865, wire_6864, wire_6855, wire_6854, wire_6845, wire_6844, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780};
    // IPIN TOTAL: 276
    assign lut_tile_2_9_ipin_in = {wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_14035, wire_14034, wire_14023, wire_14022, wire_13995, wire_13994, wire_13983, wire_13982, wire_13955, wire_13954, wire_13943, wire_13942, wire_7255, wire_7254, wire_7245, wire_7244, wire_7235, wire_7234, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13633, wire_13632, wire_13593, wire_13592, wire_13553, wire_13552, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_14039, wire_14038, wire_14011, wire_14010, wire_13999, wire_13998, wire_13971, wire_13970, wire_13959, wire_13958, wire_13931, wire_13930, wire_7259, wire_7258, wire_7249, wire_7248, wire_7239, wire_7238, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13649, wire_13648, wire_13609, wire_13608, wire_13569, wire_13568, wire_6863, wire_6862, wire_6853, wire_6852, wire_6843, wire_6842, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_14027, wire_14026, wire_14015, wire_14014, wire_13987, wire_13986, wire_13975, wire_13974, wire_13947, wire_13946, wire_13935, wire_13934, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13625, wire_13624, wire_13585, wire_13584, wire_13545, wire_13544, wire_6867, wire_6866, wire_6857, wire_6856, wire_6847, wire_6846, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_14031, wire_14030, wire_14003, wire_14002, wire_13991, wire_13990, wire_13963, wire_13962, wire_13951, wire_13950, wire_13923, wire_13922, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_13635, wire_13634, wire_13615, wire_13614, wire_13595, wire_13594, wire_13575, wire_13574, wire_13555, wire_13554, wire_13535, wire_13534, wire_6861, wire_6860, wire_6851, wire_6850, wire_6841, wire_6840, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_13631, wire_13630, wire_13611, wire_13610, wire_13591, wire_13590, wire_13571, wire_13570, wire_13551, wire_13550, wire_13531, wire_13530, wire_6865, wire_6864, wire_6855, wire_6854, wire_6845, wire_6844, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_14017, wire_14016, wire_13977, wire_13976, wire_13937, wire_13936, wire_7251, wire_7250, wire_7241, wire_7240, wire_7231, wire_7230, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174};
    // IPIN TOTAL: 276
    assign lut_tile_3_9_ipin_in = {wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_14033, wire_14032, wire_13993, wire_13992, wire_13953, wire_13952, wire_7649, wire_7648, wire_7639, wire_7638, wire_7629, wire_7628, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13643, wire_13642, wire_13603, wire_13602, wire_13563, wire_13562, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14009, wire_14008, wire_13969, wire_13968, wire_13929, wire_13928, wire_7643, wire_7642, wire_7633, wire_7632, wire_7623, wire_7622, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13619, wire_13618, wire_13579, wire_13578, wire_13539, wire_13538, wire_7259, wire_7258, wire_7249, wire_7248, wire_7239, wire_7238, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_14025, wire_14024, wire_13985, wire_13984, wire_13945, wire_13944, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13635, wire_13634, wire_13595, wire_13594, wire_13555, wire_13554, wire_7253, wire_7252, wire_7243, wire_7242, wire_7233, wire_7232, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13641, wire_13640, wire_13601, wire_13600, wire_13561, wire_13560, wire_7257, wire_7256, wire_7247, wire_7246, wire_7237, wire_7236, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14027, wire_14026, wire_13987, wire_13986, wire_13947, wire_13946, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13617, wire_13616, wire_13577, wire_13576, wire_13537, wire_13536, wire_7251, wire_7250, wire_7241, wire_7240, wire_7231, wire_7230, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_7645, wire_7644, wire_7635, wire_7634, wire_7625, wire_7624, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560};
    // IPIN TOTAL: 276
    assign lut_tile_4_9_ipin_in = {wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14019, wire_14018, wire_13979, wire_13978, wire_13939, wire_13938, wire_8035, wire_8034, wire_8025, wire_8024, wire_8015, wire_8014, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_14035, wire_14034, wire_13995, wire_13994, wire_13955, wire_13954, wire_8039, wire_8038, wire_8029, wire_8028, wire_8019, wire_8018, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_7643, wire_7642, wire_7633, wire_7632, wire_7623, wire_7622, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14011, wire_14010, wire_13971, wire_13970, wire_13931, wire_13930, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_7647, wire_7646, wire_7637, wire_7636, wire_7627, wire_7626, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14027, wire_14026, wire_13987, wire_13986, wire_13947, wire_13946, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7641, wire_7640, wire_7631, wire_7630, wire_7621, wire_7620, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13627, wire_13626, wire_13587, wire_13586, wire_13547, wire_13546, wire_7645, wire_7644, wire_7635, wire_7634, wire_7625, wire_7624, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_8031, wire_8030, wire_8021, wire_8020, wire_8011, wire_8010, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954};
    // IPIN TOTAL: 276
    assign lut_tile_5_9_ipin_in = {wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_8429, wire_8428, wire_8419, wire_8418, wire_8409, wire_8408, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_8423, wire_8422, wire_8413, wire_8412, wire_8403, wire_8402, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_8039, wire_8038, wire_8029, wire_8028, wire_8019, wire_8018, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_8033, wire_8032, wire_8023, wire_8022, wire_8013, wire_8012, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_8037, wire_8036, wire_8027, wire_8026, wire_8017, wire_8016, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_8031, wire_8030, wire_8021, wire_8020, wire_8011, wire_8010, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_8425, wire_8424, wire_8415, wire_8414, wire_8405, wire_8404, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340};
    // IPIN TOTAL: 276
    assign lut_tile_6_9_ipin_in = {wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_8815, wire_8814, wire_8805, wire_8804, wire_8795, wire_8794, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_8819, wire_8818, wire_8809, wire_8808, wire_8799, wire_8798, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_8423, wire_8422, wire_8413, wire_8412, wire_8403, wire_8402, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_8427, wire_8426, wire_8417, wire_8416, wire_8407, wire_8406, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_8421, wire_8420, wire_8411, wire_8410, wire_8401, wire_8400, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_8425, wire_8424, wire_8415, wire_8414, wire_8405, wire_8404, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_8811, wire_8810, wire_8801, wire_8800, wire_8791, wire_8790, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734};
    // IPIN TOTAL: 276
    assign lut_tile_7_9_ipin_in = {wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_9209, wire_9208, wire_9199, wire_9198, wire_9189, wire_9188, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_9203, wire_9202, wire_9193, wire_9192, wire_9183, wire_9182, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_8819, wire_8818, wire_8809, wire_8808, wire_8799, wire_8798, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_8813, wire_8812, wire_8803, wire_8802, wire_8793, wire_8792, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_8817, wire_8816, wire_8807, wire_8806, wire_8797, wire_8796, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_8811, wire_8810, wire_8801, wire_8800, wire_8791, wire_8790, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_9205, wire_9204, wire_9195, wire_9194, wire_9185, wire_9184, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120};
    // IPIN TOTAL: 276
    assign lut_tile_8_9_ipin_in = {wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_9595, wire_9594, wire_9585, wire_9584, wire_9575, wire_9574, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_9599, wire_9598, wire_9589, wire_9588, wire_9579, wire_9578, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_9203, wire_9202, wire_9193, wire_9192, wire_9183, wire_9182, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_9207, wire_9206, wire_9197, wire_9196, wire_9187, wire_9186, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_9201, wire_9200, wire_9191, wire_9190, wire_9181, wire_9180, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_9205, wire_9204, wire_9195, wire_9194, wire_9185, wire_9184, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_9591, wire_9590, wire_9581, wire_9580, wire_9571, wire_9570, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514};
    // IPIN TOTAL: 276
    assign lut_tile_9_9_ipin_in = {wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_9989, wire_9988, wire_9979, wire_9978, wire_9969, wire_9968, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_13885, wire_13884, wire_13875, wire_13874, wire_13865, wire_13864, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_9983, wire_9982, wire_9973, wire_9972, wire_9963, wire_9962, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_13889, wire_13888, wire_13879, wire_13878, wire_13869, wire_13868, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_9599, wire_9598, wire_9589, wire_9588, wire_9579, wire_9578, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_13883, wire_13882, wire_13873, wire_13872, wire_13863, wire_13862, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_9593, wire_9592, wire_9583, wire_9582, wire_9573, wire_9572, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_9597, wire_9596, wire_9587, wire_9586, wire_9577, wire_9576, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_14271, wire_14270, wire_14261, wire_14260, wire_14251, wire_14250, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_9591, wire_9590, wire_9581, wire_9580, wire_9571, wire_9570, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_14275, wire_14274, wire_14265, wire_14264, wire_14255, wire_14254, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_9985, wire_9984, wire_9975, wire_9974, wire_9965, wire_9964, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900};
    // IPIN TOTAL: 276
    assign lut_tile_10_9_ipin_in = {wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_14279, wire_14278, wire_14269, wire_14268, wire_14259, wire_14258, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_10375, wire_10374, wire_10365, wire_10364, wire_10355, wire_10354, wire_10319, wire_10318, wire_10309, wire_10308, wire_10299, wire_10298, wire_13919, wire_13918, wire_13909, wire_13908, wire_13899, wire_13898, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_14273, wire_14272, wire_14263, wire_14262, wire_14253, wire_14252, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_10379, wire_10378, wire_10369, wire_10368, wire_10359, wire_10358, wire_10313, wire_10312, wire_10303, wire_10302, wire_10293, wire_10292, wire_13913, wire_13912, wire_13903, wire_13902, wire_13893, wire_13892, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_9983, wire_9982, wire_9973, wire_9972, wire_9963, wire_9962, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_14277, wire_14276, wire_14267, wire_14266, wire_14257, wire_14256, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_10347, wire_10346, wire_10337, wire_10336, wire_10327, wire_10326, wire_10283, wire_10282, wire_10273, wire_10272, wire_10263, wire_10262, wire_13917, wire_13916, wire_13907, wire_13906, wire_13897, wire_13896, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_9987, wire_9986, wire_9977, wire_9976, wire_9967, wire_9966, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_14271, wire_14270, wire_14261, wire_14260, wire_14251, wire_14250, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_10341, wire_10340, wire_10331, wire_10330, wire_10321, wire_10320, wire_10287, wire_10286, wire_10277, wire_10276, wire_10267, wire_10266, wire_13887, wire_13886, wire_13877, wire_13876, wire_13867, wire_13866, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_9981, wire_9980, wire_9971, wire_9970, wire_9961, wire_9960, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_14307, wire_14306, wire_14297, wire_14296, wire_14287, wire_14286, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260, wire_13881, wire_13880, wire_13871, wire_13870, wire_13861, wire_13860, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_9985, wire_9984, wire_9975, wire_9974, wire_9965, wire_9964, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_14301, wire_14300, wire_14291, wire_14290, wire_14281, wire_14280, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_10371, wire_10370, wire_10361, wire_10360, wire_10351, wire_10350, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294};
    // IPIN TOTAL: 276
    assign lut_tile_1_10_ipin_in = {wire_6475, wire_6474, wire_6465, wire_6464, wire_6455, wire_6454, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_14425, wire_14424, wire_14413, wire_14412, wire_14385, wire_14384, wire_14373, wire_14372, wire_14345, wire_14344, wire_14333, wire_14332, wire_6895, wire_6894, wire_6885, wire_6884, wire_6875, wire_6874, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_14035, wire_14034, wire_14023, wire_14022, wire_13995, wire_13994, wire_13983, wire_13982, wire_13955, wire_13954, wire_13943, wire_13942, wire_6479, wire_6478, wire_6469, wire_6468, wire_6459, wire_6458, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_14429, wire_14428, wire_14401, wire_14400, wire_14389, wire_14388, wire_14361, wire_14360, wire_14349, wire_14348, wire_14321, wire_14320, wire_6899, wire_6898, wire_6889, wire_6888, wire_6879, wire_6878, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_14039, wire_14038, wire_14011, wire_14010, wire_13999, wire_13998, wire_13971, wire_13970, wire_13959, wire_13958, wire_13931, wire_13930, wire_6503, wire_6502, wire_6493, wire_6492, wire_6483, wire_6482, wire_6449, wire_6448, wire_6439, wire_6438, wire_6429, wire_6428, wire_14417, wire_14416, wire_14405, wire_14404, wire_14377, wire_14376, wire_14365, wire_14364, wire_14337, wire_14336, wire_14325, wire_14324, wire_6867, wire_6866, wire_6857, wire_6856, wire_6847, wire_6846, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_14027, wire_14026, wire_14015, wire_14014, wire_13987, wire_13986, wire_13975, wire_13974, wire_13947, wire_13946, wire_13935, wire_13934, wire_6507, wire_6506, wire_6497, wire_6496, wire_6487, wire_6486, wire_6443, wire_6442, wire_6433, wire_6432, wire_6423, wire_6422, wire_14421, wire_14420, wire_14393, wire_14392, wire_14381, wire_14380, wire_14353, wire_14352, wire_14341, wire_14340, wire_14313, wire_14312, wire_6861, wire_6860, wire_6851, wire_6850, wire_6841, wire_6840, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_14025, wire_14024, wire_14005, wire_14004, wire_13985, wire_13984, wire_13965, wire_13964, wire_13945, wire_13944, wire_13925, wire_13924, wire_6501, wire_6500, wire_6491, wire_6490, wire_6481, wire_6480, wire_6447, wire_6446, wire_6437, wire_6436, wire_6427, wire_6426, wire_14419, wire_14418, wire_14391, wire_14390, wire_14379, wire_14378, wire_14351, wire_14350, wire_14339, wire_14338, wire_14311, wire_14310, wire_6865, wire_6864, wire_6855, wire_6854, wire_6845, wire_6844, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_14021, wire_14020, wire_14001, wire_14000, wire_13981, wire_13980, wire_13961, wire_13960, wire_13941, wire_13940, wire_13921, wire_13920, wire_6505, wire_6504, wire_6495, wire_6494, wire_6485, wire_6484, wire_6441, wire_6440, wire_6431, wire_6430, wire_6421, wire_6420, wire_14407, wire_14406, wire_14395, wire_14394, wire_14367, wire_14366, wire_14355, wire_14354, wire_14327, wire_14326, wire_14315, wire_14314, wire_6891, wire_6890, wire_6881, wire_6880, wire_6871, wire_6870, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814};
    // IPIN TOTAL: 276
    assign lut_tile_2_10_ipin_in = {wire_6869, wire_6868, wire_6859, wire_6858, wire_6849, wire_6848, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_14423, wire_14422, wire_14411, wire_14410, wire_14383, wire_14382, wire_14371, wire_14370, wire_14343, wire_14342, wire_14331, wire_14330, wire_7289, wire_7288, wire_7279, wire_7278, wire_7269, wire_7268, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_14033, wire_14032, wire_13993, wire_13992, wire_13953, wire_13952, wire_6863, wire_6862, wire_6853, wire_6852, wire_6843, wire_6842, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_14427, wire_14426, wire_14399, wire_14398, wire_14387, wire_14386, wire_14359, wire_14358, wire_14347, wire_14346, wire_14319, wire_14318, wire_7283, wire_7282, wire_7273, wire_7272, wire_7263, wire_7262, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14009, wire_14008, wire_13969, wire_13968, wire_13929, wire_13928, wire_6899, wire_6898, wire_6889, wire_6888, wire_6879, wire_6878, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_14415, wire_14414, wire_14403, wire_14402, wire_14375, wire_14374, wire_14363, wire_14362, wire_14335, wire_14334, wire_14323, wire_14322, wire_7253, wire_7252, wire_7243, wire_7242, wire_7233, wire_7232, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_14025, wire_14024, wire_13985, wire_13984, wire_13945, wire_13944, wire_6893, wire_6892, wire_6883, wire_6882, wire_6873, wire_6872, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_14419, wire_14418, wire_14391, wire_14390, wire_14379, wire_14378, wire_14351, wire_14350, wire_14339, wire_14338, wire_14311, wire_14310, wire_7257, wire_7256, wire_7247, wire_7246, wire_7237, wire_7236, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_14031, wire_14030, wire_14003, wire_14002, wire_13991, wire_13990, wire_13963, wire_13962, wire_13951, wire_13950, wire_13923, wire_13922, wire_6897, wire_6896, wire_6887, wire_6886, wire_6877, wire_6876, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430, wire_14417, wire_14416, wire_14377, wire_14376, wire_14337, wire_14336, wire_7251, wire_7250, wire_7241, wire_7240, wire_7231, wire_7230, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_14019, wire_14018, wire_14007, wire_14006, wire_13979, wire_13978, wire_13967, wire_13966, wire_13939, wire_13938, wire_13927, wire_13926, wire_6891, wire_6890, wire_6881, wire_6880, wire_6871, wire_6870, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_14455, wire_14454, wire_14445, wire_14444, wire_14435, wire_14434, wire_14393, wire_14392, wire_14353, wire_14352, wire_14313, wire_14312, wire_7285, wire_7284, wire_7275, wire_7274, wire_7265, wire_7264, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200};
    // IPIN TOTAL: 276
    assign lut_tile_3_10_ipin_in = {wire_7255, wire_7254, wire_7245, wire_7244, wire_7235, wire_7234, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_14459, wire_14458, wire_14449, wire_14448, wire_14439, wire_14438, wire_14409, wire_14408, wire_14369, wire_14368, wire_14329, wire_14328, wire_7675, wire_7674, wire_7665, wire_7664, wire_7655, wire_7654, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14019, wire_14018, wire_13979, wire_13978, wire_13939, wire_13938, wire_7259, wire_7258, wire_7249, wire_7248, wire_7239, wire_7238, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_14453, wire_14452, wire_14443, wire_14442, wire_14433, wire_14432, wire_14425, wire_14424, wire_14385, wire_14384, wire_14345, wire_14344, wire_7679, wire_7678, wire_7669, wire_7668, wire_7659, wire_7658, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_14035, wire_14034, wire_13995, wire_13994, wire_13955, wire_13954, wire_7283, wire_7282, wire_7273, wire_7272, wire_7263, wire_7262, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_14401, wire_14400, wire_14361, wire_14360, wire_14321, wire_14320, wire_7647, wire_7646, wire_7637, wire_7636, wire_7627, wire_7626, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14011, wire_14010, wire_13971, wire_13970, wire_13931, wire_13930, wire_7287, wire_7286, wire_7277, wire_7276, wire_7267, wire_7266, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430, wire_14417, wire_14416, wire_14377, wire_14376, wire_14337, wire_14336, wire_7641, wire_7640, wire_7631, wire_7630, wire_7621, wire_7620, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_7281, wire_7280, wire_7271, wire_7270, wire_7261, wire_7260, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14395, wire_14394, wire_14355, wire_14354, wire_14315, wire_14314, wire_7645, wire_7644, wire_7635, wire_7634, wire_7625, wire_7624, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_14017, wire_14016, wire_13977, wire_13976, wire_13937, wire_13936, wire_7285, wire_7284, wire_7275, wire_7274, wire_7265, wire_7264, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_14411, wire_14410, wire_14371, wire_14370, wire_14331, wire_14330, wire_7671, wire_7670, wire_7661, wire_7660, wire_7651, wire_7650, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594};
    // IPIN TOTAL: 276
    assign lut_tile_4_10_ipin_in = {wire_7649, wire_7648, wire_7639, wire_7638, wire_7629, wire_7628, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_14485, wire_14484, wire_14475, wire_14474, wire_14465, wire_14464, wire_14427, wire_14426, wire_14387, wire_14386, wire_14347, wire_14346, wire_8069, wire_8068, wire_8059, wire_8058, wire_8049, wire_8048, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_7643, wire_7642, wire_7633, wire_7632, wire_7623, wire_7622, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_14489, wire_14488, wire_14479, wire_14478, wire_14469, wire_14468, wire_14403, wire_14402, wire_14363, wire_14362, wire_14323, wire_14322, wire_8063, wire_8062, wire_8053, wire_8052, wire_8043, wire_8042, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_7679, wire_7678, wire_7669, wire_7668, wire_7659, wire_7658, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_14483, wire_14482, wire_14473, wire_14472, wire_14463, wire_14462, wire_14419, wire_14418, wire_14379, wire_14378, wire_14339, wire_14338, wire_8033, wire_8032, wire_8023, wire_8022, wire_8013, wire_8012, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_7673, wire_7672, wire_7663, wire_7662, wire_7653, wire_7652, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14395, wire_14394, wire_14355, wire_14354, wire_14315, wire_14314, wire_8037, wire_8036, wire_8027, wire_8026, wire_8017, wire_8016, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14027, wire_14026, wire_13987, wire_13986, wire_13947, wire_13946, wire_7677, wire_7676, wire_7667, wire_7666, wire_7657, wire_7656, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_8031, wire_8030, wire_8021, wire_8020, wire_8011, wire_8010, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_7671, wire_7670, wire_7661, wire_7660, wire_7651, wire_7650, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_14515, wire_14514, wire_14505, wire_14504, wire_14495, wire_14494, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430, wire_8065, wire_8064, wire_8055, wire_8054, wire_8045, wire_8044, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980};
    // IPIN TOTAL: 276
    assign lut_tile_5_10_ipin_in = {wire_8035, wire_8034, wire_8025, wire_8024, wire_8015, wire_8014, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_14519, wire_14518, wire_14509, wire_14508, wire_14499, wire_14498, wire_14455, wire_14454, wire_14445, wire_14444, wire_14435, wire_14434, wire_8455, wire_8454, wire_8445, wire_8444, wire_8435, wire_8434, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_8039, wire_8038, wire_8029, wire_8028, wire_8019, wire_8018, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_14513, wire_14512, wire_14503, wire_14502, wire_14493, wire_14492, wire_14459, wire_14458, wire_14449, wire_14448, wire_14439, wire_14438, wire_8459, wire_8458, wire_8449, wire_8448, wire_8439, wire_8438, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_8063, wire_8062, wire_8053, wire_8052, wire_8043, wire_8042, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_14453, wire_14452, wire_14443, wire_14442, wire_14433, wire_14432, wire_8427, wire_8426, wire_8417, wire_8416, wire_8407, wire_8406, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_8067, wire_8066, wire_8057, wire_8056, wire_8047, wire_8046, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_8421, wire_8420, wire_8411, wire_8410, wire_8401, wire_8400, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_8061, wire_8060, wire_8051, wire_8050, wire_8041, wire_8040, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_8425, wire_8424, wire_8415, wire_8414, wire_8405, wire_8404, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_8065, wire_8064, wire_8055, wire_8054, wire_8045, wire_8044, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_14485, wire_14484, wire_14475, wire_14474, wire_14465, wire_14464, wire_8451, wire_8450, wire_8441, wire_8440, wire_8431, wire_8430, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374};
    // IPIN TOTAL: 276
    assign lut_tile_6_10_ipin_in = {wire_8429, wire_8428, wire_8419, wire_8418, wire_8409, wire_8408, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_14545, wire_14544, wire_14535, wire_14534, wire_14525, wire_14524, wire_14489, wire_14488, wire_14479, wire_14478, wire_14469, wire_14468, wire_8849, wire_8848, wire_8839, wire_8838, wire_8829, wire_8828, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_8423, wire_8422, wire_8413, wire_8412, wire_8403, wire_8402, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_14549, wire_14548, wire_14539, wire_14538, wire_14529, wire_14528, wire_14483, wire_14482, wire_14473, wire_14472, wire_14463, wire_14462, wire_8843, wire_8842, wire_8833, wire_8832, wire_8823, wire_8822, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_8459, wire_8458, wire_8449, wire_8448, wire_8439, wire_8438, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_14543, wire_14542, wire_14533, wire_14532, wire_14523, wire_14522, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_8813, wire_8812, wire_8803, wire_8802, wire_8793, wire_8792, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_8453, wire_8452, wire_8443, wire_8442, wire_8433, wire_8432, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_8817, wire_8816, wire_8807, wire_8806, wire_8797, wire_8796, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_8457, wire_8456, wire_8447, wire_8446, wire_8437, wire_8436, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_8811, wire_8810, wire_8801, wire_8800, wire_8791, wire_8790, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_8451, wire_8450, wire_8441, wire_8440, wire_8431, wire_8430, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_14575, wire_14574, wire_14565, wire_14564, wire_14555, wire_14554, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490, wire_8845, wire_8844, wire_8835, wire_8834, wire_8825, wire_8824, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760};
    // IPIN TOTAL: 276
    assign lut_tile_7_10_ipin_in = {wire_8815, wire_8814, wire_8805, wire_8804, wire_8795, wire_8794, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_14579, wire_14578, wire_14569, wire_14568, wire_14559, wire_14558, wire_14515, wire_14514, wire_14505, wire_14504, wire_14495, wire_14494, wire_9235, wire_9234, wire_9225, wire_9224, wire_9215, wire_9214, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_8819, wire_8818, wire_8809, wire_8808, wire_8799, wire_8798, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_14573, wire_14572, wire_14563, wire_14562, wire_14553, wire_14552, wire_14519, wire_14518, wire_14509, wire_14508, wire_14499, wire_14498, wire_9239, wire_9238, wire_9229, wire_9228, wire_9219, wire_9218, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_8843, wire_8842, wire_8833, wire_8832, wire_8823, wire_8822, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_14513, wire_14512, wire_14503, wire_14502, wire_14493, wire_14492, wire_9207, wire_9206, wire_9197, wire_9196, wire_9187, wire_9186, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_8847, wire_8846, wire_8837, wire_8836, wire_8827, wire_8826, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_9201, wire_9200, wire_9191, wire_9190, wire_9181, wire_9180, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_8841, wire_8840, wire_8831, wire_8830, wire_8821, wire_8820, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_9205, wire_9204, wire_9195, wire_9194, wire_9185, wire_9184, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_8845, wire_8844, wire_8835, wire_8834, wire_8825, wire_8824, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_14545, wire_14544, wire_14535, wire_14534, wire_14525, wire_14524, wire_9231, wire_9230, wire_9221, wire_9220, wire_9211, wire_9210, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154};
    // IPIN TOTAL: 276
    assign lut_tile_8_10_ipin_in = {wire_9209, wire_9208, wire_9199, wire_9198, wire_9189, wire_9188, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_14605, wire_14604, wire_14595, wire_14594, wire_14585, wire_14584, wire_14549, wire_14548, wire_14539, wire_14538, wire_14529, wire_14528, wire_9629, wire_9628, wire_9619, wire_9618, wire_9609, wire_9608, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_9203, wire_9202, wire_9193, wire_9192, wire_9183, wire_9182, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_14609, wire_14608, wire_14599, wire_14598, wire_14589, wire_14588, wire_14543, wire_14542, wire_14533, wire_14532, wire_14523, wire_14522, wire_9623, wire_9622, wire_9613, wire_9612, wire_9603, wire_9602, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_9239, wire_9238, wire_9229, wire_9228, wire_9219, wire_9218, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_14603, wire_14602, wire_14593, wire_14592, wire_14583, wire_14582, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_9593, wire_9592, wire_9583, wire_9582, wire_9573, wire_9572, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_9233, wire_9232, wire_9223, wire_9222, wire_9213, wire_9212, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_9597, wire_9596, wire_9587, wire_9586, wire_9577, wire_9576, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_9237, wire_9236, wire_9227, wire_9226, wire_9217, wire_9216, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_9591, wire_9590, wire_9581, wire_9580, wire_9571, wire_9570, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_9231, wire_9230, wire_9221, wire_9220, wire_9211, wire_9210, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_14635, wire_14634, wire_14625, wire_14624, wire_14615, wire_14614, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550, wire_9625, wire_9624, wire_9615, wire_9614, wire_9605, wire_9604, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540};
    // IPIN TOTAL: 276
    assign lut_tile_9_10_ipin_in = {wire_9595, wire_9594, wire_9585, wire_9584, wire_9575, wire_9574, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_14639, wire_14638, wire_14629, wire_14628, wire_14619, wire_14618, wire_14575, wire_14574, wire_14565, wire_14564, wire_14555, wire_14554, wire_10015, wire_10014, wire_10005, wire_10004, wire_9995, wire_9994, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_14279, wire_14278, wire_14269, wire_14268, wire_14259, wire_14258, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_9599, wire_9598, wire_9589, wire_9588, wire_9579, wire_9578, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_14633, wire_14632, wire_14623, wire_14622, wire_14613, wire_14612, wire_14579, wire_14578, wire_14569, wire_14568, wire_14559, wire_14558, wire_10019, wire_10018, wire_10009, wire_10008, wire_9999, wire_9998, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_14273, wire_14272, wire_14263, wire_14262, wire_14253, wire_14252, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_9623, wire_9622, wire_9613, wire_9612, wire_9603, wire_9602, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_14637, wire_14636, wire_14627, wire_14626, wire_14617, wire_14616, wire_14573, wire_14572, wire_14563, wire_14562, wire_14553, wire_14552, wire_9987, wire_9986, wire_9977, wire_9976, wire_9967, wire_9966, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_14277, wire_14276, wire_14267, wire_14266, wire_14257, wire_14256, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_9627, wire_9626, wire_9617, wire_9616, wire_9607, wire_9606, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_9981, wire_9980, wire_9971, wire_9970, wire_9961, wire_9960, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_9621, wire_9620, wire_9611, wire_9610, wire_9601, wire_9600, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_14667, wire_14666, wire_14657, wire_14656, wire_14647, wire_14646, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_9985, wire_9984, wire_9975, wire_9974, wire_9965, wire_9964, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_9625, wire_9624, wire_9615, wire_9614, wire_9605, wire_9604, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_14661, wire_14660, wire_14651, wire_14650, wire_14641, wire_14640, wire_14605, wire_14604, wire_14595, wire_14594, wire_14585, wire_14584, wire_10011, wire_10010, wire_10001, wire_10000, wire_9991, wire_9990, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934};
    // IPIN TOTAL: 276
    assign lut_tile_10_10_ipin_in = {wire_9989, wire_9988, wire_9979, wire_9978, wire_9969, wire_9968, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_14665, wire_14664, wire_14655, wire_14654, wire_14645, wire_14644, wire_14609, wire_14608, wire_14599, wire_14598, wire_14589, wire_14588, wire_10409, wire_10408, wire_10399, wire_10398, wire_10389, wire_10388, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_14305, wire_14304, wire_14295, wire_14294, wire_14285, wire_14284, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_9983, wire_9982, wire_9973, wire_9972, wire_9963, wire_9962, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_14669, wire_14668, wire_14659, wire_14658, wire_14649, wire_14648, wire_14603, wire_14602, wire_14593, wire_14592, wire_14583, wire_14582, wire_10403, wire_10402, wire_10393, wire_10392, wire_10383, wire_10382, wire_10349, wire_10348, wire_10339, wire_10338, wire_10329, wire_10328, wire_14309, wire_14308, wire_14299, wire_14298, wire_14289, wire_14288, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_10019, wire_10018, wire_10009, wire_10008, wire_9999, wire_9998, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_14663, wire_14662, wire_14653, wire_14652, wire_14643, wire_14642, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_10373, wire_10372, wire_10363, wire_10362, wire_10353, wire_10352, wire_10317, wire_10316, wire_10307, wire_10306, wire_10297, wire_10296, wire_14303, wire_14302, wire_14293, wire_14292, wire_14283, wire_14282, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_10013, wire_10012, wire_10003, wire_10002, wire_9993, wire_9992, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_14667, wire_14666, wire_14657, wire_14656, wire_14647, wire_14646, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_10377, wire_10376, wire_10367, wire_10366, wire_10357, wire_10356, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_14271, wire_14270, wire_14261, wire_14260, wire_14251, wire_14250, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_10017, wire_10016, wire_10007, wire_10006, wire_9997, wire_9996, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_14691, wire_14690, wire_14681, wire_14680, wire_14671, wire_14670, wire_14637, wire_14636, wire_14627, wire_14626, wire_14617, wire_14616, wire_10371, wire_10370, wire_10361, wire_10360, wire_10351, wire_10350, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294, wire_14275, wire_14274, wire_14265, wire_14264, wire_14255, wire_14254, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_10011, wire_10010, wire_10001, wire_10000, wire_9991, wire_9990, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_14695, wire_14694, wire_14685, wire_14684, wire_14675, wire_14674, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610, wire_10405, wire_10404, wire_10395, wire_10394, wire_10385, wire_10384, wire_10341, wire_10340, wire_10331, wire_10330, wire_10321, wire_10320};
    // IPIN TOTAL: 276


    // FPGA TILE OPIN
    assign wire_561 = lut_tile_1_1_opin_out[0];
    assign wire_562 = lut_tile_1_1_opin_out[1];
    assign wire_563 = lut_tile_1_1_opin_out[2];
    assign wire_564 = lut_tile_1_1_opin_out[3];
    assign wire_565 = lut_tile_1_1_opin_out[4];
    assign wire_566 = lut_tile_1_1_opin_out[5];
    assign wire_567 = lut_tile_1_1_opin_out[6];
    assign wire_568 = lut_tile_1_1_opin_out[7];
    assign wire_1077 = lut_tile_1_2_opin_out[0];
    assign wire_1078 = lut_tile_1_2_opin_out[1];
    assign wire_1079 = lut_tile_1_2_opin_out[2];
    assign wire_1080 = lut_tile_1_2_opin_out[3];
    assign wire_1081 = lut_tile_1_2_opin_out[4];
    assign wire_1082 = lut_tile_1_2_opin_out[5];
    assign wire_1083 = lut_tile_1_2_opin_out[6];
    assign wire_1084 = lut_tile_1_2_opin_out[7];
    assign wire_1593 = lut_tile_1_3_opin_out[0];
    assign wire_1594 = lut_tile_1_3_opin_out[1];
    assign wire_1595 = lut_tile_1_3_opin_out[2];
    assign wire_1596 = lut_tile_1_3_opin_out[3];
    assign wire_1597 = lut_tile_1_3_opin_out[4];
    assign wire_1598 = lut_tile_1_3_opin_out[5];
    assign wire_1599 = lut_tile_1_3_opin_out[6];
    assign wire_1600 = lut_tile_1_3_opin_out[7];
    assign wire_2109 = lut_tile_1_4_opin_out[0];
    assign wire_2110 = lut_tile_1_4_opin_out[1];
    assign wire_2111 = lut_tile_1_4_opin_out[2];
    assign wire_2112 = lut_tile_1_4_opin_out[3];
    assign wire_2113 = lut_tile_1_4_opin_out[4];
    assign wire_2114 = lut_tile_1_4_opin_out[5];
    assign wire_2115 = lut_tile_1_4_opin_out[6];
    assign wire_2116 = lut_tile_1_4_opin_out[7];
    assign wire_2625 = lut_tile_1_5_opin_out[0];
    assign wire_2626 = lut_tile_1_5_opin_out[1];
    assign wire_2627 = lut_tile_1_5_opin_out[2];
    assign wire_2628 = lut_tile_1_5_opin_out[3];
    assign wire_2629 = lut_tile_1_5_opin_out[4];
    assign wire_2630 = lut_tile_1_5_opin_out[5];
    assign wire_2631 = lut_tile_1_5_opin_out[6];
    assign wire_2632 = lut_tile_1_5_opin_out[7];
    assign wire_3141 = lut_tile_1_6_opin_out[0];
    assign wire_3142 = lut_tile_1_6_opin_out[1];
    assign wire_3143 = lut_tile_1_6_opin_out[2];
    assign wire_3144 = lut_tile_1_6_opin_out[3];
    assign wire_3145 = lut_tile_1_6_opin_out[4];
    assign wire_3146 = lut_tile_1_6_opin_out[5];
    assign wire_3147 = lut_tile_1_6_opin_out[6];
    assign wire_3148 = lut_tile_1_6_opin_out[7];
    assign wire_3657 = lut_tile_1_7_opin_out[0];
    assign wire_3658 = lut_tile_1_7_opin_out[1];
    assign wire_3659 = lut_tile_1_7_opin_out[2];
    assign wire_3660 = lut_tile_1_7_opin_out[3];
    assign wire_3661 = lut_tile_1_7_opin_out[4];
    assign wire_3662 = lut_tile_1_7_opin_out[5];
    assign wire_3663 = lut_tile_1_7_opin_out[6];
    assign wire_3664 = lut_tile_1_7_opin_out[7];
    assign wire_4173 = lut_tile_1_8_opin_out[0];
    assign wire_4174 = lut_tile_1_8_opin_out[1];
    assign wire_4175 = lut_tile_1_8_opin_out[2];
    assign wire_4176 = lut_tile_1_8_opin_out[3];
    assign wire_4177 = lut_tile_1_8_opin_out[4];
    assign wire_4178 = lut_tile_1_8_opin_out[5];
    assign wire_4179 = lut_tile_1_8_opin_out[6];
    assign wire_4180 = lut_tile_1_8_opin_out[7];
    assign wire_4689 = lut_tile_1_9_opin_out[0];
    assign wire_4690 = lut_tile_1_9_opin_out[1];
    assign wire_4691 = lut_tile_1_9_opin_out[2];
    assign wire_4692 = lut_tile_1_9_opin_out[3];
    assign wire_4693 = lut_tile_1_9_opin_out[4];
    assign wire_4694 = lut_tile_1_9_opin_out[5];
    assign wire_4695 = lut_tile_1_9_opin_out[6];
    assign wire_4696 = lut_tile_1_9_opin_out[7];
    assign wire_5205 = lut_tile_1_10_opin_out[0];
    assign wire_5206 = lut_tile_1_10_opin_out[1];
    assign wire_5207 = lut_tile_1_10_opin_out[2];
    assign wire_5208 = lut_tile_1_10_opin_out[3];
    assign wire_5209 = lut_tile_1_10_opin_out[4];
    assign wire_5210 = lut_tile_1_10_opin_out[5];
    assign wire_5211 = lut_tile_1_10_opin_out[6];
    assign wire_5212 = lut_tile_1_10_opin_out[7];
    assign wire_603 = lut_tile_2_1_opin_out[0];
    assign wire_604 = lut_tile_2_1_opin_out[1];
    assign wire_605 = lut_tile_2_1_opin_out[2];
    assign wire_606 = lut_tile_2_1_opin_out[3];
    assign wire_607 = lut_tile_2_1_opin_out[4];
    assign wire_608 = lut_tile_2_1_opin_out[5];
    assign wire_609 = lut_tile_2_1_opin_out[6];
    assign wire_610 = lut_tile_2_1_opin_out[7];
    assign wire_1119 = lut_tile_2_2_opin_out[0];
    assign wire_1120 = lut_tile_2_2_opin_out[1];
    assign wire_1121 = lut_tile_2_2_opin_out[2];
    assign wire_1122 = lut_tile_2_2_opin_out[3];
    assign wire_1123 = lut_tile_2_2_opin_out[4];
    assign wire_1124 = lut_tile_2_2_opin_out[5];
    assign wire_1125 = lut_tile_2_2_opin_out[6];
    assign wire_1126 = lut_tile_2_2_opin_out[7];
    assign wire_1635 = lut_tile_2_3_opin_out[0];
    assign wire_1636 = lut_tile_2_3_opin_out[1];
    assign wire_1637 = lut_tile_2_3_opin_out[2];
    assign wire_1638 = lut_tile_2_3_opin_out[3];
    assign wire_1639 = lut_tile_2_3_opin_out[4];
    assign wire_1640 = lut_tile_2_3_opin_out[5];
    assign wire_1641 = lut_tile_2_3_opin_out[6];
    assign wire_1642 = lut_tile_2_3_opin_out[7];
    assign wire_2151 = lut_tile_2_4_opin_out[0];
    assign wire_2152 = lut_tile_2_4_opin_out[1];
    assign wire_2153 = lut_tile_2_4_opin_out[2];
    assign wire_2154 = lut_tile_2_4_opin_out[3];
    assign wire_2155 = lut_tile_2_4_opin_out[4];
    assign wire_2156 = lut_tile_2_4_opin_out[5];
    assign wire_2157 = lut_tile_2_4_opin_out[6];
    assign wire_2158 = lut_tile_2_4_opin_out[7];
    assign wire_2667 = lut_tile_2_5_opin_out[0];
    assign wire_2668 = lut_tile_2_5_opin_out[1];
    assign wire_2669 = lut_tile_2_5_opin_out[2];
    assign wire_2670 = lut_tile_2_5_opin_out[3];
    assign wire_2671 = lut_tile_2_5_opin_out[4];
    assign wire_2672 = lut_tile_2_5_opin_out[5];
    assign wire_2673 = lut_tile_2_5_opin_out[6];
    assign wire_2674 = lut_tile_2_5_opin_out[7];
    assign wire_3183 = lut_tile_2_6_opin_out[0];
    assign wire_3184 = lut_tile_2_6_opin_out[1];
    assign wire_3185 = lut_tile_2_6_opin_out[2];
    assign wire_3186 = lut_tile_2_6_opin_out[3];
    assign wire_3187 = lut_tile_2_6_opin_out[4];
    assign wire_3188 = lut_tile_2_6_opin_out[5];
    assign wire_3189 = lut_tile_2_6_opin_out[6];
    assign wire_3190 = lut_tile_2_6_opin_out[7];
    assign wire_3699 = lut_tile_2_7_opin_out[0];
    assign wire_3700 = lut_tile_2_7_opin_out[1];
    assign wire_3701 = lut_tile_2_7_opin_out[2];
    assign wire_3702 = lut_tile_2_7_opin_out[3];
    assign wire_3703 = lut_tile_2_7_opin_out[4];
    assign wire_3704 = lut_tile_2_7_opin_out[5];
    assign wire_3705 = lut_tile_2_7_opin_out[6];
    assign wire_3706 = lut_tile_2_7_opin_out[7];
    assign wire_4215 = lut_tile_2_8_opin_out[0];
    assign wire_4216 = lut_tile_2_8_opin_out[1];
    assign wire_4217 = lut_tile_2_8_opin_out[2];
    assign wire_4218 = lut_tile_2_8_opin_out[3];
    assign wire_4219 = lut_tile_2_8_opin_out[4];
    assign wire_4220 = lut_tile_2_8_opin_out[5];
    assign wire_4221 = lut_tile_2_8_opin_out[6];
    assign wire_4222 = lut_tile_2_8_opin_out[7];
    assign wire_4731 = lut_tile_2_9_opin_out[0];
    assign wire_4732 = lut_tile_2_9_opin_out[1];
    assign wire_4733 = lut_tile_2_9_opin_out[2];
    assign wire_4734 = lut_tile_2_9_opin_out[3];
    assign wire_4735 = lut_tile_2_9_opin_out[4];
    assign wire_4736 = lut_tile_2_9_opin_out[5];
    assign wire_4737 = lut_tile_2_9_opin_out[6];
    assign wire_4738 = lut_tile_2_9_opin_out[7];
    assign wire_5247 = lut_tile_2_10_opin_out[0];
    assign wire_5248 = lut_tile_2_10_opin_out[1];
    assign wire_5249 = lut_tile_2_10_opin_out[2];
    assign wire_5250 = lut_tile_2_10_opin_out[3];
    assign wire_5251 = lut_tile_2_10_opin_out[4];
    assign wire_5252 = lut_tile_2_10_opin_out[5];
    assign wire_5253 = lut_tile_2_10_opin_out[6];
    assign wire_5254 = lut_tile_2_10_opin_out[7];
    assign wire_645 = lut_tile_3_1_opin_out[0];
    assign wire_646 = lut_tile_3_1_opin_out[1];
    assign wire_647 = lut_tile_3_1_opin_out[2];
    assign wire_648 = lut_tile_3_1_opin_out[3];
    assign wire_649 = lut_tile_3_1_opin_out[4];
    assign wire_650 = lut_tile_3_1_opin_out[5];
    assign wire_651 = lut_tile_3_1_opin_out[6];
    assign wire_652 = lut_tile_3_1_opin_out[7];
    assign wire_1161 = lut_tile_3_2_opin_out[0];
    assign wire_1162 = lut_tile_3_2_opin_out[1];
    assign wire_1163 = lut_tile_3_2_opin_out[2];
    assign wire_1164 = lut_tile_3_2_opin_out[3];
    assign wire_1165 = lut_tile_3_2_opin_out[4];
    assign wire_1166 = lut_tile_3_2_opin_out[5];
    assign wire_1167 = lut_tile_3_2_opin_out[6];
    assign wire_1168 = lut_tile_3_2_opin_out[7];
    assign wire_1677 = lut_tile_3_3_opin_out[0];
    assign wire_1678 = lut_tile_3_3_opin_out[1];
    assign wire_1679 = lut_tile_3_3_opin_out[2];
    assign wire_1680 = lut_tile_3_3_opin_out[3];
    assign wire_1681 = lut_tile_3_3_opin_out[4];
    assign wire_1682 = lut_tile_3_3_opin_out[5];
    assign wire_1683 = lut_tile_3_3_opin_out[6];
    assign wire_1684 = lut_tile_3_3_opin_out[7];
    assign wire_2193 = lut_tile_3_4_opin_out[0];
    assign wire_2194 = lut_tile_3_4_opin_out[1];
    assign wire_2195 = lut_tile_3_4_opin_out[2];
    assign wire_2196 = lut_tile_3_4_opin_out[3];
    assign wire_2197 = lut_tile_3_4_opin_out[4];
    assign wire_2198 = lut_tile_3_4_opin_out[5];
    assign wire_2199 = lut_tile_3_4_opin_out[6];
    assign wire_2200 = lut_tile_3_4_opin_out[7];
    assign wire_2709 = lut_tile_3_5_opin_out[0];
    assign wire_2710 = lut_tile_3_5_opin_out[1];
    assign wire_2711 = lut_tile_3_5_opin_out[2];
    assign wire_2712 = lut_tile_3_5_opin_out[3];
    assign wire_2713 = lut_tile_3_5_opin_out[4];
    assign wire_2714 = lut_tile_3_5_opin_out[5];
    assign wire_2715 = lut_tile_3_5_opin_out[6];
    assign wire_2716 = lut_tile_3_5_opin_out[7];
    assign wire_3225 = lut_tile_3_6_opin_out[0];
    assign wire_3226 = lut_tile_3_6_opin_out[1];
    assign wire_3227 = lut_tile_3_6_opin_out[2];
    assign wire_3228 = lut_tile_3_6_opin_out[3];
    assign wire_3229 = lut_tile_3_6_opin_out[4];
    assign wire_3230 = lut_tile_3_6_opin_out[5];
    assign wire_3231 = lut_tile_3_6_opin_out[6];
    assign wire_3232 = lut_tile_3_6_opin_out[7];
    assign wire_3741 = lut_tile_3_7_opin_out[0];
    assign wire_3742 = lut_tile_3_7_opin_out[1];
    assign wire_3743 = lut_tile_3_7_opin_out[2];
    assign wire_3744 = lut_tile_3_7_opin_out[3];
    assign wire_3745 = lut_tile_3_7_opin_out[4];
    assign wire_3746 = lut_tile_3_7_opin_out[5];
    assign wire_3747 = lut_tile_3_7_opin_out[6];
    assign wire_3748 = lut_tile_3_7_opin_out[7];
    assign wire_4257 = lut_tile_3_8_opin_out[0];
    assign wire_4258 = lut_tile_3_8_opin_out[1];
    assign wire_4259 = lut_tile_3_8_opin_out[2];
    assign wire_4260 = lut_tile_3_8_opin_out[3];
    assign wire_4261 = lut_tile_3_8_opin_out[4];
    assign wire_4262 = lut_tile_3_8_opin_out[5];
    assign wire_4263 = lut_tile_3_8_opin_out[6];
    assign wire_4264 = lut_tile_3_8_opin_out[7];
    assign wire_4773 = lut_tile_3_9_opin_out[0];
    assign wire_4774 = lut_tile_3_9_opin_out[1];
    assign wire_4775 = lut_tile_3_9_opin_out[2];
    assign wire_4776 = lut_tile_3_9_opin_out[3];
    assign wire_4777 = lut_tile_3_9_opin_out[4];
    assign wire_4778 = lut_tile_3_9_opin_out[5];
    assign wire_4779 = lut_tile_3_9_opin_out[6];
    assign wire_4780 = lut_tile_3_9_opin_out[7];
    assign wire_5289 = lut_tile_3_10_opin_out[0];
    assign wire_5290 = lut_tile_3_10_opin_out[1];
    assign wire_5291 = lut_tile_3_10_opin_out[2];
    assign wire_5292 = lut_tile_3_10_opin_out[3];
    assign wire_5293 = lut_tile_3_10_opin_out[4];
    assign wire_5294 = lut_tile_3_10_opin_out[5];
    assign wire_5295 = lut_tile_3_10_opin_out[6];
    assign wire_5296 = lut_tile_3_10_opin_out[7];
    assign wire_687 = lut_tile_4_1_opin_out[0];
    assign wire_688 = lut_tile_4_1_opin_out[1];
    assign wire_689 = lut_tile_4_1_opin_out[2];
    assign wire_690 = lut_tile_4_1_opin_out[3];
    assign wire_691 = lut_tile_4_1_opin_out[4];
    assign wire_692 = lut_tile_4_1_opin_out[5];
    assign wire_693 = lut_tile_4_1_opin_out[6];
    assign wire_694 = lut_tile_4_1_opin_out[7];
    assign wire_1203 = lut_tile_4_2_opin_out[0];
    assign wire_1204 = lut_tile_4_2_opin_out[1];
    assign wire_1205 = lut_tile_4_2_opin_out[2];
    assign wire_1206 = lut_tile_4_2_opin_out[3];
    assign wire_1207 = lut_tile_4_2_opin_out[4];
    assign wire_1208 = lut_tile_4_2_opin_out[5];
    assign wire_1209 = lut_tile_4_2_opin_out[6];
    assign wire_1210 = lut_tile_4_2_opin_out[7];
    assign wire_1719 = lut_tile_4_3_opin_out[0];
    assign wire_1720 = lut_tile_4_3_opin_out[1];
    assign wire_1721 = lut_tile_4_3_opin_out[2];
    assign wire_1722 = lut_tile_4_3_opin_out[3];
    assign wire_1723 = lut_tile_4_3_opin_out[4];
    assign wire_1724 = lut_tile_4_3_opin_out[5];
    assign wire_1725 = lut_tile_4_3_opin_out[6];
    assign wire_1726 = lut_tile_4_3_opin_out[7];
    assign wire_2235 = lut_tile_4_4_opin_out[0];
    assign wire_2236 = lut_tile_4_4_opin_out[1];
    assign wire_2237 = lut_tile_4_4_opin_out[2];
    assign wire_2238 = lut_tile_4_4_opin_out[3];
    assign wire_2239 = lut_tile_4_4_opin_out[4];
    assign wire_2240 = lut_tile_4_4_opin_out[5];
    assign wire_2241 = lut_tile_4_4_opin_out[6];
    assign wire_2242 = lut_tile_4_4_opin_out[7];
    assign wire_2751 = lut_tile_4_5_opin_out[0];
    assign wire_2752 = lut_tile_4_5_opin_out[1];
    assign wire_2753 = lut_tile_4_5_opin_out[2];
    assign wire_2754 = lut_tile_4_5_opin_out[3];
    assign wire_2755 = lut_tile_4_5_opin_out[4];
    assign wire_2756 = lut_tile_4_5_opin_out[5];
    assign wire_2757 = lut_tile_4_5_opin_out[6];
    assign wire_2758 = lut_tile_4_5_opin_out[7];
    assign wire_3267 = lut_tile_4_6_opin_out[0];
    assign wire_3268 = lut_tile_4_6_opin_out[1];
    assign wire_3269 = lut_tile_4_6_opin_out[2];
    assign wire_3270 = lut_tile_4_6_opin_out[3];
    assign wire_3271 = lut_tile_4_6_opin_out[4];
    assign wire_3272 = lut_tile_4_6_opin_out[5];
    assign wire_3273 = lut_tile_4_6_opin_out[6];
    assign wire_3274 = lut_tile_4_6_opin_out[7];
    assign wire_3783 = lut_tile_4_7_opin_out[0];
    assign wire_3784 = lut_tile_4_7_opin_out[1];
    assign wire_3785 = lut_tile_4_7_opin_out[2];
    assign wire_3786 = lut_tile_4_7_opin_out[3];
    assign wire_3787 = lut_tile_4_7_opin_out[4];
    assign wire_3788 = lut_tile_4_7_opin_out[5];
    assign wire_3789 = lut_tile_4_7_opin_out[6];
    assign wire_3790 = lut_tile_4_7_opin_out[7];
    assign wire_4299 = lut_tile_4_8_opin_out[0];
    assign wire_4300 = lut_tile_4_8_opin_out[1];
    assign wire_4301 = lut_tile_4_8_opin_out[2];
    assign wire_4302 = lut_tile_4_8_opin_out[3];
    assign wire_4303 = lut_tile_4_8_opin_out[4];
    assign wire_4304 = lut_tile_4_8_opin_out[5];
    assign wire_4305 = lut_tile_4_8_opin_out[6];
    assign wire_4306 = lut_tile_4_8_opin_out[7];
    assign wire_4815 = lut_tile_4_9_opin_out[0];
    assign wire_4816 = lut_tile_4_9_opin_out[1];
    assign wire_4817 = lut_tile_4_9_opin_out[2];
    assign wire_4818 = lut_tile_4_9_opin_out[3];
    assign wire_4819 = lut_tile_4_9_opin_out[4];
    assign wire_4820 = lut_tile_4_9_opin_out[5];
    assign wire_4821 = lut_tile_4_9_opin_out[6];
    assign wire_4822 = lut_tile_4_9_opin_out[7];
    assign wire_5331 = lut_tile_4_10_opin_out[0];
    assign wire_5332 = lut_tile_4_10_opin_out[1];
    assign wire_5333 = lut_tile_4_10_opin_out[2];
    assign wire_5334 = lut_tile_4_10_opin_out[3];
    assign wire_5335 = lut_tile_4_10_opin_out[4];
    assign wire_5336 = lut_tile_4_10_opin_out[5];
    assign wire_5337 = lut_tile_4_10_opin_out[6];
    assign wire_5338 = lut_tile_4_10_opin_out[7];
    assign wire_729 = lut_tile_5_1_opin_out[0];
    assign wire_730 = lut_tile_5_1_opin_out[1];
    assign wire_731 = lut_tile_5_1_opin_out[2];
    assign wire_732 = lut_tile_5_1_opin_out[3];
    assign wire_733 = lut_tile_5_1_opin_out[4];
    assign wire_734 = lut_tile_5_1_opin_out[5];
    assign wire_735 = lut_tile_5_1_opin_out[6];
    assign wire_736 = lut_tile_5_1_opin_out[7];
    assign wire_1245 = lut_tile_5_2_opin_out[0];
    assign wire_1246 = lut_tile_5_2_opin_out[1];
    assign wire_1247 = lut_tile_5_2_opin_out[2];
    assign wire_1248 = lut_tile_5_2_opin_out[3];
    assign wire_1249 = lut_tile_5_2_opin_out[4];
    assign wire_1250 = lut_tile_5_2_opin_out[5];
    assign wire_1251 = lut_tile_5_2_opin_out[6];
    assign wire_1252 = lut_tile_5_2_opin_out[7];
    assign wire_1761 = lut_tile_5_3_opin_out[0];
    assign wire_1762 = lut_tile_5_3_opin_out[1];
    assign wire_1763 = lut_tile_5_3_opin_out[2];
    assign wire_1764 = lut_tile_5_3_opin_out[3];
    assign wire_1765 = lut_tile_5_3_opin_out[4];
    assign wire_1766 = lut_tile_5_3_opin_out[5];
    assign wire_1767 = lut_tile_5_3_opin_out[6];
    assign wire_1768 = lut_tile_5_3_opin_out[7];
    assign wire_2277 = lut_tile_5_4_opin_out[0];
    assign wire_2278 = lut_tile_5_4_opin_out[1];
    assign wire_2279 = lut_tile_5_4_opin_out[2];
    assign wire_2280 = lut_tile_5_4_opin_out[3];
    assign wire_2281 = lut_tile_5_4_opin_out[4];
    assign wire_2282 = lut_tile_5_4_opin_out[5];
    assign wire_2283 = lut_tile_5_4_opin_out[6];
    assign wire_2284 = lut_tile_5_4_opin_out[7];
    assign wire_2793 = lut_tile_5_5_opin_out[0];
    assign wire_2794 = lut_tile_5_5_opin_out[1];
    assign wire_2795 = lut_tile_5_5_opin_out[2];
    assign wire_2796 = lut_tile_5_5_opin_out[3];
    assign wire_2797 = lut_tile_5_5_opin_out[4];
    assign wire_2798 = lut_tile_5_5_opin_out[5];
    assign wire_2799 = lut_tile_5_5_opin_out[6];
    assign wire_2800 = lut_tile_5_5_opin_out[7];
    assign wire_3309 = lut_tile_5_6_opin_out[0];
    assign wire_3310 = lut_tile_5_6_opin_out[1];
    assign wire_3311 = lut_tile_5_6_opin_out[2];
    assign wire_3312 = lut_tile_5_6_opin_out[3];
    assign wire_3313 = lut_tile_5_6_opin_out[4];
    assign wire_3314 = lut_tile_5_6_opin_out[5];
    assign wire_3315 = lut_tile_5_6_opin_out[6];
    assign wire_3316 = lut_tile_5_6_opin_out[7];
    assign wire_3825 = lut_tile_5_7_opin_out[0];
    assign wire_3826 = lut_tile_5_7_opin_out[1];
    assign wire_3827 = lut_tile_5_7_opin_out[2];
    assign wire_3828 = lut_tile_5_7_opin_out[3];
    assign wire_3829 = lut_tile_5_7_opin_out[4];
    assign wire_3830 = lut_tile_5_7_opin_out[5];
    assign wire_3831 = lut_tile_5_7_opin_out[6];
    assign wire_3832 = lut_tile_5_7_opin_out[7];
    assign wire_4341 = lut_tile_5_8_opin_out[0];
    assign wire_4342 = lut_tile_5_8_opin_out[1];
    assign wire_4343 = lut_tile_5_8_opin_out[2];
    assign wire_4344 = lut_tile_5_8_opin_out[3];
    assign wire_4345 = lut_tile_5_8_opin_out[4];
    assign wire_4346 = lut_tile_5_8_opin_out[5];
    assign wire_4347 = lut_tile_5_8_opin_out[6];
    assign wire_4348 = lut_tile_5_8_opin_out[7];
    assign wire_4857 = lut_tile_5_9_opin_out[0];
    assign wire_4858 = lut_tile_5_9_opin_out[1];
    assign wire_4859 = lut_tile_5_9_opin_out[2];
    assign wire_4860 = lut_tile_5_9_opin_out[3];
    assign wire_4861 = lut_tile_5_9_opin_out[4];
    assign wire_4862 = lut_tile_5_9_opin_out[5];
    assign wire_4863 = lut_tile_5_9_opin_out[6];
    assign wire_4864 = lut_tile_5_9_opin_out[7];
    assign wire_5373 = lut_tile_5_10_opin_out[0];
    assign wire_5374 = lut_tile_5_10_opin_out[1];
    assign wire_5375 = lut_tile_5_10_opin_out[2];
    assign wire_5376 = lut_tile_5_10_opin_out[3];
    assign wire_5377 = lut_tile_5_10_opin_out[4];
    assign wire_5378 = lut_tile_5_10_opin_out[5];
    assign wire_5379 = lut_tile_5_10_opin_out[6];
    assign wire_5380 = lut_tile_5_10_opin_out[7];
    assign wire_771 = lut_tile_6_1_opin_out[0];
    assign wire_772 = lut_tile_6_1_opin_out[1];
    assign wire_773 = lut_tile_6_1_opin_out[2];
    assign wire_774 = lut_tile_6_1_opin_out[3];
    assign wire_775 = lut_tile_6_1_opin_out[4];
    assign wire_776 = lut_tile_6_1_opin_out[5];
    assign wire_777 = lut_tile_6_1_opin_out[6];
    assign wire_778 = lut_tile_6_1_opin_out[7];
    assign wire_1287 = lut_tile_6_2_opin_out[0];
    assign wire_1288 = lut_tile_6_2_opin_out[1];
    assign wire_1289 = lut_tile_6_2_opin_out[2];
    assign wire_1290 = lut_tile_6_2_opin_out[3];
    assign wire_1291 = lut_tile_6_2_opin_out[4];
    assign wire_1292 = lut_tile_6_2_opin_out[5];
    assign wire_1293 = lut_tile_6_2_opin_out[6];
    assign wire_1294 = lut_tile_6_2_opin_out[7];
    assign wire_1803 = lut_tile_6_3_opin_out[0];
    assign wire_1804 = lut_tile_6_3_opin_out[1];
    assign wire_1805 = lut_tile_6_3_opin_out[2];
    assign wire_1806 = lut_tile_6_3_opin_out[3];
    assign wire_1807 = lut_tile_6_3_opin_out[4];
    assign wire_1808 = lut_tile_6_3_opin_out[5];
    assign wire_1809 = lut_tile_6_3_opin_out[6];
    assign wire_1810 = lut_tile_6_3_opin_out[7];
    assign wire_2319 = lut_tile_6_4_opin_out[0];
    assign wire_2320 = lut_tile_6_4_opin_out[1];
    assign wire_2321 = lut_tile_6_4_opin_out[2];
    assign wire_2322 = lut_tile_6_4_opin_out[3];
    assign wire_2323 = lut_tile_6_4_opin_out[4];
    assign wire_2324 = lut_tile_6_4_opin_out[5];
    assign wire_2325 = lut_tile_6_4_opin_out[6];
    assign wire_2326 = lut_tile_6_4_opin_out[7];
    assign wire_2835 = lut_tile_6_5_opin_out[0];
    assign wire_2836 = lut_tile_6_5_opin_out[1];
    assign wire_2837 = lut_tile_6_5_opin_out[2];
    assign wire_2838 = lut_tile_6_5_opin_out[3];
    assign wire_2839 = lut_tile_6_5_opin_out[4];
    assign wire_2840 = lut_tile_6_5_opin_out[5];
    assign wire_2841 = lut_tile_6_5_opin_out[6];
    assign wire_2842 = lut_tile_6_5_opin_out[7];
    assign wire_3351 = lut_tile_6_6_opin_out[0];
    assign wire_3352 = lut_tile_6_6_opin_out[1];
    assign wire_3353 = lut_tile_6_6_opin_out[2];
    assign wire_3354 = lut_tile_6_6_opin_out[3];
    assign wire_3355 = lut_tile_6_6_opin_out[4];
    assign wire_3356 = lut_tile_6_6_opin_out[5];
    assign wire_3357 = lut_tile_6_6_opin_out[6];
    assign wire_3358 = lut_tile_6_6_opin_out[7];
    assign wire_3867 = lut_tile_6_7_opin_out[0];
    assign wire_3868 = lut_tile_6_7_opin_out[1];
    assign wire_3869 = lut_tile_6_7_opin_out[2];
    assign wire_3870 = lut_tile_6_7_opin_out[3];
    assign wire_3871 = lut_tile_6_7_opin_out[4];
    assign wire_3872 = lut_tile_6_7_opin_out[5];
    assign wire_3873 = lut_tile_6_7_opin_out[6];
    assign wire_3874 = lut_tile_6_7_opin_out[7];
    assign wire_4383 = lut_tile_6_8_opin_out[0];
    assign wire_4384 = lut_tile_6_8_opin_out[1];
    assign wire_4385 = lut_tile_6_8_opin_out[2];
    assign wire_4386 = lut_tile_6_8_opin_out[3];
    assign wire_4387 = lut_tile_6_8_opin_out[4];
    assign wire_4388 = lut_tile_6_8_opin_out[5];
    assign wire_4389 = lut_tile_6_8_opin_out[6];
    assign wire_4390 = lut_tile_6_8_opin_out[7];
    assign wire_4899 = lut_tile_6_9_opin_out[0];
    assign wire_4900 = lut_tile_6_9_opin_out[1];
    assign wire_4901 = lut_tile_6_9_opin_out[2];
    assign wire_4902 = lut_tile_6_9_opin_out[3];
    assign wire_4903 = lut_tile_6_9_opin_out[4];
    assign wire_4904 = lut_tile_6_9_opin_out[5];
    assign wire_4905 = lut_tile_6_9_opin_out[6];
    assign wire_4906 = lut_tile_6_9_opin_out[7];
    assign wire_5415 = lut_tile_6_10_opin_out[0];
    assign wire_5416 = lut_tile_6_10_opin_out[1];
    assign wire_5417 = lut_tile_6_10_opin_out[2];
    assign wire_5418 = lut_tile_6_10_opin_out[3];
    assign wire_5419 = lut_tile_6_10_opin_out[4];
    assign wire_5420 = lut_tile_6_10_opin_out[5];
    assign wire_5421 = lut_tile_6_10_opin_out[6];
    assign wire_5422 = lut_tile_6_10_opin_out[7];
    assign wire_813 = lut_tile_7_1_opin_out[0];
    assign wire_814 = lut_tile_7_1_opin_out[1];
    assign wire_815 = lut_tile_7_1_opin_out[2];
    assign wire_816 = lut_tile_7_1_opin_out[3];
    assign wire_817 = lut_tile_7_1_opin_out[4];
    assign wire_818 = lut_tile_7_1_opin_out[5];
    assign wire_819 = lut_tile_7_1_opin_out[6];
    assign wire_820 = lut_tile_7_1_opin_out[7];
    assign wire_1329 = lut_tile_7_2_opin_out[0];
    assign wire_1330 = lut_tile_7_2_opin_out[1];
    assign wire_1331 = lut_tile_7_2_opin_out[2];
    assign wire_1332 = lut_tile_7_2_opin_out[3];
    assign wire_1333 = lut_tile_7_2_opin_out[4];
    assign wire_1334 = lut_tile_7_2_opin_out[5];
    assign wire_1335 = lut_tile_7_2_opin_out[6];
    assign wire_1336 = lut_tile_7_2_opin_out[7];
    assign wire_1845 = lut_tile_7_3_opin_out[0];
    assign wire_1846 = lut_tile_7_3_opin_out[1];
    assign wire_1847 = lut_tile_7_3_opin_out[2];
    assign wire_1848 = lut_tile_7_3_opin_out[3];
    assign wire_1849 = lut_tile_7_3_opin_out[4];
    assign wire_1850 = lut_tile_7_3_opin_out[5];
    assign wire_1851 = lut_tile_7_3_opin_out[6];
    assign wire_1852 = lut_tile_7_3_opin_out[7];
    assign wire_2361 = lut_tile_7_4_opin_out[0];
    assign wire_2362 = lut_tile_7_4_opin_out[1];
    assign wire_2363 = lut_tile_7_4_opin_out[2];
    assign wire_2364 = lut_tile_7_4_opin_out[3];
    assign wire_2365 = lut_tile_7_4_opin_out[4];
    assign wire_2366 = lut_tile_7_4_opin_out[5];
    assign wire_2367 = lut_tile_7_4_opin_out[6];
    assign wire_2368 = lut_tile_7_4_opin_out[7];
    assign wire_2877 = lut_tile_7_5_opin_out[0];
    assign wire_2878 = lut_tile_7_5_opin_out[1];
    assign wire_2879 = lut_tile_7_5_opin_out[2];
    assign wire_2880 = lut_tile_7_5_opin_out[3];
    assign wire_2881 = lut_tile_7_5_opin_out[4];
    assign wire_2882 = lut_tile_7_5_opin_out[5];
    assign wire_2883 = lut_tile_7_5_opin_out[6];
    assign wire_2884 = lut_tile_7_5_opin_out[7];
    assign wire_3393 = lut_tile_7_6_opin_out[0];
    assign wire_3394 = lut_tile_7_6_opin_out[1];
    assign wire_3395 = lut_tile_7_6_opin_out[2];
    assign wire_3396 = lut_tile_7_6_opin_out[3];
    assign wire_3397 = lut_tile_7_6_opin_out[4];
    assign wire_3398 = lut_tile_7_6_opin_out[5];
    assign wire_3399 = lut_tile_7_6_opin_out[6];
    assign wire_3400 = lut_tile_7_6_opin_out[7];
    assign wire_3909 = lut_tile_7_7_opin_out[0];
    assign wire_3910 = lut_tile_7_7_opin_out[1];
    assign wire_3911 = lut_tile_7_7_opin_out[2];
    assign wire_3912 = lut_tile_7_7_opin_out[3];
    assign wire_3913 = lut_tile_7_7_opin_out[4];
    assign wire_3914 = lut_tile_7_7_opin_out[5];
    assign wire_3915 = lut_tile_7_7_opin_out[6];
    assign wire_3916 = lut_tile_7_7_opin_out[7];
    assign wire_4425 = lut_tile_7_8_opin_out[0];
    assign wire_4426 = lut_tile_7_8_opin_out[1];
    assign wire_4427 = lut_tile_7_8_opin_out[2];
    assign wire_4428 = lut_tile_7_8_opin_out[3];
    assign wire_4429 = lut_tile_7_8_opin_out[4];
    assign wire_4430 = lut_tile_7_8_opin_out[5];
    assign wire_4431 = lut_tile_7_8_opin_out[6];
    assign wire_4432 = lut_tile_7_8_opin_out[7];
    assign wire_4941 = lut_tile_7_9_opin_out[0];
    assign wire_4942 = lut_tile_7_9_opin_out[1];
    assign wire_4943 = lut_tile_7_9_opin_out[2];
    assign wire_4944 = lut_tile_7_9_opin_out[3];
    assign wire_4945 = lut_tile_7_9_opin_out[4];
    assign wire_4946 = lut_tile_7_9_opin_out[5];
    assign wire_4947 = lut_tile_7_9_opin_out[6];
    assign wire_4948 = lut_tile_7_9_opin_out[7];
    assign wire_5457 = lut_tile_7_10_opin_out[0];
    assign wire_5458 = lut_tile_7_10_opin_out[1];
    assign wire_5459 = lut_tile_7_10_opin_out[2];
    assign wire_5460 = lut_tile_7_10_opin_out[3];
    assign wire_5461 = lut_tile_7_10_opin_out[4];
    assign wire_5462 = lut_tile_7_10_opin_out[5];
    assign wire_5463 = lut_tile_7_10_opin_out[6];
    assign wire_5464 = lut_tile_7_10_opin_out[7];
    assign wire_855 = lut_tile_8_1_opin_out[0];
    assign wire_856 = lut_tile_8_1_opin_out[1];
    assign wire_857 = lut_tile_8_1_opin_out[2];
    assign wire_858 = lut_tile_8_1_opin_out[3];
    assign wire_859 = lut_tile_8_1_opin_out[4];
    assign wire_860 = lut_tile_8_1_opin_out[5];
    assign wire_861 = lut_tile_8_1_opin_out[6];
    assign wire_862 = lut_tile_8_1_opin_out[7];
    assign wire_1371 = lut_tile_8_2_opin_out[0];
    assign wire_1372 = lut_tile_8_2_opin_out[1];
    assign wire_1373 = lut_tile_8_2_opin_out[2];
    assign wire_1374 = lut_tile_8_2_opin_out[3];
    assign wire_1375 = lut_tile_8_2_opin_out[4];
    assign wire_1376 = lut_tile_8_2_opin_out[5];
    assign wire_1377 = lut_tile_8_2_opin_out[6];
    assign wire_1378 = lut_tile_8_2_opin_out[7];
    assign wire_1887 = lut_tile_8_3_opin_out[0];
    assign wire_1888 = lut_tile_8_3_opin_out[1];
    assign wire_1889 = lut_tile_8_3_opin_out[2];
    assign wire_1890 = lut_tile_8_3_opin_out[3];
    assign wire_1891 = lut_tile_8_3_opin_out[4];
    assign wire_1892 = lut_tile_8_3_opin_out[5];
    assign wire_1893 = lut_tile_8_3_opin_out[6];
    assign wire_1894 = lut_tile_8_3_opin_out[7];
    assign wire_2403 = lut_tile_8_4_opin_out[0];
    assign wire_2404 = lut_tile_8_4_opin_out[1];
    assign wire_2405 = lut_tile_8_4_opin_out[2];
    assign wire_2406 = lut_tile_8_4_opin_out[3];
    assign wire_2407 = lut_tile_8_4_opin_out[4];
    assign wire_2408 = lut_tile_8_4_opin_out[5];
    assign wire_2409 = lut_tile_8_4_opin_out[6];
    assign wire_2410 = lut_tile_8_4_opin_out[7];
    assign wire_2919 = lut_tile_8_5_opin_out[0];
    assign wire_2920 = lut_tile_8_5_opin_out[1];
    assign wire_2921 = lut_tile_8_5_opin_out[2];
    assign wire_2922 = lut_tile_8_5_opin_out[3];
    assign wire_2923 = lut_tile_8_5_opin_out[4];
    assign wire_2924 = lut_tile_8_5_opin_out[5];
    assign wire_2925 = lut_tile_8_5_opin_out[6];
    assign wire_2926 = lut_tile_8_5_opin_out[7];
    assign wire_3435 = lut_tile_8_6_opin_out[0];
    assign wire_3436 = lut_tile_8_6_opin_out[1];
    assign wire_3437 = lut_tile_8_6_opin_out[2];
    assign wire_3438 = lut_tile_8_6_opin_out[3];
    assign wire_3439 = lut_tile_8_6_opin_out[4];
    assign wire_3440 = lut_tile_8_6_opin_out[5];
    assign wire_3441 = lut_tile_8_6_opin_out[6];
    assign wire_3442 = lut_tile_8_6_opin_out[7];
    assign wire_3951 = lut_tile_8_7_opin_out[0];
    assign wire_3952 = lut_tile_8_7_opin_out[1];
    assign wire_3953 = lut_tile_8_7_opin_out[2];
    assign wire_3954 = lut_tile_8_7_opin_out[3];
    assign wire_3955 = lut_tile_8_7_opin_out[4];
    assign wire_3956 = lut_tile_8_7_opin_out[5];
    assign wire_3957 = lut_tile_8_7_opin_out[6];
    assign wire_3958 = lut_tile_8_7_opin_out[7];
    assign wire_4467 = lut_tile_8_8_opin_out[0];
    assign wire_4468 = lut_tile_8_8_opin_out[1];
    assign wire_4469 = lut_tile_8_8_opin_out[2];
    assign wire_4470 = lut_tile_8_8_opin_out[3];
    assign wire_4471 = lut_tile_8_8_opin_out[4];
    assign wire_4472 = lut_tile_8_8_opin_out[5];
    assign wire_4473 = lut_tile_8_8_opin_out[6];
    assign wire_4474 = lut_tile_8_8_opin_out[7];
    assign wire_4983 = lut_tile_8_9_opin_out[0];
    assign wire_4984 = lut_tile_8_9_opin_out[1];
    assign wire_4985 = lut_tile_8_9_opin_out[2];
    assign wire_4986 = lut_tile_8_9_opin_out[3];
    assign wire_4987 = lut_tile_8_9_opin_out[4];
    assign wire_4988 = lut_tile_8_9_opin_out[5];
    assign wire_4989 = lut_tile_8_9_opin_out[6];
    assign wire_4990 = lut_tile_8_9_opin_out[7];
    assign wire_5499 = lut_tile_8_10_opin_out[0];
    assign wire_5500 = lut_tile_8_10_opin_out[1];
    assign wire_5501 = lut_tile_8_10_opin_out[2];
    assign wire_5502 = lut_tile_8_10_opin_out[3];
    assign wire_5503 = lut_tile_8_10_opin_out[4];
    assign wire_5504 = lut_tile_8_10_opin_out[5];
    assign wire_5505 = lut_tile_8_10_opin_out[6];
    assign wire_5506 = lut_tile_8_10_opin_out[7];
    assign wire_897 = lut_tile_9_1_opin_out[0];
    assign wire_898 = lut_tile_9_1_opin_out[1];
    assign wire_899 = lut_tile_9_1_opin_out[2];
    assign wire_900 = lut_tile_9_1_opin_out[3];
    assign wire_901 = lut_tile_9_1_opin_out[4];
    assign wire_902 = lut_tile_9_1_opin_out[5];
    assign wire_903 = lut_tile_9_1_opin_out[6];
    assign wire_904 = lut_tile_9_1_opin_out[7];
    assign wire_1413 = lut_tile_9_2_opin_out[0];
    assign wire_1414 = lut_tile_9_2_opin_out[1];
    assign wire_1415 = lut_tile_9_2_opin_out[2];
    assign wire_1416 = lut_tile_9_2_opin_out[3];
    assign wire_1417 = lut_tile_9_2_opin_out[4];
    assign wire_1418 = lut_tile_9_2_opin_out[5];
    assign wire_1419 = lut_tile_9_2_opin_out[6];
    assign wire_1420 = lut_tile_9_2_opin_out[7];
    assign wire_1929 = lut_tile_9_3_opin_out[0];
    assign wire_1930 = lut_tile_9_3_opin_out[1];
    assign wire_1931 = lut_tile_9_3_opin_out[2];
    assign wire_1932 = lut_tile_9_3_opin_out[3];
    assign wire_1933 = lut_tile_9_3_opin_out[4];
    assign wire_1934 = lut_tile_9_3_opin_out[5];
    assign wire_1935 = lut_tile_9_3_opin_out[6];
    assign wire_1936 = lut_tile_9_3_opin_out[7];
    assign wire_2445 = lut_tile_9_4_opin_out[0];
    assign wire_2446 = lut_tile_9_4_opin_out[1];
    assign wire_2447 = lut_tile_9_4_opin_out[2];
    assign wire_2448 = lut_tile_9_4_opin_out[3];
    assign wire_2449 = lut_tile_9_4_opin_out[4];
    assign wire_2450 = lut_tile_9_4_opin_out[5];
    assign wire_2451 = lut_tile_9_4_opin_out[6];
    assign wire_2452 = lut_tile_9_4_opin_out[7];
    assign wire_2961 = lut_tile_9_5_opin_out[0];
    assign wire_2962 = lut_tile_9_5_opin_out[1];
    assign wire_2963 = lut_tile_9_5_opin_out[2];
    assign wire_2964 = lut_tile_9_5_opin_out[3];
    assign wire_2965 = lut_tile_9_5_opin_out[4];
    assign wire_2966 = lut_tile_9_5_opin_out[5];
    assign wire_2967 = lut_tile_9_5_opin_out[6];
    assign wire_2968 = lut_tile_9_5_opin_out[7];
    assign wire_3477 = lut_tile_9_6_opin_out[0];
    assign wire_3478 = lut_tile_9_6_opin_out[1];
    assign wire_3479 = lut_tile_9_6_opin_out[2];
    assign wire_3480 = lut_tile_9_6_opin_out[3];
    assign wire_3481 = lut_tile_9_6_opin_out[4];
    assign wire_3482 = lut_tile_9_6_opin_out[5];
    assign wire_3483 = lut_tile_9_6_opin_out[6];
    assign wire_3484 = lut_tile_9_6_opin_out[7];
    assign wire_3993 = lut_tile_9_7_opin_out[0];
    assign wire_3994 = lut_tile_9_7_opin_out[1];
    assign wire_3995 = lut_tile_9_7_opin_out[2];
    assign wire_3996 = lut_tile_9_7_opin_out[3];
    assign wire_3997 = lut_tile_9_7_opin_out[4];
    assign wire_3998 = lut_tile_9_7_opin_out[5];
    assign wire_3999 = lut_tile_9_7_opin_out[6];
    assign wire_4000 = lut_tile_9_7_opin_out[7];
    assign wire_4509 = lut_tile_9_8_opin_out[0];
    assign wire_4510 = lut_tile_9_8_opin_out[1];
    assign wire_4511 = lut_tile_9_8_opin_out[2];
    assign wire_4512 = lut_tile_9_8_opin_out[3];
    assign wire_4513 = lut_tile_9_8_opin_out[4];
    assign wire_4514 = lut_tile_9_8_opin_out[5];
    assign wire_4515 = lut_tile_9_8_opin_out[6];
    assign wire_4516 = lut_tile_9_8_opin_out[7];
    assign wire_5025 = lut_tile_9_9_opin_out[0];
    assign wire_5026 = lut_tile_9_9_opin_out[1];
    assign wire_5027 = lut_tile_9_9_opin_out[2];
    assign wire_5028 = lut_tile_9_9_opin_out[3];
    assign wire_5029 = lut_tile_9_9_opin_out[4];
    assign wire_5030 = lut_tile_9_9_opin_out[5];
    assign wire_5031 = lut_tile_9_9_opin_out[6];
    assign wire_5032 = lut_tile_9_9_opin_out[7];
    assign wire_5541 = lut_tile_9_10_opin_out[0];
    assign wire_5542 = lut_tile_9_10_opin_out[1];
    assign wire_5543 = lut_tile_9_10_opin_out[2];
    assign wire_5544 = lut_tile_9_10_opin_out[3];
    assign wire_5545 = lut_tile_9_10_opin_out[4];
    assign wire_5546 = lut_tile_9_10_opin_out[5];
    assign wire_5547 = lut_tile_9_10_opin_out[6];
    assign wire_5548 = lut_tile_9_10_opin_out[7];
    assign wire_939 = lut_tile_10_1_opin_out[0];
    assign wire_940 = lut_tile_10_1_opin_out[1];
    assign wire_941 = lut_tile_10_1_opin_out[2];
    assign wire_942 = lut_tile_10_1_opin_out[3];
    assign wire_943 = lut_tile_10_1_opin_out[4];
    assign wire_944 = lut_tile_10_1_opin_out[5];
    assign wire_945 = lut_tile_10_1_opin_out[6];
    assign wire_946 = lut_tile_10_1_opin_out[7];
    assign wire_1455 = lut_tile_10_2_opin_out[0];
    assign wire_1456 = lut_tile_10_2_opin_out[1];
    assign wire_1457 = lut_tile_10_2_opin_out[2];
    assign wire_1458 = lut_tile_10_2_opin_out[3];
    assign wire_1459 = lut_tile_10_2_opin_out[4];
    assign wire_1460 = lut_tile_10_2_opin_out[5];
    assign wire_1461 = lut_tile_10_2_opin_out[6];
    assign wire_1462 = lut_tile_10_2_opin_out[7];
    assign wire_1971 = lut_tile_10_3_opin_out[0];
    assign wire_1972 = lut_tile_10_3_opin_out[1];
    assign wire_1973 = lut_tile_10_3_opin_out[2];
    assign wire_1974 = lut_tile_10_3_opin_out[3];
    assign wire_1975 = lut_tile_10_3_opin_out[4];
    assign wire_1976 = lut_tile_10_3_opin_out[5];
    assign wire_1977 = lut_tile_10_3_opin_out[6];
    assign wire_1978 = lut_tile_10_3_opin_out[7];
    assign wire_2487 = lut_tile_10_4_opin_out[0];
    assign wire_2488 = lut_tile_10_4_opin_out[1];
    assign wire_2489 = lut_tile_10_4_opin_out[2];
    assign wire_2490 = lut_tile_10_4_opin_out[3];
    assign wire_2491 = lut_tile_10_4_opin_out[4];
    assign wire_2492 = lut_tile_10_4_opin_out[5];
    assign wire_2493 = lut_tile_10_4_opin_out[6];
    assign wire_2494 = lut_tile_10_4_opin_out[7];
    assign wire_3003 = lut_tile_10_5_opin_out[0];
    assign wire_3004 = lut_tile_10_5_opin_out[1];
    assign wire_3005 = lut_tile_10_5_opin_out[2];
    assign wire_3006 = lut_tile_10_5_opin_out[3];
    assign wire_3007 = lut_tile_10_5_opin_out[4];
    assign wire_3008 = lut_tile_10_5_opin_out[5];
    assign wire_3009 = lut_tile_10_5_opin_out[6];
    assign wire_3010 = lut_tile_10_5_opin_out[7];
    assign wire_3519 = lut_tile_10_6_opin_out[0];
    assign wire_3520 = lut_tile_10_6_opin_out[1];
    assign wire_3521 = lut_tile_10_6_opin_out[2];
    assign wire_3522 = lut_tile_10_6_opin_out[3];
    assign wire_3523 = lut_tile_10_6_opin_out[4];
    assign wire_3524 = lut_tile_10_6_opin_out[5];
    assign wire_3525 = lut_tile_10_6_opin_out[6];
    assign wire_3526 = lut_tile_10_6_opin_out[7];
    assign wire_4035 = lut_tile_10_7_opin_out[0];
    assign wire_4036 = lut_tile_10_7_opin_out[1];
    assign wire_4037 = lut_tile_10_7_opin_out[2];
    assign wire_4038 = lut_tile_10_7_opin_out[3];
    assign wire_4039 = lut_tile_10_7_opin_out[4];
    assign wire_4040 = lut_tile_10_7_opin_out[5];
    assign wire_4041 = lut_tile_10_7_opin_out[6];
    assign wire_4042 = lut_tile_10_7_opin_out[7];
    assign wire_4551 = lut_tile_10_8_opin_out[0];
    assign wire_4552 = lut_tile_10_8_opin_out[1];
    assign wire_4553 = lut_tile_10_8_opin_out[2];
    assign wire_4554 = lut_tile_10_8_opin_out[3];
    assign wire_4555 = lut_tile_10_8_opin_out[4];
    assign wire_4556 = lut_tile_10_8_opin_out[5];
    assign wire_4557 = lut_tile_10_8_opin_out[6];
    assign wire_4558 = lut_tile_10_8_opin_out[7];
    assign wire_5067 = lut_tile_10_9_opin_out[0];
    assign wire_5068 = lut_tile_10_9_opin_out[1];
    assign wire_5069 = lut_tile_10_9_opin_out[2];
    assign wire_5070 = lut_tile_10_9_opin_out[3];
    assign wire_5071 = lut_tile_10_9_opin_out[4];
    assign wire_5072 = lut_tile_10_9_opin_out[5];
    assign wire_5073 = lut_tile_10_9_opin_out[6];
    assign wire_5074 = lut_tile_10_9_opin_out[7];
    assign wire_5583 = lut_tile_10_10_opin_out[0];
    assign wire_5584 = lut_tile_10_10_opin_out[1];
    assign wire_5585 = lut_tile_10_10_opin_out[2];
    assign wire_5586 = lut_tile_10_10_opin_out[3];
    assign wire_5587 = lut_tile_10_10_opin_out[4];
    assign wire_5588 = lut_tile_10_10_opin_out[5];
    assign wire_5589 = lut_tile_10_10_opin_out[6];
    assign wire_5590 = lut_tile_10_10_opin_out[7];
    // LUT TILE CHANXY 
    assign lut_tile_1_1_chanxy_in = {wire_6175, wire_6174, wire_10949, wire_6659, wire_6629, wire_6628, wire_6589, wire_6588, wire_6549, wire_6548, wire_6514, wire_1077, wire_6239, wire_6238, wire_6237, wire_6236, wire_6173, wire_6172, wire_6269, wire_6234, wire_10947, wire_6631, wire_6626, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_1077, wire_6233, wire_6232, wire_6253, wire_6170, wire_6231, wire_6230, wire_6229, wire_6228, wire_10945, wire_6633, wire_6623, wire_6622, wire_6618, wire_6583, wire_6582, wire_6543, wire_6542, wire_1077, wire_6169, wire_6168, wire_6267, wire_6226, wire_6225, wire_6224, wire_6223, wire_6222, wire_10943, wire_6635, wire_6621, wire_6620, wire_6610, wire_6581, wire_6580, wire_6541, wire_6540, wire_567, wire_6167, wire_6166, wire_6165, wire_6164, wire_6221, wire_6220, wire_6251, wire_6162, wire_10941, wire_6637, wire_6617, wire_6616, wire_6602, wire_6577, wire_6576, wire_6537, wire_6536, wire_567, wire_6161, wire_6160, wire_6265, wire_6218, wire_6159, wire_6158, wire_6157, wire_6156, wire_10939, wire_6639, wire_6615, wire_6614, wire_6594, wire_6575, wire_6574, wire_6535, wire_6534, wire_567, wire_6217, wire_6216, wire_6249, wire_6154, wire_6153, wire_6152, wire_6151, wire_6150, wire_10937, wire_6641, wire_6613, wire_6612, wire_6586, wire_6573, wire_6572, wire_6533, wire_6532, wire_1081, wire_567, wire_6215, wire_6214, wire_6213, wire_6212, wire_6149, wire_6148, wire_6263, wire_6210, wire_10935, wire_6643, wire_6609, wire_6608, wire_6578, wire_6569, wire_6568, wire_6529, wire_6528, wire_1081, wire_567, wire_6209, wire_6208, wire_6247, wire_6146, wire_6207, wire_6206, wire_6205, wire_6204, wire_10933, wire_6645, wire_6607, wire_6606, wire_6570, wire_6567, wire_6566, wire_6527, wire_6526, wire_1081, wire_567, wire_6145, wire_6144, wire_6261, wire_6202, wire_6201, wire_6200, wire_6199, wire_6198, wire_1081, wire_10931, wire_6647, wire_6605, wire_6604, wire_6565, wire_6564, wire_6562, wire_6525, wire_6524, wire_1081, wire_563, wire_6143, wire_6142, wire_1081, wire_6141, wire_6140, wire_1081, wire_6197, wire_6196, wire_1081, wire_6245, wire_6138, wire_1081, wire_10929, wire_6649, wire_6601, wire_6600, wire_6561, wire_6560, wire_6554, wire_6521, wire_6520, wire_1081, wire_563, wire_6137, wire_6136, wire_1081, wire_6259, wire_6194, wire_1077, wire_6135, wire_6134, wire_1077, wire_6133, wire_6132, wire_1077, wire_10927, wire_6651, wire_6599, wire_6598, wire_6559, wire_6558, wire_6546, wire_6519, wire_6518, wire_1081, wire_563, wire_6193, wire_6192, wire_1077, wire_6243, wire_6130, wire_1077, wire_6129, wire_6128, wire_1077, wire_6127, wire_6126, wire_567, wire_10925, wire_6653, wire_6597, wire_6596, wire_6557, wire_6556, wire_6538, wire_6517, wire_6516, wire_1077, wire_563, wire_6191, wire_6190, wire_567, wire_6189, wire_6188, wire_567, wire_6125, wire_6124, wire_567, wire_6257, wire_6186, wire_567, wire_10923, wire_6655, wire_6593, wire_6592, wire_6553, wire_6552, wire_6530, wire_6513, wire_6512, wire_1077, wire_563, wire_6185, wire_6184, wire_567, wire_6241, wire_6122, wire_563, wire_6183, wire_6182, wire_563, wire_6181, wire_6180, wire_563, wire_10921, wire_6657, wire_6591, wire_6590, wire_6551, wire_6550, wire_6522, wire_6511, wire_6510, wire_1077, wire_563, wire_6121, wire_6120, wire_563, wire_6255, wire_6178, wire_563, wire_6177, wire_6176, wire_563, wire_10465, wire_10464, wire_10923, wire_10919, wire_10918, wire_10908, wire_10879, wire_10878, wire_10839, wire_10838, wire_6659, wire_606, wire_10529, wire_10528, wire_10527, wire_10526, wire_10463, wire_10462, wire_10559, wire_10524, wire_10925, wire_10915, wire_10914, wire_10900, wire_10875, wire_10874, wire_10835, wire_10834, wire_6657, wire_606, wire_10523, wire_10522, wire_10543, wire_10460, wire_10521, wire_10520, wire_10519, wire_10518, wire_10927, wire_10913, wire_10912, wire_10892, wire_10873, wire_10872, wire_10833, wire_10832, wire_6655, wire_606, wire_10459, wire_10458, wire_10557, wire_10516, wire_10515, wire_10514, wire_10513, wire_10512, wire_10929, wire_10911, wire_10910, wire_10884, wire_10871, wire_10870, wire_10831, wire_10830, wire_6653, wire_566, wire_10457, wire_10456, wire_10455, wire_10454, wire_10511, wire_10510, wire_10541, wire_10452, wire_10931, wire_10907, wire_10906, wire_10876, wire_10867, wire_10866, wire_10827, wire_10826, wire_6651, wire_566, wire_10451, wire_10450, wire_10555, wire_10508, wire_10449, wire_10448, wire_10447, wire_10446, wire_10933, wire_10905, wire_10904, wire_10868, wire_10865, wire_10864, wire_10825, wire_10824, wire_6649, wire_566, wire_10507, wire_10506, wire_10539, wire_10444, wire_10443, wire_10442, wire_10441, wire_10440, wire_10935, wire_10903, wire_10902, wire_10863, wire_10862, wire_10860, wire_10823, wire_10822, wire_6647, wire_610, wire_566, wire_10505, wire_10504, wire_10503, wire_10502, wire_10439, wire_10438, wire_10553, wire_10500, wire_10937, wire_10899, wire_10898, wire_10859, wire_10858, wire_10852, wire_10819, wire_10818, wire_6645, wire_610, wire_566, wire_10499, wire_10498, wire_10537, wire_10436, wire_10497, wire_10496, wire_10495, wire_10494, wire_10939, wire_10897, wire_10896, wire_10857, wire_10856, wire_10844, wire_10817, wire_10816, wire_6643, wire_610, wire_566, wire_10435, wire_10434, wire_10551, wire_10492, wire_10491, wire_10490, wire_10489, wire_10488, wire_610, wire_10941, wire_10895, wire_10894, wire_10855, wire_10854, wire_10836, wire_10815, wire_10814, wire_6641, wire_610, wire_562, wire_10433, wire_10432, wire_610, wire_10431, wire_10430, wire_610, wire_10487, wire_10486, wire_610, wire_10535, wire_10428, wire_610, wire_10943, wire_10891, wire_10890, wire_10851, wire_10850, wire_10828, wire_10811, wire_10810, wire_6639, wire_610, wire_562, wire_10427, wire_10426, wire_610, wire_10549, wire_10484, wire_606, wire_10425, wire_10424, wire_606, wire_10423, wire_10422, wire_606, wire_10945, wire_10889, wire_10888, wire_10849, wire_10848, wire_10820, wire_10809, wire_10808, wire_6637, wire_610, wire_562, wire_10483, wire_10482, wire_606, wire_10533, wire_10420, wire_606, wire_10419, wire_10418, wire_606, wire_10417, wire_10416, wire_566, wire_10947, wire_10887, wire_10886, wire_10847, wire_10846, wire_10812, wire_10807, wire_10806, wire_6635, wire_606, wire_562, wire_10481, wire_10480, wire_566, wire_10479, wire_10478, wire_566, wire_10415, wire_10414, wire_566, wire_10547, wire_10476, wire_566, wire_10949, wire_10883, wire_10882, wire_10843, wire_10842, wire_10804, wire_10803, wire_10802, wire_6633, wire_606, wire_562, wire_10475, wire_10474, wire_566, wire_10531, wire_10412, wire_562, wire_10473, wire_10472, wire_562, wire_10471, wire_10470, wire_562, wire_10921, wire_10916, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_6631, wire_606, wire_562, wire_10411, wire_10410, wire_562, wire_10545, wire_10468, wire_562, wire_10467, wire_10466, wire_562};
    // CHNAXY TOTAL: 606
    assign wire_6510 = lut_tile_1_1_chanxy_out[0];
    assign wire_6512 = lut_tile_1_1_chanxy_out[1];
    assign wire_6514 = lut_tile_1_1_chanxy_out[2];
    assign wire_6515 = lut_tile_1_1_chanxy_out[3];
    assign wire_6516 = lut_tile_1_1_chanxy_out[4];
    assign wire_6518 = lut_tile_1_1_chanxy_out[5];
    assign wire_6520 = lut_tile_1_1_chanxy_out[6];
    assign wire_6522 = lut_tile_1_1_chanxy_out[7];
    assign wire_6523 = lut_tile_1_1_chanxy_out[8];
    assign wire_6524 = lut_tile_1_1_chanxy_out[9];
    assign wire_6526 = lut_tile_1_1_chanxy_out[10];
    assign wire_6528 = lut_tile_1_1_chanxy_out[11];
    assign wire_6530 = lut_tile_1_1_chanxy_out[12];
    assign wire_6531 = lut_tile_1_1_chanxy_out[13];
    assign wire_6532 = lut_tile_1_1_chanxy_out[14];
    assign wire_6534 = lut_tile_1_1_chanxy_out[15];
    assign wire_6536 = lut_tile_1_1_chanxy_out[16];
    assign wire_6538 = lut_tile_1_1_chanxy_out[17];
    assign wire_6539 = lut_tile_1_1_chanxy_out[18];
    assign wire_6540 = lut_tile_1_1_chanxy_out[19];
    assign wire_6542 = lut_tile_1_1_chanxy_out[20];
    assign wire_6544 = lut_tile_1_1_chanxy_out[21];
    assign wire_6546 = lut_tile_1_1_chanxy_out[22];
    assign wire_6547 = lut_tile_1_1_chanxy_out[23];
    assign wire_6548 = lut_tile_1_1_chanxy_out[24];
    assign wire_6550 = lut_tile_1_1_chanxy_out[25];
    assign wire_6552 = lut_tile_1_1_chanxy_out[26];
    assign wire_6554 = lut_tile_1_1_chanxy_out[27];
    assign wire_6555 = lut_tile_1_1_chanxy_out[28];
    assign wire_6556 = lut_tile_1_1_chanxy_out[29];
    assign wire_6558 = lut_tile_1_1_chanxy_out[30];
    assign wire_6560 = lut_tile_1_1_chanxy_out[31];
    assign wire_6562 = lut_tile_1_1_chanxy_out[32];
    assign wire_6563 = lut_tile_1_1_chanxy_out[33];
    assign wire_6564 = lut_tile_1_1_chanxy_out[34];
    assign wire_6566 = lut_tile_1_1_chanxy_out[35];
    assign wire_6568 = lut_tile_1_1_chanxy_out[36];
    assign wire_6570 = lut_tile_1_1_chanxy_out[37];
    assign wire_6571 = lut_tile_1_1_chanxy_out[38];
    assign wire_6572 = lut_tile_1_1_chanxy_out[39];
    assign wire_6574 = lut_tile_1_1_chanxy_out[40];
    assign wire_6576 = lut_tile_1_1_chanxy_out[41];
    assign wire_6578 = lut_tile_1_1_chanxy_out[42];
    assign wire_6579 = lut_tile_1_1_chanxy_out[43];
    assign wire_6580 = lut_tile_1_1_chanxy_out[44];
    assign wire_6582 = lut_tile_1_1_chanxy_out[45];
    assign wire_6584 = lut_tile_1_1_chanxy_out[46];
    assign wire_6586 = lut_tile_1_1_chanxy_out[47];
    assign wire_6587 = lut_tile_1_1_chanxy_out[48];
    assign wire_6588 = lut_tile_1_1_chanxy_out[49];
    assign wire_6590 = lut_tile_1_1_chanxy_out[50];
    assign wire_6592 = lut_tile_1_1_chanxy_out[51];
    assign wire_6594 = lut_tile_1_1_chanxy_out[52];
    assign wire_6595 = lut_tile_1_1_chanxy_out[53];
    assign wire_6596 = lut_tile_1_1_chanxy_out[54];
    assign wire_6598 = lut_tile_1_1_chanxy_out[55];
    assign wire_6600 = lut_tile_1_1_chanxy_out[56];
    assign wire_6602 = lut_tile_1_1_chanxy_out[57];
    assign wire_6603 = lut_tile_1_1_chanxy_out[58];
    assign wire_6604 = lut_tile_1_1_chanxy_out[59];
    assign wire_6606 = lut_tile_1_1_chanxy_out[60];
    assign wire_6608 = lut_tile_1_1_chanxy_out[61];
    assign wire_6610 = lut_tile_1_1_chanxy_out[62];
    assign wire_6611 = lut_tile_1_1_chanxy_out[63];
    assign wire_6612 = lut_tile_1_1_chanxy_out[64];
    assign wire_6614 = lut_tile_1_1_chanxy_out[65];
    assign wire_6616 = lut_tile_1_1_chanxy_out[66];
    assign wire_6618 = lut_tile_1_1_chanxy_out[67];
    assign wire_6619 = lut_tile_1_1_chanxy_out[68];
    assign wire_6620 = lut_tile_1_1_chanxy_out[69];
    assign wire_6622 = lut_tile_1_1_chanxy_out[70];
    assign wire_6624 = lut_tile_1_1_chanxy_out[71];
    assign wire_6626 = lut_tile_1_1_chanxy_out[72];
    assign wire_6627 = lut_tile_1_1_chanxy_out[73];
    assign wire_6628 = lut_tile_1_1_chanxy_out[74];
    assign wire_10800 = lut_tile_1_1_chanxy_out[75];
    assign wire_10802 = lut_tile_1_1_chanxy_out[76];
    assign wire_10804 = lut_tile_1_1_chanxy_out[77];
    assign wire_10805 = lut_tile_1_1_chanxy_out[78];
    assign wire_10806 = lut_tile_1_1_chanxy_out[79];
    assign wire_10808 = lut_tile_1_1_chanxy_out[80];
    assign wire_10810 = lut_tile_1_1_chanxy_out[81];
    assign wire_10812 = lut_tile_1_1_chanxy_out[82];
    assign wire_10813 = lut_tile_1_1_chanxy_out[83];
    assign wire_10814 = lut_tile_1_1_chanxy_out[84];
    assign wire_10816 = lut_tile_1_1_chanxy_out[85];
    assign wire_10818 = lut_tile_1_1_chanxy_out[86];
    assign wire_10820 = lut_tile_1_1_chanxy_out[87];
    assign wire_10821 = lut_tile_1_1_chanxy_out[88];
    assign wire_10822 = lut_tile_1_1_chanxy_out[89];
    assign wire_10824 = lut_tile_1_1_chanxy_out[90];
    assign wire_10826 = lut_tile_1_1_chanxy_out[91];
    assign wire_10828 = lut_tile_1_1_chanxy_out[92];
    assign wire_10829 = lut_tile_1_1_chanxy_out[93];
    assign wire_10830 = lut_tile_1_1_chanxy_out[94];
    assign wire_10832 = lut_tile_1_1_chanxy_out[95];
    assign wire_10834 = lut_tile_1_1_chanxy_out[96];
    assign wire_10836 = lut_tile_1_1_chanxy_out[97];
    assign wire_10837 = lut_tile_1_1_chanxy_out[98];
    assign wire_10838 = lut_tile_1_1_chanxy_out[99];
    assign wire_10840 = lut_tile_1_1_chanxy_out[100];
    assign wire_10842 = lut_tile_1_1_chanxy_out[101];
    assign wire_10844 = lut_tile_1_1_chanxy_out[102];
    assign wire_10845 = lut_tile_1_1_chanxy_out[103];
    assign wire_10846 = lut_tile_1_1_chanxy_out[104];
    assign wire_10848 = lut_tile_1_1_chanxy_out[105];
    assign wire_10850 = lut_tile_1_1_chanxy_out[106];
    assign wire_10852 = lut_tile_1_1_chanxy_out[107];
    assign wire_10853 = lut_tile_1_1_chanxy_out[108];
    assign wire_10854 = lut_tile_1_1_chanxy_out[109];
    assign wire_10856 = lut_tile_1_1_chanxy_out[110];
    assign wire_10858 = lut_tile_1_1_chanxy_out[111];
    assign wire_10860 = lut_tile_1_1_chanxy_out[112];
    assign wire_10861 = lut_tile_1_1_chanxy_out[113];
    assign wire_10862 = lut_tile_1_1_chanxy_out[114];
    assign wire_10864 = lut_tile_1_1_chanxy_out[115];
    assign wire_10866 = lut_tile_1_1_chanxy_out[116];
    assign wire_10868 = lut_tile_1_1_chanxy_out[117];
    assign wire_10869 = lut_tile_1_1_chanxy_out[118];
    assign wire_10870 = lut_tile_1_1_chanxy_out[119];
    assign wire_10872 = lut_tile_1_1_chanxy_out[120];
    assign wire_10874 = lut_tile_1_1_chanxy_out[121];
    assign wire_10876 = lut_tile_1_1_chanxy_out[122];
    assign wire_10877 = lut_tile_1_1_chanxy_out[123];
    assign wire_10878 = lut_tile_1_1_chanxy_out[124];
    assign wire_10880 = lut_tile_1_1_chanxy_out[125];
    assign wire_10882 = lut_tile_1_1_chanxy_out[126];
    assign wire_10884 = lut_tile_1_1_chanxy_out[127];
    assign wire_10885 = lut_tile_1_1_chanxy_out[128];
    assign wire_10886 = lut_tile_1_1_chanxy_out[129];
    assign wire_10888 = lut_tile_1_1_chanxy_out[130];
    assign wire_10890 = lut_tile_1_1_chanxy_out[131];
    assign wire_10892 = lut_tile_1_1_chanxy_out[132];
    assign wire_10893 = lut_tile_1_1_chanxy_out[133];
    assign wire_10894 = lut_tile_1_1_chanxy_out[134];
    assign wire_10896 = lut_tile_1_1_chanxy_out[135];
    assign wire_10898 = lut_tile_1_1_chanxy_out[136];
    assign wire_10900 = lut_tile_1_1_chanxy_out[137];
    assign wire_10901 = lut_tile_1_1_chanxy_out[138];
    assign wire_10902 = lut_tile_1_1_chanxy_out[139];
    assign wire_10904 = lut_tile_1_1_chanxy_out[140];
    assign wire_10906 = lut_tile_1_1_chanxy_out[141];
    assign wire_10908 = lut_tile_1_1_chanxy_out[142];
    assign wire_10909 = lut_tile_1_1_chanxy_out[143];
    assign wire_10910 = lut_tile_1_1_chanxy_out[144];
    assign wire_10912 = lut_tile_1_1_chanxy_out[145];
    assign wire_10914 = lut_tile_1_1_chanxy_out[146];
    assign wire_10916 = lut_tile_1_1_chanxy_out[147];
    assign wire_10917 = lut_tile_1_1_chanxy_out[148];
    assign wire_10918 = lut_tile_1_1_chanxy_out[149];
   // CHANXY OUT
    assign lut_tile_1_2_chanxy_in = {wire_11339, wire_6689, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6516, wire_1593, wire_6175, wire_6174, wire_6239, wire_6238, wire_6299, wire_6236, wire_6283, wire_6172, wire_11337, wire_6661, wire_6628, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_1593, wire_6269, wire_6268, wire_6233, wire_6232, wire_6253, wire_6252, wire_6231, wire_6230, wire_11335, wire_6663, wire_6623, wire_6622, wire_6620, wire_6583, wire_6582, wire_6543, wire_6542, wire_1593, wire_6297, wire_6228, wire_6169, wire_6168, wire_6267, wire_6266, wire_6225, wire_6224, wire_11333, wire_6665, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6612, wire_1083, wire_6223, wire_6222, wire_6167, wire_6166, wire_6281, wire_6164, wire_6295, wire_6220, wire_11331, wire_6667, wire_6617, wire_6616, wire_6604, wire_6577, wire_6576, wire_6537, wire_6536, wire_1083, wire_6251, wire_6250, wire_6161, wire_6160, wire_6265, wire_6264, wire_6159, wire_6158, wire_11329, wire_6669, wire_6615, wire_6614, wire_6596, wire_6575, wire_6574, wire_6535, wire_6534, wire_1083, wire_6279, wire_6156, wire_6217, wire_6216, wire_6249, wire_6248, wire_6153, wire_6152, wire_11327, wire_6671, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6588, wire_1597, wire_1083, wire_6151, wire_6150, wire_6215, wire_6214, wire_6293, wire_6212, wire_6277, wire_6148, wire_11325, wire_6673, wire_6609, wire_6608, wire_6580, wire_6569, wire_6568, wire_6529, wire_6528, wire_1597, wire_1083, wire_6263, wire_6262, wire_6209, wire_6208, wire_6247, wire_6246, wire_6207, wire_6206, wire_11323, wire_6675, wire_6607, wire_6606, wire_6572, wire_6567, wire_6566, wire_6527, wire_6526, wire_1597, wire_1083, wire_6291, wire_6204, wire_6145, wire_6144, wire_6261, wire_6260, wire_6201, wire_6200, wire_11321, wire_6677, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6564, wire_1597, wire_1079, wire_6199, wire_6198, wire_1597, wire_6143, wire_6142, wire_1597, wire_6275, wire_6140, wire_1597, wire_6289, wire_6196, wire_1597, wire_11319, wire_6679, wire_6601, wire_6600, wire_6561, wire_6560, wire_6556, wire_6521, wire_6520, wire_1597, wire_1079, wire_6245, wire_6244, wire_1597, wire_6137, wire_6136, wire_1597, wire_6259, wire_6258, wire_1593, wire_6135, wire_6134, wire_1593, wire_11317, wire_6681, wire_6599, wire_6598, wire_6559, wire_6558, wire_6548, wire_6519, wire_6518, wire_1597, wire_1079, wire_6273, wire_6132, wire_1593, wire_6193, wire_6192, wire_1593, wire_6243, wire_6242, wire_1593, wire_6129, wire_6128, wire_1593, wire_11315, wire_6683, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6540, wire_1593, wire_1079, wire_6127, wire_6126, wire_1083, wire_6191, wire_6190, wire_1083, wire_6287, wire_6188, wire_1083, wire_6271, wire_6124, wire_1083, wire_11313, wire_6685, wire_6593, wire_6592, wire_6553, wire_6552, wire_6532, wire_6513, wire_6512, wire_1593, wire_1079, wire_6257, wire_6256, wire_1083, wire_6185, wire_6184, wire_1083, wire_6241, wire_6240, wire_1079, wire_6183, wire_6182, wire_1079, wire_11311, wire_6687, wire_6591, wire_6590, wire_6551, wire_6550, wire_6524, wire_6511, wire_6510, wire_1593, wire_1079, wire_6285, wire_6180, wire_1079, wire_6121, wire_6120, wire_1079, wire_6255, wire_6254, wire_1079, wire_6177, wire_6176, wire_1079, wire_10947, wire_10919, wire_10918, wire_10916, wire_10879, wire_10878, wire_10839, wire_10838, wire_6626, wire_1122, wire_10945, wire_10915, wire_10914, wire_10875, wire_10874, wire_10835, wire_10834, wire_10804, wire_6618, wire_1122, wire_10943, wire_10913, wire_10912, wire_10873, wire_10872, wire_10833, wire_10832, wire_10812, wire_6610, wire_1122, wire_10941, wire_10911, wire_10910, wire_10871, wire_10870, wire_10831, wire_10830, wire_10820, wire_6602, wire_1082, wire_10939, wire_10907, wire_10906, wire_10867, wire_10866, wire_10828, wire_10827, wire_10826, wire_6594, wire_1082, wire_10937, wire_10905, wire_10904, wire_10865, wire_10864, wire_10836, wire_10825, wire_10824, wire_6586, wire_1082, wire_10935, wire_10903, wire_10902, wire_10863, wire_10862, wire_10844, wire_10823, wire_10822, wire_6578, wire_1126, wire_1082, wire_10933, wire_10899, wire_10898, wire_10859, wire_10858, wire_10852, wire_10819, wire_10818, wire_6570, wire_1126, wire_1082, wire_10931, wire_10897, wire_10896, wire_10860, wire_10857, wire_10856, wire_10817, wire_10816, wire_6562, wire_1126, wire_1082, wire_10929, wire_10895, wire_10894, wire_10868, wire_10855, wire_10854, wire_10815, wire_10814, wire_6554, wire_1126, wire_1078, wire_10927, wire_10891, wire_10890, wire_10876, wire_10851, wire_10850, wire_10811, wire_10810, wire_6546, wire_1126, wire_1078, wire_10925, wire_10889, wire_10888, wire_10884, wire_10849, wire_10848, wire_10809, wire_10808, wire_6538, wire_1126, wire_1078, wire_10923, wire_10892, wire_10887, wire_10886, wire_10847, wire_10846, wire_10807, wire_10806, wire_6530, wire_1122, wire_1078, wire_10921, wire_10900, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_6522, wire_1122, wire_1078, wire_10949, wire_10908, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_6514, wire_1122, wire_1078, wire_11313, wire_11307, wire_11306, wire_11300, wire_11267, wire_11266, wire_11227, wire_11226, wire_6689, wire_1122, wire_11315, wire_11305, wire_11304, wire_11292, wire_11265, wire_11264, wire_11225, wire_11224, wire_6687, wire_1122, wire_11317, wire_11303, wire_11302, wire_11284, wire_11263, wire_11262, wire_11223, wire_11222, wire_6685, wire_1122, wire_11319, wire_11299, wire_11298, wire_11276, wire_11259, wire_11258, wire_11219, wire_11218, wire_6683, wire_1082, wire_11321, wire_11297, wire_11296, wire_11268, wire_11257, wire_11256, wire_11217, wire_11216, wire_6681, wire_1082, wire_11323, wire_11295, wire_11294, wire_11260, wire_11255, wire_11254, wire_11215, wire_11214, wire_6679, wire_1082, wire_11325, wire_11291, wire_11290, wire_11252, wire_11251, wire_11250, wire_11211, wire_11210, wire_6677, wire_1126, wire_1082, wire_11327, wire_11289, wire_11288, wire_11249, wire_11248, wire_11244, wire_11209, wire_11208, wire_6675, wire_1126, wire_1082, wire_11329, wire_11287, wire_11286, wire_11247, wire_11246, wire_11236, wire_11207, wire_11206, wire_6673, wire_1126, wire_1082, wire_11331, wire_11283, wire_11282, wire_11243, wire_11242, wire_11228, wire_11203, wire_11202, wire_6671, wire_1126, wire_1078, wire_11333, wire_11281, wire_11280, wire_11241, wire_11240, wire_11220, wire_11201, wire_11200, wire_6669, wire_1126, wire_1078, wire_11335, wire_11279, wire_11278, wire_11239, wire_11238, wire_11212, wire_11199, wire_11198, wire_6667, wire_1126, wire_1078, wire_11337, wire_11275, wire_11274, wire_11235, wire_11234, wire_11204, wire_11195, wire_11194, wire_6665, wire_1122, wire_1078, wire_11339, wire_11273, wire_11272, wire_11233, wire_11232, wire_11196, wire_11193, wire_11192, wire_6663, wire_1122, wire_1078, wire_11311, wire_11308, wire_11271, wire_11270, wire_11231, wire_11230, wire_11191, wire_11190, wire_6661, wire_1122, wire_1078};
    // CHNAXY TOTAL: 621
    assign wire_6517 = lut_tile_1_2_chanxy_out[0];
    assign wire_6525 = lut_tile_1_2_chanxy_out[1];
    assign wire_6533 = lut_tile_1_2_chanxy_out[2];
    assign wire_6541 = lut_tile_1_2_chanxy_out[3];
    assign wire_6549 = lut_tile_1_2_chanxy_out[4];
    assign wire_6557 = lut_tile_1_2_chanxy_out[5];
    assign wire_6565 = lut_tile_1_2_chanxy_out[6];
    assign wire_6573 = lut_tile_1_2_chanxy_out[7];
    assign wire_6581 = lut_tile_1_2_chanxy_out[8];
    assign wire_6589 = lut_tile_1_2_chanxy_out[9];
    assign wire_6597 = lut_tile_1_2_chanxy_out[10];
    assign wire_6605 = lut_tile_1_2_chanxy_out[11];
    assign wire_6613 = lut_tile_1_2_chanxy_out[12];
    assign wire_6621 = lut_tile_1_2_chanxy_out[13];
    assign wire_6629 = lut_tile_1_2_chanxy_out[14];
    assign wire_6630 = lut_tile_1_2_chanxy_out[15];
    assign wire_6632 = lut_tile_1_2_chanxy_out[16];
    assign wire_6634 = lut_tile_1_2_chanxy_out[17];
    assign wire_6636 = lut_tile_1_2_chanxy_out[18];
    assign wire_6638 = lut_tile_1_2_chanxy_out[19];
    assign wire_6640 = lut_tile_1_2_chanxy_out[20];
    assign wire_6642 = lut_tile_1_2_chanxy_out[21];
    assign wire_6644 = lut_tile_1_2_chanxy_out[22];
    assign wire_6646 = lut_tile_1_2_chanxy_out[23];
    assign wire_6648 = lut_tile_1_2_chanxy_out[24];
    assign wire_6650 = lut_tile_1_2_chanxy_out[25];
    assign wire_6652 = lut_tile_1_2_chanxy_out[26];
    assign wire_6654 = lut_tile_1_2_chanxy_out[27];
    assign wire_6656 = lut_tile_1_2_chanxy_out[28];
    assign wire_6658 = lut_tile_1_2_chanxy_out[29];
    assign wire_11190 = lut_tile_1_2_chanxy_out[30];
    assign wire_11192 = lut_tile_1_2_chanxy_out[31];
    assign wire_11194 = lut_tile_1_2_chanxy_out[32];
    assign wire_11196 = lut_tile_1_2_chanxy_out[33];
    assign wire_11197 = lut_tile_1_2_chanxy_out[34];
    assign wire_11198 = lut_tile_1_2_chanxy_out[35];
    assign wire_11200 = lut_tile_1_2_chanxy_out[36];
    assign wire_11202 = lut_tile_1_2_chanxy_out[37];
    assign wire_11204 = lut_tile_1_2_chanxy_out[38];
    assign wire_11205 = lut_tile_1_2_chanxy_out[39];
    assign wire_11206 = lut_tile_1_2_chanxy_out[40];
    assign wire_11208 = lut_tile_1_2_chanxy_out[41];
    assign wire_11210 = lut_tile_1_2_chanxy_out[42];
    assign wire_11212 = lut_tile_1_2_chanxy_out[43];
    assign wire_11213 = lut_tile_1_2_chanxy_out[44];
    assign wire_11214 = lut_tile_1_2_chanxy_out[45];
    assign wire_11216 = lut_tile_1_2_chanxy_out[46];
    assign wire_11218 = lut_tile_1_2_chanxy_out[47];
    assign wire_11220 = lut_tile_1_2_chanxy_out[48];
    assign wire_11221 = lut_tile_1_2_chanxy_out[49];
    assign wire_11222 = lut_tile_1_2_chanxy_out[50];
    assign wire_11224 = lut_tile_1_2_chanxy_out[51];
    assign wire_11226 = lut_tile_1_2_chanxy_out[52];
    assign wire_11228 = lut_tile_1_2_chanxy_out[53];
    assign wire_11229 = lut_tile_1_2_chanxy_out[54];
    assign wire_11230 = lut_tile_1_2_chanxy_out[55];
    assign wire_11232 = lut_tile_1_2_chanxy_out[56];
    assign wire_11234 = lut_tile_1_2_chanxy_out[57];
    assign wire_11236 = lut_tile_1_2_chanxy_out[58];
    assign wire_11237 = lut_tile_1_2_chanxy_out[59];
    assign wire_11238 = lut_tile_1_2_chanxy_out[60];
    assign wire_11240 = lut_tile_1_2_chanxy_out[61];
    assign wire_11242 = lut_tile_1_2_chanxy_out[62];
    assign wire_11244 = lut_tile_1_2_chanxy_out[63];
    assign wire_11245 = lut_tile_1_2_chanxy_out[64];
    assign wire_11246 = lut_tile_1_2_chanxy_out[65];
    assign wire_11248 = lut_tile_1_2_chanxy_out[66];
    assign wire_11250 = lut_tile_1_2_chanxy_out[67];
    assign wire_11252 = lut_tile_1_2_chanxy_out[68];
    assign wire_11253 = lut_tile_1_2_chanxy_out[69];
    assign wire_11254 = lut_tile_1_2_chanxy_out[70];
    assign wire_11256 = lut_tile_1_2_chanxy_out[71];
    assign wire_11258 = lut_tile_1_2_chanxy_out[72];
    assign wire_11260 = lut_tile_1_2_chanxy_out[73];
    assign wire_11261 = lut_tile_1_2_chanxy_out[74];
    assign wire_11262 = lut_tile_1_2_chanxy_out[75];
    assign wire_11264 = lut_tile_1_2_chanxy_out[76];
    assign wire_11266 = lut_tile_1_2_chanxy_out[77];
    assign wire_11268 = lut_tile_1_2_chanxy_out[78];
    assign wire_11269 = lut_tile_1_2_chanxy_out[79];
    assign wire_11270 = lut_tile_1_2_chanxy_out[80];
    assign wire_11272 = lut_tile_1_2_chanxy_out[81];
    assign wire_11274 = lut_tile_1_2_chanxy_out[82];
    assign wire_11276 = lut_tile_1_2_chanxy_out[83];
    assign wire_11277 = lut_tile_1_2_chanxy_out[84];
    assign wire_11278 = lut_tile_1_2_chanxy_out[85];
    assign wire_11280 = lut_tile_1_2_chanxy_out[86];
    assign wire_11282 = lut_tile_1_2_chanxy_out[87];
    assign wire_11284 = lut_tile_1_2_chanxy_out[88];
    assign wire_11285 = lut_tile_1_2_chanxy_out[89];
    assign wire_11286 = lut_tile_1_2_chanxy_out[90];
    assign wire_11288 = lut_tile_1_2_chanxy_out[91];
    assign wire_11290 = lut_tile_1_2_chanxy_out[92];
    assign wire_11292 = lut_tile_1_2_chanxy_out[93];
    assign wire_11293 = lut_tile_1_2_chanxy_out[94];
    assign wire_11294 = lut_tile_1_2_chanxy_out[95];
    assign wire_11296 = lut_tile_1_2_chanxy_out[96];
    assign wire_11298 = lut_tile_1_2_chanxy_out[97];
    assign wire_11300 = lut_tile_1_2_chanxy_out[98];
    assign wire_11301 = lut_tile_1_2_chanxy_out[99];
    assign wire_11302 = lut_tile_1_2_chanxy_out[100];
    assign wire_11304 = lut_tile_1_2_chanxy_out[101];
    assign wire_11306 = lut_tile_1_2_chanxy_out[102];
    assign wire_11308 = lut_tile_1_2_chanxy_out[103];
    assign wire_11309 = lut_tile_1_2_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_3_chanxy_in = {wire_6313, wire_6174, wire_6329, wire_6238, wire_6299, wire_6298, wire_11729, wire_6719, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6510, wire_2109, wire_6283, wire_6282, wire_6269, wire_6268, wire_6233, wire_6232, wire_6253, wire_6252, wire_11727, wire_6691, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6622, wire_2109, wire_6327, wire_6230, wire_6297, wire_6296, wire_6169, wire_6168, wire_6267, wire_6266, wire_11725, wire_6693, wire_6625, wire_6624, wire_6614, wire_6585, wire_6584, wire_6545, wire_6544, wire_2109, wire_6225, wire_6224, wire_6325, wire_6222, wire_6311, wire_6166, wire_6281, wire_6280, wire_11723, wire_6695, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6606, wire_1599, wire_6295, wire_6294, wire_6251, wire_6250, wire_6161, wire_6160, wire_6265, wire_6264, wire_11721, wire_6697, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6598, wire_1599, wire_6309, wire_6158, wire_6279, wire_6278, wire_6217, wire_6216, wire_6249, wire_6248, wire_11719, wire_6699, wire_6617, wire_6616, wire_6590, wire_6577, wire_6576, wire_6537, wire_6536, wire_1599, wire_6153, wire_6152, wire_6307, wire_6150, wire_6323, wire_6214, wire_6293, wire_6292, wire_11717, wire_6701, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6582, wire_2113, wire_1599, wire_6277, wire_6276, wire_6263, wire_6262, wire_6209, wire_6208, wire_6247, wire_6246, wire_11715, wire_6703, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6574, wire_2113, wire_1599, wire_6321, wire_6206, wire_6291, wire_6290, wire_6145, wire_6144, wire_6261, wire_6260, wire_11713, wire_6705, wire_6609, wire_6608, wire_6569, wire_6568, wire_6566, wire_6529, wire_6528, wire_2113, wire_1599, wire_6201, wire_6200, wire_6319, wire_6198, wire_2113, wire_6305, wire_6142, wire_2113, wire_6275, wire_6274, wire_2113, wire_11711, wire_6707, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6558, wire_2113, wire_1595, wire_6289, wire_6288, wire_2113, wire_6245, wire_6244, wire_2113, wire_6137, wire_6136, wire_2113, wire_6259, wire_6258, wire_2109, wire_11709, wire_6709, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6550, wire_2113, wire_1595, wire_6303, wire_6134, wire_2109, wire_6273, wire_6272, wire_2109, wire_6193, wire_6192, wire_2109, wire_6243, wire_6242, wire_2109, wire_11707, wire_6711, wire_6601, wire_6600, wire_6561, wire_6560, wire_6542, wire_6521, wire_6520, wire_2113, wire_1595, wire_6129, wire_6128, wire_2109, wire_6301, wire_6126, wire_1599, wire_6317, wire_6190, wire_1599, wire_6287, wire_6286, wire_1599, wire_11705, wire_6713, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6534, wire_2109, wire_1595, wire_6271, wire_6270, wire_1599, wire_6257, wire_6256, wire_1599, wire_6185, wire_6184, wire_1599, wire_6241, wire_6240, wire_1595, wire_11703, wire_6715, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6526, wire_2109, wire_1595, wire_6315, wire_6182, wire_1595, wire_6285, wire_6284, wire_1595, wire_6121, wire_6120, wire_1595, wire_6255, wire_6254, wire_1595, wire_11701, wire_6717, wire_6593, wire_6592, wire_6553, wire_6552, wire_6518, wire_6513, wire_6512, wire_2109, wire_1595, wire_6177, wire_6176, wire_1595, wire_11337, wire_11308, wire_11307, wire_11306, wire_11267, wire_11266, wire_11227, wire_11226, wire_6628, wire_1638, wire_11335, wire_11305, wire_11304, wire_11265, wire_11264, wire_11225, wire_11224, wire_11196, wire_6620, wire_1638, wire_11333, wire_11303, wire_11302, wire_11263, wire_11262, wire_11223, wire_11222, wire_11204, wire_6612, wire_1638, wire_11331, wire_11299, wire_11298, wire_11259, wire_11258, wire_11219, wire_11218, wire_11212, wire_6604, wire_1598, wire_11329, wire_11297, wire_11296, wire_11257, wire_11256, wire_11220, wire_11217, wire_11216, wire_6596, wire_1598, wire_11327, wire_11295, wire_11294, wire_11255, wire_11254, wire_11228, wire_11215, wire_11214, wire_6588, wire_1598, wire_11325, wire_11291, wire_11290, wire_11251, wire_11250, wire_11236, wire_11211, wire_11210, wire_6580, wire_1642, wire_1598, wire_11323, wire_11289, wire_11288, wire_11249, wire_11248, wire_11244, wire_11209, wire_11208, wire_6572, wire_1642, wire_1598, wire_11321, wire_11287, wire_11286, wire_11252, wire_11247, wire_11246, wire_11207, wire_11206, wire_6564, wire_1642, wire_1598, wire_11319, wire_11283, wire_11282, wire_11260, wire_11243, wire_11242, wire_11203, wire_11202, wire_6556, wire_1642, wire_1594, wire_11317, wire_11281, wire_11280, wire_11268, wire_11241, wire_11240, wire_11201, wire_11200, wire_6548, wire_1642, wire_1594, wire_11315, wire_11279, wire_11278, wire_11276, wire_11239, wire_11238, wire_11199, wire_11198, wire_6540, wire_1642, wire_1594, wire_11313, wire_11284, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_6532, wire_1638, wire_1594, wire_11311, wire_11292, wire_11273, wire_11272, wire_11233, wire_11232, wire_11193, wire_11192, wire_6524, wire_1638, wire_1594, wire_11339, wire_11300, wire_11271, wire_11270, wire_11231, wire_11230, wire_11191, wire_11190, wire_6516, wire_1638, wire_1594, wire_11703, wire_11699, wire_11698, wire_11684, wire_11659, wire_11658, wire_11619, wire_11618, wire_6719, wire_1638, wire_11705, wire_11697, wire_11696, wire_11676, wire_11657, wire_11656, wire_11617, wire_11616, wire_6717, wire_1638, wire_11707, wire_11695, wire_11694, wire_11668, wire_11655, wire_11654, wire_11615, wire_11614, wire_6715, wire_1638, wire_11709, wire_11691, wire_11690, wire_11660, wire_11651, wire_11650, wire_11611, wire_11610, wire_6713, wire_1598, wire_11711, wire_11689, wire_11688, wire_11652, wire_11649, wire_11648, wire_11609, wire_11608, wire_6711, wire_1598, wire_11713, wire_11687, wire_11686, wire_11647, wire_11646, wire_11644, wire_11607, wire_11606, wire_6709, wire_1598, wire_11715, wire_11683, wire_11682, wire_11643, wire_11642, wire_11636, wire_11603, wire_11602, wire_6707, wire_1642, wire_1598, wire_11717, wire_11681, wire_11680, wire_11641, wire_11640, wire_11628, wire_11601, wire_11600, wire_6705, wire_1642, wire_1598, wire_11719, wire_11679, wire_11678, wire_11639, wire_11638, wire_11620, wire_11599, wire_11598, wire_6703, wire_1642, wire_1598, wire_11721, wire_11675, wire_11674, wire_11635, wire_11634, wire_11612, wire_11595, wire_11594, wire_6701, wire_1642, wire_1594, wire_11723, wire_11673, wire_11672, wire_11633, wire_11632, wire_11604, wire_11593, wire_11592, wire_6699, wire_1642, wire_1594, wire_11725, wire_11671, wire_11670, wire_11631, wire_11630, wire_11596, wire_11591, wire_11590, wire_6697, wire_1642, wire_1594, wire_11727, wire_11667, wire_11666, wire_11627, wire_11626, wire_11588, wire_11587, wire_11586, wire_6695, wire_1638, wire_1594, wire_11729, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_11580, wire_6693, wire_1638, wire_1594, wire_11701, wire_11692, wire_11663, wire_11662, wire_11623, wire_11622, wire_11583, wire_11582, wire_6691, wire_1638, wire_1594};
    // CHNAXY TOTAL: 621
    assign wire_6511 = lut_tile_1_3_chanxy_out[0];
    assign wire_6519 = lut_tile_1_3_chanxy_out[1];
    assign wire_6527 = lut_tile_1_3_chanxy_out[2];
    assign wire_6535 = lut_tile_1_3_chanxy_out[3];
    assign wire_6543 = lut_tile_1_3_chanxy_out[4];
    assign wire_6551 = lut_tile_1_3_chanxy_out[5];
    assign wire_6559 = lut_tile_1_3_chanxy_out[6];
    assign wire_6567 = lut_tile_1_3_chanxy_out[7];
    assign wire_6575 = lut_tile_1_3_chanxy_out[8];
    assign wire_6583 = lut_tile_1_3_chanxy_out[9];
    assign wire_6591 = lut_tile_1_3_chanxy_out[10];
    assign wire_6599 = lut_tile_1_3_chanxy_out[11];
    assign wire_6607 = lut_tile_1_3_chanxy_out[12];
    assign wire_6615 = lut_tile_1_3_chanxy_out[13];
    assign wire_6623 = lut_tile_1_3_chanxy_out[14];
    assign wire_6660 = lut_tile_1_3_chanxy_out[15];
    assign wire_6662 = lut_tile_1_3_chanxy_out[16];
    assign wire_6664 = lut_tile_1_3_chanxy_out[17];
    assign wire_6666 = lut_tile_1_3_chanxy_out[18];
    assign wire_6668 = lut_tile_1_3_chanxy_out[19];
    assign wire_6670 = lut_tile_1_3_chanxy_out[20];
    assign wire_6672 = lut_tile_1_3_chanxy_out[21];
    assign wire_6674 = lut_tile_1_3_chanxy_out[22];
    assign wire_6676 = lut_tile_1_3_chanxy_out[23];
    assign wire_6678 = lut_tile_1_3_chanxy_out[24];
    assign wire_6680 = lut_tile_1_3_chanxy_out[25];
    assign wire_6682 = lut_tile_1_3_chanxy_out[26];
    assign wire_6684 = lut_tile_1_3_chanxy_out[27];
    assign wire_6686 = lut_tile_1_3_chanxy_out[28];
    assign wire_6688 = lut_tile_1_3_chanxy_out[29];
    assign wire_11580 = lut_tile_1_3_chanxy_out[30];
    assign wire_11581 = lut_tile_1_3_chanxy_out[31];
    assign wire_11582 = lut_tile_1_3_chanxy_out[32];
    assign wire_11584 = lut_tile_1_3_chanxy_out[33];
    assign wire_11586 = lut_tile_1_3_chanxy_out[34];
    assign wire_11588 = lut_tile_1_3_chanxy_out[35];
    assign wire_11589 = lut_tile_1_3_chanxy_out[36];
    assign wire_11590 = lut_tile_1_3_chanxy_out[37];
    assign wire_11592 = lut_tile_1_3_chanxy_out[38];
    assign wire_11594 = lut_tile_1_3_chanxy_out[39];
    assign wire_11596 = lut_tile_1_3_chanxy_out[40];
    assign wire_11597 = lut_tile_1_3_chanxy_out[41];
    assign wire_11598 = lut_tile_1_3_chanxy_out[42];
    assign wire_11600 = lut_tile_1_3_chanxy_out[43];
    assign wire_11602 = lut_tile_1_3_chanxy_out[44];
    assign wire_11604 = lut_tile_1_3_chanxy_out[45];
    assign wire_11605 = lut_tile_1_3_chanxy_out[46];
    assign wire_11606 = lut_tile_1_3_chanxy_out[47];
    assign wire_11608 = lut_tile_1_3_chanxy_out[48];
    assign wire_11610 = lut_tile_1_3_chanxy_out[49];
    assign wire_11612 = lut_tile_1_3_chanxy_out[50];
    assign wire_11613 = lut_tile_1_3_chanxy_out[51];
    assign wire_11614 = lut_tile_1_3_chanxy_out[52];
    assign wire_11616 = lut_tile_1_3_chanxy_out[53];
    assign wire_11618 = lut_tile_1_3_chanxy_out[54];
    assign wire_11620 = lut_tile_1_3_chanxy_out[55];
    assign wire_11621 = lut_tile_1_3_chanxy_out[56];
    assign wire_11622 = lut_tile_1_3_chanxy_out[57];
    assign wire_11624 = lut_tile_1_3_chanxy_out[58];
    assign wire_11626 = lut_tile_1_3_chanxy_out[59];
    assign wire_11628 = lut_tile_1_3_chanxy_out[60];
    assign wire_11629 = lut_tile_1_3_chanxy_out[61];
    assign wire_11630 = lut_tile_1_3_chanxy_out[62];
    assign wire_11632 = lut_tile_1_3_chanxy_out[63];
    assign wire_11634 = lut_tile_1_3_chanxy_out[64];
    assign wire_11636 = lut_tile_1_3_chanxy_out[65];
    assign wire_11637 = lut_tile_1_3_chanxy_out[66];
    assign wire_11638 = lut_tile_1_3_chanxy_out[67];
    assign wire_11640 = lut_tile_1_3_chanxy_out[68];
    assign wire_11642 = lut_tile_1_3_chanxy_out[69];
    assign wire_11644 = lut_tile_1_3_chanxy_out[70];
    assign wire_11645 = lut_tile_1_3_chanxy_out[71];
    assign wire_11646 = lut_tile_1_3_chanxy_out[72];
    assign wire_11648 = lut_tile_1_3_chanxy_out[73];
    assign wire_11650 = lut_tile_1_3_chanxy_out[74];
    assign wire_11652 = lut_tile_1_3_chanxy_out[75];
    assign wire_11653 = lut_tile_1_3_chanxy_out[76];
    assign wire_11654 = lut_tile_1_3_chanxy_out[77];
    assign wire_11656 = lut_tile_1_3_chanxy_out[78];
    assign wire_11658 = lut_tile_1_3_chanxy_out[79];
    assign wire_11660 = lut_tile_1_3_chanxy_out[80];
    assign wire_11661 = lut_tile_1_3_chanxy_out[81];
    assign wire_11662 = lut_tile_1_3_chanxy_out[82];
    assign wire_11664 = lut_tile_1_3_chanxy_out[83];
    assign wire_11666 = lut_tile_1_3_chanxy_out[84];
    assign wire_11668 = lut_tile_1_3_chanxy_out[85];
    assign wire_11669 = lut_tile_1_3_chanxy_out[86];
    assign wire_11670 = lut_tile_1_3_chanxy_out[87];
    assign wire_11672 = lut_tile_1_3_chanxy_out[88];
    assign wire_11674 = lut_tile_1_3_chanxy_out[89];
    assign wire_11676 = lut_tile_1_3_chanxy_out[90];
    assign wire_11677 = lut_tile_1_3_chanxy_out[91];
    assign wire_11678 = lut_tile_1_3_chanxy_out[92];
    assign wire_11680 = lut_tile_1_3_chanxy_out[93];
    assign wire_11682 = lut_tile_1_3_chanxy_out[94];
    assign wire_11684 = lut_tile_1_3_chanxy_out[95];
    assign wire_11685 = lut_tile_1_3_chanxy_out[96];
    assign wire_11686 = lut_tile_1_3_chanxy_out[97];
    assign wire_11688 = lut_tile_1_3_chanxy_out[98];
    assign wire_11690 = lut_tile_1_3_chanxy_out[99];
    assign wire_11692 = lut_tile_1_3_chanxy_out[100];
    assign wire_11693 = lut_tile_1_3_chanxy_out[101];
    assign wire_11694 = lut_tile_1_3_chanxy_out[102];
    assign wire_11696 = lut_tile_1_3_chanxy_out[103];
    assign wire_11698 = lut_tile_1_3_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_4_chanxy_in = {wire_6313, wire_6312, wire_6329, wire_6328, wire_12119, wire_6749, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6512, wire_2625, wire_6299, wire_6298, wire_6283, wire_6282, wire_6269, wire_6268, wire_6359, wire_6232, wire_12117, wire_6721, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6624, wire_2625, wire_6253, wire_6252, wire_6327, wire_6326, wire_6297, wire_6296, wire_6343, wire_6168, wire_12115, wire_6723, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6616, wire_2625, wire_6267, wire_6266, wire_6357, wire_6224, wire_6325, wire_6324, wire_6311, wire_6310, wire_12113, wire_6725, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6608, wire_2115, wire_6281, wire_6280, wire_6295, wire_6294, wire_6251, wire_6250, wire_6341, wire_6160, wire_12111, wire_6727, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6600, wire_2115, wire_6265, wire_6264, wire_6309, wire_6308, wire_6279, wire_6278, wire_6355, wire_6216, wire_12109, wire_6729, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6592, wire_2115, wire_6249, wire_6248, wire_6339, wire_6152, wire_6307, wire_6306, wire_6323, wire_6322, wire_12107, wire_6731, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6584, wire_2629, wire_2115, wire_6293, wire_6292, wire_6277, wire_6276, wire_6263, wire_6262, wire_6353, wire_6208, wire_12105, wire_6733, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6576, wire_2629, wire_2115, wire_6247, wire_6246, wire_6321, wire_6320, wire_6291, wire_6290, wire_6337, wire_6144, wire_12103, wire_6735, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6568, wire_2629, wire_2115, wire_6261, wire_6260, wire_6351, wire_6200, wire_6319, wire_6318, wire_2629, wire_6305, wire_6304, wire_2629, wire_12101, wire_6737, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6560, wire_2629, wire_2111, wire_6275, wire_6274, wire_2629, wire_6289, wire_6288, wire_2629, wire_6245, wire_6244, wire_2629, wire_6335, wire_6136, wire_2629, wire_12099, wire_6739, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6552, wire_2629, wire_2111, wire_6259, wire_6258, wire_2625, wire_6303, wire_6302, wire_2625, wire_6273, wire_6272, wire_2625, wire_6349, wire_6192, wire_2625, wire_12097, wire_6741, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6544, wire_2629, wire_2111, wire_6243, wire_6242, wire_2625, wire_6333, wire_6128, wire_2625, wire_6301, wire_6300, wire_2115, wire_6317, wire_6316, wire_2115, wire_12095, wire_6743, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6536, wire_2625, wire_2111, wire_6287, wire_6286, wire_2115, wire_6271, wire_6270, wire_2115, wire_6257, wire_6256, wire_2115, wire_6347, wire_6184, wire_2115, wire_12093, wire_6745, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6528, wire_2625, wire_2111, wire_6241, wire_6240, wire_2111, wire_6315, wire_6314, wire_2111, wire_6285, wire_6284, wire_2111, wire_6331, wire_6120, wire_2111, wire_12091, wire_6747, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6520, wire_2625, wire_2111, wire_6255, wire_6254, wire_2111, wire_6345, wire_6176, wire_2111, wire_11727, wire_11699, wire_11698, wire_11692, wire_11659, wire_11658, wire_11619, wire_11618, wire_6622, wire_2154, wire_11725, wire_11697, wire_11696, wire_11657, wire_11656, wire_11617, wire_11616, wire_11580, wire_6614, wire_2154, wire_11723, wire_11695, wire_11694, wire_11655, wire_11654, wire_11615, wire_11614, wire_11588, wire_6606, wire_2154, wire_11721, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_11596, wire_6598, wire_2114, wire_11719, wire_11689, wire_11688, wire_11649, wire_11648, wire_11609, wire_11608, wire_11604, wire_6590, wire_2114, wire_11717, wire_11687, wire_11686, wire_11647, wire_11646, wire_11612, wire_11607, wire_11606, wire_6582, wire_2114, wire_11715, wire_11683, wire_11682, wire_11643, wire_11642, wire_11620, wire_11603, wire_11602, wire_6574, wire_2158, wire_2114, wire_11713, wire_11681, wire_11680, wire_11641, wire_11640, wire_11628, wire_11601, wire_11600, wire_6566, wire_2158, wire_2114, wire_11711, wire_11679, wire_11678, wire_11639, wire_11638, wire_11636, wire_11599, wire_11598, wire_6558, wire_2158, wire_2114, wire_11709, wire_11675, wire_11674, wire_11644, wire_11635, wire_11634, wire_11595, wire_11594, wire_6550, wire_2158, wire_2110, wire_11707, wire_11673, wire_11672, wire_11652, wire_11633, wire_11632, wire_11593, wire_11592, wire_6542, wire_2158, wire_2110, wire_11705, wire_11671, wire_11670, wire_11660, wire_11631, wire_11630, wire_11591, wire_11590, wire_6534, wire_2158, wire_2110, wire_11703, wire_11668, wire_11667, wire_11666, wire_11627, wire_11626, wire_11587, wire_11586, wire_6526, wire_2154, wire_2110, wire_11701, wire_11676, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_6518, wire_2154, wire_2110, wire_11729, wire_11684, wire_11663, wire_11662, wire_11623, wire_11622, wire_11583, wire_11582, wire_6510, wire_2154, wire_2110, wire_12093, wire_12089, wire_12088, wire_12076, wire_12049, wire_12048, wire_12009, wire_12008, wire_6749, wire_2154, wire_12095, wire_12087, wire_12086, wire_12068, wire_12047, wire_12046, wire_12007, wire_12006, wire_6747, wire_2154, wire_12097, wire_12083, wire_12082, wire_12060, wire_12043, wire_12042, wire_12003, wire_12002, wire_6745, wire_2154, wire_12099, wire_12081, wire_12080, wire_12052, wire_12041, wire_12040, wire_12001, wire_12000, wire_6743, wire_2114, wire_12101, wire_12079, wire_12078, wire_12044, wire_12039, wire_12038, wire_11999, wire_11998, wire_6741, wire_2114, wire_12103, wire_12075, wire_12074, wire_12036, wire_12035, wire_12034, wire_11995, wire_11994, wire_6739, wire_2114, wire_12105, wire_12073, wire_12072, wire_12033, wire_12032, wire_12028, wire_11993, wire_11992, wire_6737, wire_2158, wire_2114, wire_12107, wire_12071, wire_12070, wire_12031, wire_12030, wire_12020, wire_11991, wire_11990, wire_6735, wire_2158, wire_2114, wire_12109, wire_12067, wire_12066, wire_12027, wire_12026, wire_12012, wire_11987, wire_11986, wire_6733, wire_2158, wire_2114, wire_12111, wire_12065, wire_12064, wire_12025, wire_12024, wire_12004, wire_11985, wire_11984, wire_6731, wire_2158, wire_2110, wire_12113, wire_12063, wire_12062, wire_12023, wire_12022, wire_11996, wire_11983, wire_11982, wire_6729, wire_2158, wire_2110, wire_12115, wire_12059, wire_12058, wire_12019, wire_12018, wire_11988, wire_11979, wire_11978, wire_6727, wire_2158, wire_2110, wire_12117, wire_12057, wire_12056, wire_12017, wire_12016, wire_11980, wire_11977, wire_11976, wire_6725, wire_2154, wire_2110, wire_12119, wire_12055, wire_12054, wire_12015, wire_12014, wire_11975, wire_11974, wire_11972, wire_6723, wire_2154, wire_2110, wire_12091, wire_12084, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_6721, wire_2154, wire_2110};
    // CHNAXY TOTAL: 621
    assign wire_6513 = lut_tile_1_4_chanxy_out[0];
    assign wire_6521 = lut_tile_1_4_chanxy_out[1];
    assign wire_6529 = lut_tile_1_4_chanxy_out[2];
    assign wire_6537 = lut_tile_1_4_chanxy_out[3];
    assign wire_6545 = lut_tile_1_4_chanxy_out[4];
    assign wire_6553 = lut_tile_1_4_chanxy_out[5];
    assign wire_6561 = lut_tile_1_4_chanxy_out[6];
    assign wire_6569 = lut_tile_1_4_chanxy_out[7];
    assign wire_6577 = lut_tile_1_4_chanxy_out[8];
    assign wire_6585 = lut_tile_1_4_chanxy_out[9];
    assign wire_6593 = lut_tile_1_4_chanxy_out[10];
    assign wire_6601 = lut_tile_1_4_chanxy_out[11];
    assign wire_6609 = lut_tile_1_4_chanxy_out[12];
    assign wire_6617 = lut_tile_1_4_chanxy_out[13];
    assign wire_6625 = lut_tile_1_4_chanxy_out[14];
    assign wire_6690 = lut_tile_1_4_chanxy_out[15];
    assign wire_6692 = lut_tile_1_4_chanxy_out[16];
    assign wire_6694 = lut_tile_1_4_chanxy_out[17];
    assign wire_6696 = lut_tile_1_4_chanxy_out[18];
    assign wire_6698 = lut_tile_1_4_chanxy_out[19];
    assign wire_6700 = lut_tile_1_4_chanxy_out[20];
    assign wire_6702 = lut_tile_1_4_chanxy_out[21];
    assign wire_6704 = lut_tile_1_4_chanxy_out[22];
    assign wire_6706 = lut_tile_1_4_chanxy_out[23];
    assign wire_6708 = lut_tile_1_4_chanxy_out[24];
    assign wire_6710 = lut_tile_1_4_chanxy_out[25];
    assign wire_6712 = lut_tile_1_4_chanxy_out[26];
    assign wire_6714 = lut_tile_1_4_chanxy_out[27];
    assign wire_6716 = lut_tile_1_4_chanxy_out[28];
    assign wire_6718 = lut_tile_1_4_chanxy_out[29];
    assign wire_11970 = lut_tile_1_4_chanxy_out[30];
    assign wire_11972 = lut_tile_1_4_chanxy_out[31];
    assign wire_11973 = lut_tile_1_4_chanxy_out[32];
    assign wire_11974 = lut_tile_1_4_chanxy_out[33];
    assign wire_11976 = lut_tile_1_4_chanxy_out[34];
    assign wire_11978 = lut_tile_1_4_chanxy_out[35];
    assign wire_11980 = lut_tile_1_4_chanxy_out[36];
    assign wire_11981 = lut_tile_1_4_chanxy_out[37];
    assign wire_11982 = lut_tile_1_4_chanxy_out[38];
    assign wire_11984 = lut_tile_1_4_chanxy_out[39];
    assign wire_11986 = lut_tile_1_4_chanxy_out[40];
    assign wire_11988 = lut_tile_1_4_chanxy_out[41];
    assign wire_11989 = lut_tile_1_4_chanxy_out[42];
    assign wire_11990 = lut_tile_1_4_chanxy_out[43];
    assign wire_11992 = lut_tile_1_4_chanxy_out[44];
    assign wire_11994 = lut_tile_1_4_chanxy_out[45];
    assign wire_11996 = lut_tile_1_4_chanxy_out[46];
    assign wire_11997 = lut_tile_1_4_chanxy_out[47];
    assign wire_11998 = lut_tile_1_4_chanxy_out[48];
    assign wire_12000 = lut_tile_1_4_chanxy_out[49];
    assign wire_12002 = lut_tile_1_4_chanxy_out[50];
    assign wire_12004 = lut_tile_1_4_chanxy_out[51];
    assign wire_12005 = lut_tile_1_4_chanxy_out[52];
    assign wire_12006 = lut_tile_1_4_chanxy_out[53];
    assign wire_12008 = lut_tile_1_4_chanxy_out[54];
    assign wire_12010 = lut_tile_1_4_chanxy_out[55];
    assign wire_12012 = lut_tile_1_4_chanxy_out[56];
    assign wire_12013 = lut_tile_1_4_chanxy_out[57];
    assign wire_12014 = lut_tile_1_4_chanxy_out[58];
    assign wire_12016 = lut_tile_1_4_chanxy_out[59];
    assign wire_12018 = lut_tile_1_4_chanxy_out[60];
    assign wire_12020 = lut_tile_1_4_chanxy_out[61];
    assign wire_12021 = lut_tile_1_4_chanxy_out[62];
    assign wire_12022 = lut_tile_1_4_chanxy_out[63];
    assign wire_12024 = lut_tile_1_4_chanxy_out[64];
    assign wire_12026 = lut_tile_1_4_chanxy_out[65];
    assign wire_12028 = lut_tile_1_4_chanxy_out[66];
    assign wire_12029 = lut_tile_1_4_chanxy_out[67];
    assign wire_12030 = lut_tile_1_4_chanxy_out[68];
    assign wire_12032 = lut_tile_1_4_chanxy_out[69];
    assign wire_12034 = lut_tile_1_4_chanxy_out[70];
    assign wire_12036 = lut_tile_1_4_chanxy_out[71];
    assign wire_12037 = lut_tile_1_4_chanxy_out[72];
    assign wire_12038 = lut_tile_1_4_chanxy_out[73];
    assign wire_12040 = lut_tile_1_4_chanxy_out[74];
    assign wire_12042 = lut_tile_1_4_chanxy_out[75];
    assign wire_12044 = lut_tile_1_4_chanxy_out[76];
    assign wire_12045 = lut_tile_1_4_chanxy_out[77];
    assign wire_12046 = lut_tile_1_4_chanxy_out[78];
    assign wire_12048 = lut_tile_1_4_chanxy_out[79];
    assign wire_12050 = lut_tile_1_4_chanxy_out[80];
    assign wire_12052 = lut_tile_1_4_chanxy_out[81];
    assign wire_12053 = lut_tile_1_4_chanxy_out[82];
    assign wire_12054 = lut_tile_1_4_chanxy_out[83];
    assign wire_12056 = lut_tile_1_4_chanxy_out[84];
    assign wire_12058 = lut_tile_1_4_chanxy_out[85];
    assign wire_12060 = lut_tile_1_4_chanxy_out[86];
    assign wire_12061 = lut_tile_1_4_chanxy_out[87];
    assign wire_12062 = lut_tile_1_4_chanxy_out[88];
    assign wire_12064 = lut_tile_1_4_chanxy_out[89];
    assign wire_12066 = lut_tile_1_4_chanxy_out[90];
    assign wire_12068 = lut_tile_1_4_chanxy_out[91];
    assign wire_12069 = lut_tile_1_4_chanxy_out[92];
    assign wire_12070 = lut_tile_1_4_chanxy_out[93];
    assign wire_12072 = lut_tile_1_4_chanxy_out[94];
    assign wire_12074 = lut_tile_1_4_chanxy_out[95];
    assign wire_12076 = lut_tile_1_4_chanxy_out[96];
    assign wire_12077 = lut_tile_1_4_chanxy_out[97];
    assign wire_12078 = lut_tile_1_4_chanxy_out[98];
    assign wire_12080 = lut_tile_1_4_chanxy_out[99];
    assign wire_12082 = lut_tile_1_4_chanxy_out[100];
    assign wire_12084 = lut_tile_1_4_chanxy_out[101];
    assign wire_12085 = lut_tile_1_4_chanxy_out[102];
    assign wire_12086 = lut_tile_1_4_chanxy_out[103];
    assign wire_12088 = lut_tile_1_4_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_5_chanxy_in = {wire_6313, wire_6312, wire_12509, wire_6779, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6630, wire_3141, wire_6329, wire_6328, wire_6299, wire_6298, wire_6283, wire_6282, wire_6389, wire_6268, wire_12507, wire_6751, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6658, wire_3141, wire_6359, wire_6358, wire_6373, wire_6252, wire_6327, wire_6326, wire_6297, wire_6296, wire_12505, wire_6753, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6656, wire_3141, wire_6343, wire_6342, wire_6387, wire_6266, wire_6357, wire_6356, wire_6325, wire_6324, wire_12503, wire_6755, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6654, wire_2631, wire_6311, wire_6310, wire_6281, wire_6280, wire_6295, wire_6294, wire_6371, wire_6250, wire_12501, wire_6757, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6652, wire_2631, wire_6341, wire_6340, wire_6385, wire_6264, wire_6309, wire_6308, wire_6279, wire_6278, wire_12499, wire_6759, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6650, wire_2631, wire_6355, wire_6354, wire_6369, wire_6248, wire_6339, wire_6338, wire_6307, wire_6306, wire_12497, wire_6761, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6648, wire_3145, wire_2631, wire_6323, wire_6322, wire_6293, wire_6292, wire_6277, wire_6276, wire_6383, wire_6262, wire_12495, wire_6763, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6646, wire_3145, wire_2631, wire_6353, wire_6352, wire_6367, wire_6246, wire_6321, wire_6320, wire_6291, wire_6290, wire_12493, wire_6765, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6644, wire_3145, wire_2631, wire_6337, wire_6336, wire_6381, wire_6260, wire_6351, wire_6350, wire_6319, wire_6318, wire_3145, wire_12491, wire_6767, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6642, wire_3145, wire_2627, wire_6305, wire_6304, wire_3145, wire_6275, wire_6274, wire_3145, wire_6289, wire_6288, wire_3145, wire_6365, wire_6244, wire_3145, wire_12489, wire_6769, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6640, wire_3145, wire_2627, wire_6335, wire_6334, wire_3145, wire_6379, wire_6258, wire_3141, wire_6303, wire_6302, wire_3141, wire_6273, wire_6272, wire_3141, wire_12487, wire_6771, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6638, wire_3145, wire_2627, wire_6349, wire_6348, wire_3141, wire_6363, wire_6242, wire_3141, wire_6333, wire_6332, wire_3141, wire_6301, wire_6300, wire_2631, wire_12485, wire_6773, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6636, wire_3141, wire_2627, wire_6317, wire_6316, wire_2631, wire_6287, wire_6286, wire_2631, wire_6271, wire_6270, wire_2631, wire_6377, wire_6256, wire_2631, wire_12483, wire_6775, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6634, wire_3141, wire_2627, wire_6347, wire_6346, wire_2631, wire_6361, wire_6240, wire_2627, wire_6315, wire_6314, wire_2627, wire_6285, wire_6284, wire_2627, wire_12481, wire_6777, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6632, wire_3141, wire_2627, wire_6331, wire_6330, wire_2627, wire_6375, wire_6254, wire_2627, wire_6345, wire_6344, wire_2627, wire_12117, wire_12089, wire_12088, wire_12084, wire_12049, wire_12048, wire_12009, wire_12008, wire_6624, wire_2670, wire_12115, wire_12087, wire_12086, wire_12047, wire_12046, wire_12007, wire_12006, wire_11972, wire_6616, wire_2670, wire_12113, wire_12083, wire_12082, wire_12043, wire_12042, wire_12003, wire_12002, wire_11980, wire_6608, wire_2670, wire_12111, wire_12081, wire_12080, wire_12041, wire_12040, wire_12001, wire_12000, wire_11988, wire_6600, wire_2630, wire_12109, wire_12079, wire_12078, wire_12039, wire_12038, wire_11999, wire_11998, wire_11996, wire_6592, wire_2630, wire_12107, wire_12075, wire_12074, wire_12035, wire_12034, wire_12004, wire_11995, wire_11994, wire_6584, wire_2630, wire_12105, wire_12073, wire_12072, wire_12033, wire_12032, wire_12012, wire_11993, wire_11992, wire_6576, wire_2674, wire_2630, wire_12103, wire_12071, wire_12070, wire_12031, wire_12030, wire_12020, wire_11991, wire_11990, wire_6568, wire_2674, wire_2630, wire_12101, wire_12067, wire_12066, wire_12028, wire_12027, wire_12026, wire_11987, wire_11986, wire_6560, wire_2674, wire_2630, wire_12099, wire_12065, wire_12064, wire_12036, wire_12025, wire_12024, wire_11985, wire_11984, wire_6552, wire_2674, wire_2626, wire_12097, wire_12063, wire_12062, wire_12044, wire_12023, wire_12022, wire_11983, wire_11982, wire_6544, wire_2674, wire_2626, wire_12095, wire_12059, wire_12058, wire_12052, wire_12019, wire_12018, wire_11979, wire_11978, wire_6536, wire_2674, wire_2626, wire_12093, wire_12060, wire_12057, wire_12056, wire_12017, wire_12016, wire_11977, wire_11976, wire_6528, wire_2670, wire_2626, wire_12091, wire_12068, wire_12055, wire_12054, wire_12015, wire_12014, wire_11975, wire_11974, wire_6520, wire_2670, wire_2626, wire_12119, wire_12076, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_6512, wire_2670, wire_2626, wire_12483, wire_12479, wire_12478, wire_12468, wire_12439, wire_12438, wire_12399, wire_12398, wire_6779, wire_2670, wire_12485, wire_12475, wire_12474, wire_12460, wire_12435, wire_12434, wire_12395, wire_12394, wire_6777, wire_2670, wire_12487, wire_12473, wire_12472, wire_12452, wire_12433, wire_12432, wire_12393, wire_12392, wire_6775, wire_2670, wire_12489, wire_12471, wire_12470, wire_12444, wire_12431, wire_12430, wire_12391, wire_12390, wire_6773, wire_2630, wire_12491, wire_12467, wire_12466, wire_12436, wire_12427, wire_12426, wire_12387, wire_12386, wire_6771, wire_2630, wire_12493, wire_12465, wire_12464, wire_12428, wire_12425, wire_12424, wire_12385, wire_12384, wire_6769, wire_2630, wire_12495, wire_12463, wire_12462, wire_12423, wire_12422, wire_12420, wire_12383, wire_12382, wire_6767, wire_2674, wire_2630, wire_12497, wire_12459, wire_12458, wire_12419, wire_12418, wire_12412, wire_12379, wire_12378, wire_6765, wire_2674, wire_2630, wire_12499, wire_12457, wire_12456, wire_12417, wire_12416, wire_12404, wire_12377, wire_12376, wire_6763, wire_2674, wire_2630, wire_12501, wire_12455, wire_12454, wire_12415, wire_12414, wire_12396, wire_12375, wire_12374, wire_6761, wire_2674, wire_2626, wire_12503, wire_12451, wire_12450, wire_12411, wire_12410, wire_12388, wire_12371, wire_12370, wire_6759, wire_2674, wire_2626, wire_12505, wire_12449, wire_12448, wire_12409, wire_12408, wire_12380, wire_12369, wire_12368, wire_6757, wire_2674, wire_2626, wire_12507, wire_12447, wire_12446, wire_12407, wire_12406, wire_12372, wire_12367, wire_12366, wire_6755, wire_2670, wire_2626, wire_12509, wire_12443, wire_12442, wire_12403, wire_12402, wire_12364, wire_12363, wire_12362, wire_6753, wire_2670, wire_2626, wire_12481, wire_12476, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_6751, wire_2670, wire_2626};
    // CHNAXY TOTAL: 621
    assign wire_6631 = lut_tile_1_5_chanxy_out[0];
    assign wire_6633 = lut_tile_1_5_chanxy_out[1];
    assign wire_6635 = lut_tile_1_5_chanxy_out[2];
    assign wire_6637 = lut_tile_1_5_chanxy_out[3];
    assign wire_6639 = lut_tile_1_5_chanxy_out[4];
    assign wire_6641 = lut_tile_1_5_chanxy_out[5];
    assign wire_6643 = lut_tile_1_5_chanxy_out[6];
    assign wire_6645 = lut_tile_1_5_chanxy_out[7];
    assign wire_6647 = lut_tile_1_5_chanxy_out[8];
    assign wire_6649 = lut_tile_1_5_chanxy_out[9];
    assign wire_6651 = lut_tile_1_5_chanxy_out[10];
    assign wire_6653 = lut_tile_1_5_chanxy_out[11];
    assign wire_6655 = lut_tile_1_5_chanxy_out[12];
    assign wire_6657 = lut_tile_1_5_chanxy_out[13];
    assign wire_6659 = lut_tile_1_5_chanxy_out[14];
    assign wire_6720 = lut_tile_1_5_chanxy_out[15];
    assign wire_6722 = lut_tile_1_5_chanxy_out[16];
    assign wire_6724 = lut_tile_1_5_chanxy_out[17];
    assign wire_6726 = lut_tile_1_5_chanxy_out[18];
    assign wire_6728 = lut_tile_1_5_chanxy_out[19];
    assign wire_6730 = lut_tile_1_5_chanxy_out[20];
    assign wire_6732 = lut_tile_1_5_chanxy_out[21];
    assign wire_6734 = lut_tile_1_5_chanxy_out[22];
    assign wire_6736 = lut_tile_1_5_chanxy_out[23];
    assign wire_6738 = lut_tile_1_5_chanxy_out[24];
    assign wire_6740 = lut_tile_1_5_chanxy_out[25];
    assign wire_6742 = lut_tile_1_5_chanxy_out[26];
    assign wire_6744 = lut_tile_1_5_chanxy_out[27];
    assign wire_6746 = lut_tile_1_5_chanxy_out[28];
    assign wire_6748 = lut_tile_1_5_chanxy_out[29];
    assign wire_12360 = lut_tile_1_5_chanxy_out[30];
    assign wire_12362 = lut_tile_1_5_chanxy_out[31];
    assign wire_12364 = lut_tile_1_5_chanxy_out[32];
    assign wire_12365 = lut_tile_1_5_chanxy_out[33];
    assign wire_12366 = lut_tile_1_5_chanxy_out[34];
    assign wire_12368 = lut_tile_1_5_chanxy_out[35];
    assign wire_12370 = lut_tile_1_5_chanxy_out[36];
    assign wire_12372 = lut_tile_1_5_chanxy_out[37];
    assign wire_12373 = lut_tile_1_5_chanxy_out[38];
    assign wire_12374 = lut_tile_1_5_chanxy_out[39];
    assign wire_12376 = lut_tile_1_5_chanxy_out[40];
    assign wire_12378 = lut_tile_1_5_chanxy_out[41];
    assign wire_12380 = lut_tile_1_5_chanxy_out[42];
    assign wire_12381 = lut_tile_1_5_chanxy_out[43];
    assign wire_12382 = lut_tile_1_5_chanxy_out[44];
    assign wire_12384 = lut_tile_1_5_chanxy_out[45];
    assign wire_12386 = lut_tile_1_5_chanxy_out[46];
    assign wire_12388 = lut_tile_1_5_chanxy_out[47];
    assign wire_12389 = lut_tile_1_5_chanxy_out[48];
    assign wire_12390 = lut_tile_1_5_chanxy_out[49];
    assign wire_12392 = lut_tile_1_5_chanxy_out[50];
    assign wire_12394 = lut_tile_1_5_chanxy_out[51];
    assign wire_12396 = lut_tile_1_5_chanxy_out[52];
    assign wire_12397 = lut_tile_1_5_chanxy_out[53];
    assign wire_12398 = lut_tile_1_5_chanxy_out[54];
    assign wire_12400 = lut_tile_1_5_chanxy_out[55];
    assign wire_12402 = lut_tile_1_5_chanxy_out[56];
    assign wire_12404 = lut_tile_1_5_chanxy_out[57];
    assign wire_12405 = lut_tile_1_5_chanxy_out[58];
    assign wire_12406 = lut_tile_1_5_chanxy_out[59];
    assign wire_12408 = lut_tile_1_5_chanxy_out[60];
    assign wire_12410 = lut_tile_1_5_chanxy_out[61];
    assign wire_12412 = lut_tile_1_5_chanxy_out[62];
    assign wire_12413 = lut_tile_1_5_chanxy_out[63];
    assign wire_12414 = lut_tile_1_5_chanxy_out[64];
    assign wire_12416 = lut_tile_1_5_chanxy_out[65];
    assign wire_12418 = lut_tile_1_5_chanxy_out[66];
    assign wire_12420 = lut_tile_1_5_chanxy_out[67];
    assign wire_12421 = lut_tile_1_5_chanxy_out[68];
    assign wire_12422 = lut_tile_1_5_chanxy_out[69];
    assign wire_12424 = lut_tile_1_5_chanxy_out[70];
    assign wire_12426 = lut_tile_1_5_chanxy_out[71];
    assign wire_12428 = lut_tile_1_5_chanxy_out[72];
    assign wire_12429 = lut_tile_1_5_chanxy_out[73];
    assign wire_12430 = lut_tile_1_5_chanxy_out[74];
    assign wire_12432 = lut_tile_1_5_chanxy_out[75];
    assign wire_12434 = lut_tile_1_5_chanxy_out[76];
    assign wire_12436 = lut_tile_1_5_chanxy_out[77];
    assign wire_12437 = lut_tile_1_5_chanxy_out[78];
    assign wire_12438 = lut_tile_1_5_chanxy_out[79];
    assign wire_12440 = lut_tile_1_5_chanxy_out[80];
    assign wire_12442 = lut_tile_1_5_chanxy_out[81];
    assign wire_12444 = lut_tile_1_5_chanxy_out[82];
    assign wire_12445 = lut_tile_1_5_chanxy_out[83];
    assign wire_12446 = lut_tile_1_5_chanxy_out[84];
    assign wire_12448 = lut_tile_1_5_chanxy_out[85];
    assign wire_12450 = lut_tile_1_5_chanxy_out[86];
    assign wire_12452 = lut_tile_1_5_chanxy_out[87];
    assign wire_12453 = lut_tile_1_5_chanxy_out[88];
    assign wire_12454 = lut_tile_1_5_chanxy_out[89];
    assign wire_12456 = lut_tile_1_5_chanxy_out[90];
    assign wire_12458 = lut_tile_1_5_chanxy_out[91];
    assign wire_12460 = lut_tile_1_5_chanxy_out[92];
    assign wire_12461 = lut_tile_1_5_chanxy_out[93];
    assign wire_12462 = lut_tile_1_5_chanxy_out[94];
    assign wire_12464 = lut_tile_1_5_chanxy_out[95];
    assign wire_12466 = lut_tile_1_5_chanxy_out[96];
    assign wire_12468 = lut_tile_1_5_chanxy_out[97];
    assign wire_12469 = lut_tile_1_5_chanxy_out[98];
    assign wire_12470 = lut_tile_1_5_chanxy_out[99];
    assign wire_12472 = lut_tile_1_5_chanxy_out[100];
    assign wire_12474 = lut_tile_1_5_chanxy_out[101];
    assign wire_12476 = lut_tile_1_5_chanxy_out[102];
    assign wire_12477 = lut_tile_1_5_chanxy_out[103];
    assign wire_12478 = lut_tile_1_5_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_6_chanxy_in = {wire_12899, wire_6809, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6660, wire_3657, wire_6313, wire_6312, wire_6329, wire_6328, wire_6419, wire_6298, wire_6403, wire_6282, wire_12897, wire_6781, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6688, wire_3657, wire_6389, wire_6388, wire_6359, wire_6358, wire_6373, wire_6372, wire_6327, wire_6326, wire_12895, wire_6783, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6686, wire_3657, wire_6417, wire_6296, wire_6343, wire_6342, wire_6387, wire_6386, wire_6357, wire_6356, wire_12893, wire_6785, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6684, wire_3147, wire_6325, wire_6324, wire_6311, wire_6310, wire_6401, wire_6280, wire_6415, wire_6294, wire_12891, wire_6787, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6682, wire_3147, wire_6371, wire_6370, wire_6341, wire_6340, wire_6385, wire_6384, wire_6309, wire_6308, wire_12889, wire_6789, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6680, wire_3147, wire_6399, wire_6278, wire_6355, wire_6354, wire_6369, wire_6368, wire_6339, wire_6338, wire_12887, wire_6791, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6678, wire_3661, wire_3147, wire_6307, wire_6306, wire_6323, wire_6322, wire_6413, wire_6292, wire_6397, wire_6276, wire_12885, wire_6793, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6676, wire_3661, wire_3147, wire_6383, wire_6382, wire_6353, wire_6352, wire_6367, wire_6366, wire_6321, wire_6320, wire_12883, wire_6795, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6674, wire_3661, wire_3147, wire_6411, wire_6290, wire_6337, wire_6336, wire_6381, wire_6380, wire_6351, wire_6350, wire_12881, wire_6797, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6672, wire_3661, wire_3143, wire_6319, wire_6318, wire_3661, wire_6305, wire_6304, wire_3661, wire_6395, wire_6274, wire_3661, wire_6409, wire_6288, wire_3661, wire_12879, wire_6799, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6670, wire_3661, wire_3143, wire_6365, wire_6364, wire_3661, wire_6335, wire_6334, wire_3661, wire_6379, wire_6378, wire_3657, wire_6303, wire_6302, wire_3657, wire_12877, wire_6801, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6668, wire_3661, wire_3143, wire_6393, wire_6272, wire_3657, wire_6349, wire_6348, wire_3657, wire_6363, wire_6362, wire_3657, wire_6333, wire_6332, wire_3657, wire_12875, wire_6803, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6666, wire_3657, wire_3143, wire_6301, wire_6300, wire_3147, wire_6317, wire_6316, wire_3147, wire_6407, wire_6286, wire_3147, wire_6391, wire_6270, wire_3147, wire_12873, wire_6805, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6664, wire_3657, wire_3143, wire_6377, wire_6376, wire_3147, wire_6347, wire_6346, wire_3147, wire_6361, wire_6360, wire_3143, wire_6315, wire_6314, wire_3143, wire_12871, wire_6807, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6662, wire_3657, wire_3143, wire_6405, wire_6284, wire_3143, wire_6331, wire_6330, wire_3143, wire_6375, wire_6374, wire_3143, wire_6345, wire_6344, wire_3143, wire_12507, wire_12479, wire_12478, wire_12476, wire_12439, wire_12438, wire_12399, wire_12398, wire_6658, wire_3186, wire_12505, wire_12475, wire_12474, wire_12435, wire_12434, wire_12395, wire_12394, wire_12364, wire_6656, wire_3186, wire_12503, wire_12473, wire_12472, wire_12433, wire_12432, wire_12393, wire_12392, wire_12372, wire_6654, wire_3186, wire_12501, wire_12471, wire_12470, wire_12431, wire_12430, wire_12391, wire_12390, wire_12380, wire_6652, wire_3146, wire_12499, wire_12467, wire_12466, wire_12427, wire_12426, wire_12388, wire_12387, wire_12386, wire_6650, wire_3146, wire_12497, wire_12465, wire_12464, wire_12425, wire_12424, wire_12396, wire_12385, wire_12384, wire_6648, wire_3146, wire_12495, wire_12463, wire_12462, wire_12423, wire_12422, wire_12404, wire_12383, wire_12382, wire_6646, wire_3190, wire_3146, wire_12493, wire_12459, wire_12458, wire_12419, wire_12418, wire_12412, wire_12379, wire_12378, wire_6644, wire_3190, wire_3146, wire_12491, wire_12457, wire_12456, wire_12420, wire_12417, wire_12416, wire_12377, wire_12376, wire_6642, wire_3190, wire_3146, wire_12489, wire_12455, wire_12454, wire_12428, wire_12415, wire_12414, wire_12375, wire_12374, wire_6640, wire_3190, wire_3142, wire_12487, wire_12451, wire_12450, wire_12436, wire_12411, wire_12410, wire_12371, wire_12370, wire_6638, wire_3190, wire_3142, wire_12485, wire_12449, wire_12448, wire_12444, wire_12409, wire_12408, wire_12369, wire_12368, wire_6636, wire_3190, wire_3142, wire_12483, wire_12452, wire_12447, wire_12446, wire_12407, wire_12406, wire_12367, wire_12366, wire_6634, wire_3186, wire_3142, wire_12481, wire_12460, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_6632, wire_3186, wire_3142, wire_12509, wire_12468, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_6630, wire_3186, wire_3142, wire_12873, wire_12867, wire_12866, wire_12860, wire_12827, wire_12826, wire_12787, wire_12786, wire_6809, wire_3186, wire_12875, wire_12865, wire_12864, wire_12852, wire_12825, wire_12824, wire_12785, wire_12784, wire_6807, wire_3186, wire_12877, wire_12863, wire_12862, wire_12844, wire_12823, wire_12822, wire_12783, wire_12782, wire_6805, wire_3186, wire_12879, wire_12859, wire_12858, wire_12836, wire_12819, wire_12818, wire_12779, wire_12778, wire_6803, wire_3146, wire_12881, wire_12857, wire_12856, wire_12828, wire_12817, wire_12816, wire_12777, wire_12776, wire_6801, wire_3146, wire_12883, wire_12855, wire_12854, wire_12820, wire_12815, wire_12814, wire_12775, wire_12774, wire_6799, wire_3146, wire_12885, wire_12851, wire_12850, wire_12812, wire_12811, wire_12810, wire_12771, wire_12770, wire_6797, wire_3190, wire_3146, wire_12887, wire_12849, wire_12848, wire_12809, wire_12808, wire_12804, wire_12769, wire_12768, wire_6795, wire_3190, wire_3146, wire_12889, wire_12847, wire_12846, wire_12807, wire_12806, wire_12796, wire_12767, wire_12766, wire_6793, wire_3190, wire_3146, wire_12891, wire_12843, wire_12842, wire_12803, wire_12802, wire_12788, wire_12763, wire_12762, wire_6791, wire_3190, wire_3142, wire_12893, wire_12841, wire_12840, wire_12801, wire_12800, wire_12780, wire_12761, wire_12760, wire_6789, wire_3190, wire_3142, wire_12895, wire_12839, wire_12838, wire_12799, wire_12798, wire_12772, wire_12759, wire_12758, wire_6787, wire_3190, wire_3142, wire_12897, wire_12835, wire_12834, wire_12795, wire_12794, wire_12764, wire_12755, wire_12754, wire_6785, wire_3186, wire_3142, wire_12899, wire_12833, wire_12832, wire_12793, wire_12792, wire_12756, wire_12753, wire_12752, wire_6783, wire_3186, wire_3142, wire_12871, wire_12868, wire_12831, wire_12830, wire_12791, wire_12790, wire_12751, wire_12750, wire_6781, wire_3186, wire_3142};
    // CHNAXY TOTAL: 621
    assign wire_6661 = lut_tile_1_6_chanxy_out[0];
    assign wire_6663 = lut_tile_1_6_chanxy_out[1];
    assign wire_6665 = lut_tile_1_6_chanxy_out[2];
    assign wire_6667 = lut_tile_1_6_chanxy_out[3];
    assign wire_6669 = lut_tile_1_6_chanxy_out[4];
    assign wire_6671 = lut_tile_1_6_chanxy_out[5];
    assign wire_6673 = lut_tile_1_6_chanxy_out[6];
    assign wire_6675 = lut_tile_1_6_chanxy_out[7];
    assign wire_6677 = lut_tile_1_6_chanxy_out[8];
    assign wire_6679 = lut_tile_1_6_chanxy_out[9];
    assign wire_6681 = lut_tile_1_6_chanxy_out[10];
    assign wire_6683 = lut_tile_1_6_chanxy_out[11];
    assign wire_6685 = lut_tile_1_6_chanxy_out[12];
    assign wire_6687 = lut_tile_1_6_chanxy_out[13];
    assign wire_6689 = lut_tile_1_6_chanxy_out[14];
    assign wire_6750 = lut_tile_1_6_chanxy_out[15];
    assign wire_6752 = lut_tile_1_6_chanxy_out[16];
    assign wire_6754 = lut_tile_1_6_chanxy_out[17];
    assign wire_6756 = lut_tile_1_6_chanxy_out[18];
    assign wire_6758 = lut_tile_1_6_chanxy_out[19];
    assign wire_6760 = lut_tile_1_6_chanxy_out[20];
    assign wire_6762 = lut_tile_1_6_chanxy_out[21];
    assign wire_6764 = lut_tile_1_6_chanxy_out[22];
    assign wire_6766 = lut_tile_1_6_chanxy_out[23];
    assign wire_6768 = lut_tile_1_6_chanxy_out[24];
    assign wire_6770 = lut_tile_1_6_chanxy_out[25];
    assign wire_6772 = lut_tile_1_6_chanxy_out[26];
    assign wire_6774 = lut_tile_1_6_chanxy_out[27];
    assign wire_6776 = lut_tile_1_6_chanxy_out[28];
    assign wire_6778 = lut_tile_1_6_chanxy_out[29];
    assign wire_12750 = lut_tile_1_6_chanxy_out[30];
    assign wire_12752 = lut_tile_1_6_chanxy_out[31];
    assign wire_12754 = lut_tile_1_6_chanxy_out[32];
    assign wire_12756 = lut_tile_1_6_chanxy_out[33];
    assign wire_12757 = lut_tile_1_6_chanxy_out[34];
    assign wire_12758 = lut_tile_1_6_chanxy_out[35];
    assign wire_12760 = lut_tile_1_6_chanxy_out[36];
    assign wire_12762 = lut_tile_1_6_chanxy_out[37];
    assign wire_12764 = lut_tile_1_6_chanxy_out[38];
    assign wire_12765 = lut_tile_1_6_chanxy_out[39];
    assign wire_12766 = lut_tile_1_6_chanxy_out[40];
    assign wire_12768 = lut_tile_1_6_chanxy_out[41];
    assign wire_12770 = lut_tile_1_6_chanxy_out[42];
    assign wire_12772 = lut_tile_1_6_chanxy_out[43];
    assign wire_12773 = lut_tile_1_6_chanxy_out[44];
    assign wire_12774 = lut_tile_1_6_chanxy_out[45];
    assign wire_12776 = lut_tile_1_6_chanxy_out[46];
    assign wire_12778 = lut_tile_1_6_chanxy_out[47];
    assign wire_12780 = lut_tile_1_6_chanxy_out[48];
    assign wire_12781 = lut_tile_1_6_chanxy_out[49];
    assign wire_12782 = lut_tile_1_6_chanxy_out[50];
    assign wire_12784 = lut_tile_1_6_chanxy_out[51];
    assign wire_12786 = lut_tile_1_6_chanxy_out[52];
    assign wire_12788 = lut_tile_1_6_chanxy_out[53];
    assign wire_12789 = lut_tile_1_6_chanxy_out[54];
    assign wire_12790 = lut_tile_1_6_chanxy_out[55];
    assign wire_12792 = lut_tile_1_6_chanxy_out[56];
    assign wire_12794 = lut_tile_1_6_chanxy_out[57];
    assign wire_12796 = lut_tile_1_6_chanxy_out[58];
    assign wire_12797 = lut_tile_1_6_chanxy_out[59];
    assign wire_12798 = lut_tile_1_6_chanxy_out[60];
    assign wire_12800 = lut_tile_1_6_chanxy_out[61];
    assign wire_12802 = lut_tile_1_6_chanxy_out[62];
    assign wire_12804 = lut_tile_1_6_chanxy_out[63];
    assign wire_12805 = lut_tile_1_6_chanxy_out[64];
    assign wire_12806 = lut_tile_1_6_chanxy_out[65];
    assign wire_12808 = lut_tile_1_6_chanxy_out[66];
    assign wire_12810 = lut_tile_1_6_chanxy_out[67];
    assign wire_12812 = lut_tile_1_6_chanxy_out[68];
    assign wire_12813 = lut_tile_1_6_chanxy_out[69];
    assign wire_12814 = lut_tile_1_6_chanxy_out[70];
    assign wire_12816 = lut_tile_1_6_chanxy_out[71];
    assign wire_12818 = lut_tile_1_6_chanxy_out[72];
    assign wire_12820 = lut_tile_1_6_chanxy_out[73];
    assign wire_12821 = lut_tile_1_6_chanxy_out[74];
    assign wire_12822 = lut_tile_1_6_chanxy_out[75];
    assign wire_12824 = lut_tile_1_6_chanxy_out[76];
    assign wire_12826 = lut_tile_1_6_chanxy_out[77];
    assign wire_12828 = lut_tile_1_6_chanxy_out[78];
    assign wire_12829 = lut_tile_1_6_chanxy_out[79];
    assign wire_12830 = lut_tile_1_6_chanxy_out[80];
    assign wire_12832 = lut_tile_1_6_chanxy_out[81];
    assign wire_12834 = lut_tile_1_6_chanxy_out[82];
    assign wire_12836 = lut_tile_1_6_chanxy_out[83];
    assign wire_12837 = lut_tile_1_6_chanxy_out[84];
    assign wire_12838 = lut_tile_1_6_chanxy_out[85];
    assign wire_12840 = lut_tile_1_6_chanxy_out[86];
    assign wire_12842 = lut_tile_1_6_chanxy_out[87];
    assign wire_12844 = lut_tile_1_6_chanxy_out[88];
    assign wire_12845 = lut_tile_1_6_chanxy_out[89];
    assign wire_12846 = lut_tile_1_6_chanxy_out[90];
    assign wire_12848 = lut_tile_1_6_chanxy_out[91];
    assign wire_12850 = lut_tile_1_6_chanxy_out[92];
    assign wire_12852 = lut_tile_1_6_chanxy_out[93];
    assign wire_12853 = lut_tile_1_6_chanxy_out[94];
    assign wire_12854 = lut_tile_1_6_chanxy_out[95];
    assign wire_12856 = lut_tile_1_6_chanxy_out[96];
    assign wire_12858 = lut_tile_1_6_chanxy_out[97];
    assign wire_12860 = lut_tile_1_6_chanxy_out[98];
    assign wire_12861 = lut_tile_1_6_chanxy_out[99];
    assign wire_12862 = lut_tile_1_6_chanxy_out[100];
    assign wire_12864 = lut_tile_1_6_chanxy_out[101];
    assign wire_12866 = lut_tile_1_6_chanxy_out[102];
    assign wire_12868 = lut_tile_1_6_chanxy_out[103];
    assign wire_12869 = lut_tile_1_6_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_7_chanxy_in = {wire_6433, wire_6312, wire_6449, wire_6328, wire_6419, wire_6418, wire_13289, wire_6839, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6690, wire_4173, wire_6403, wire_6402, wire_6389, wire_6388, wire_6359, wire_6358, wire_6373, wire_6372, wire_13287, wire_6811, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6718, wire_4173, wire_6447, wire_6326, wire_6417, wire_6416, wire_6343, wire_6342, wire_6387, wire_6386, wire_13285, wire_6813, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6716, wire_4173, wire_6357, wire_6356, wire_6445, wire_6324, wire_6431, wire_6310, wire_6401, wire_6400, wire_13283, wire_6815, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6714, wire_3663, wire_6415, wire_6414, wire_6371, wire_6370, wire_6341, wire_6340, wire_6385, wire_6384, wire_13281, wire_6817, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6712, wire_3663, wire_6429, wire_6308, wire_6399, wire_6398, wire_6355, wire_6354, wire_6369, wire_6368, wire_13279, wire_6819, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6710, wire_3663, wire_6339, wire_6338, wire_6427, wire_6306, wire_6443, wire_6322, wire_6413, wire_6412, wire_13277, wire_6821, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6708, wire_4177, wire_3663, wire_6397, wire_6396, wire_6383, wire_6382, wire_6353, wire_6352, wire_6367, wire_6366, wire_13275, wire_6823, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6706, wire_4177, wire_3663, wire_6441, wire_6320, wire_6411, wire_6410, wire_6337, wire_6336, wire_6381, wire_6380, wire_13273, wire_6825, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6704, wire_4177, wire_3663, wire_6351, wire_6350, wire_6439, wire_6318, wire_4177, wire_6425, wire_6304, wire_4177, wire_6395, wire_6394, wire_4177, wire_13271, wire_6827, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6702, wire_4177, wire_3659, wire_6409, wire_6408, wire_4177, wire_6365, wire_6364, wire_4177, wire_6335, wire_6334, wire_4177, wire_6379, wire_6378, wire_4173, wire_13269, wire_6829, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6700, wire_4177, wire_3659, wire_6423, wire_6302, wire_4173, wire_6393, wire_6392, wire_4173, wire_6349, wire_6348, wire_4173, wire_6363, wire_6362, wire_4173, wire_13267, wire_6831, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6698, wire_4177, wire_3659, wire_6333, wire_6332, wire_4173, wire_6421, wire_6300, wire_3663, wire_6437, wire_6316, wire_3663, wire_6407, wire_6406, wire_3663, wire_13265, wire_6833, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6696, wire_4173, wire_3659, wire_6391, wire_6390, wire_3663, wire_6377, wire_6376, wire_3663, wire_6347, wire_6346, wire_3663, wire_6361, wire_6360, wire_3659, wire_13263, wire_6835, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6694, wire_4173, wire_3659, wire_6435, wire_6314, wire_3659, wire_6405, wire_6404, wire_3659, wire_6331, wire_6330, wire_3659, wire_6375, wire_6374, wire_3659, wire_13261, wire_6837, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6692, wire_4173, wire_3659, wire_6345, wire_6344, wire_3659, wire_12897, wire_12868, wire_12867, wire_12866, wire_12827, wire_12826, wire_12787, wire_12786, wire_6688, wire_3702, wire_12895, wire_12865, wire_12864, wire_12825, wire_12824, wire_12785, wire_12784, wire_12756, wire_6686, wire_3702, wire_12893, wire_12863, wire_12862, wire_12823, wire_12822, wire_12783, wire_12782, wire_12764, wire_6684, wire_3702, wire_12891, wire_12859, wire_12858, wire_12819, wire_12818, wire_12779, wire_12778, wire_12772, wire_6682, wire_3662, wire_12889, wire_12857, wire_12856, wire_12817, wire_12816, wire_12780, wire_12777, wire_12776, wire_6680, wire_3662, wire_12887, wire_12855, wire_12854, wire_12815, wire_12814, wire_12788, wire_12775, wire_12774, wire_6678, wire_3662, wire_12885, wire_12851, wire_12850, wire_12811, wire_12810, wire_12796, wire_12771, wire_12770, wire_6676, wire_3706, wire_3662, wire_12883, wire_12849, wire_12848, wire_12809, wire_12808, wire_12804, wire_12769, wire_12768, wire_6674, wire_3706, wire_3662, wire_12881, wire_12847, wire_12846, wire_12812, wire_12807, wire_12806, wire_12767, wire_12766, wire_6672, wire_3706, wire_3662, wire_12879, wire_12843, wire_12842, wire_12820, wire_12803, wire_12802, wire_12763, wire_12762, wire_6670, wire_3706, wire_3658, wire_12877, wire_12841, wire_12840, wire_12828, wire_12801, wire_12800, wire_12761, wire_12760, wire_6668, wire_3706, wire_3658, wire_12875, wire_12839, wire_12838, wire_12836, wire_12799, wire_12798, wire_12759, wire_12758, wire_6666, wire_3706, wire_3658, wire_12873, wire_12844, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_6664, wire_3702, wire_3658, wire_12871, wire_12852, wire_12833, wire_12832, wire_12793, wire_12792, wire_12753, wire_12752, wire_6662, wire_3702, wire_3658, wire_12899, wire_12860, wire_12831, wire_12830, wire_12791, wire_12790, wire_12751, wire_12750, wire_6660, wire_3702, wire_3658, wire_13263, wire_13259, wire_13258, wire_13244, wire_13219, wire_13218, wire_13179, wire_13178, wire_6839, wire_3702, wire_13265, wire_13257, wire_13256, wire_13236, wire_13217, wire_13216, wire_13177, wire_13176, wire_6837, wire_3702, wire_13267, wire_13255, wire_13254, wire_13228, wire_13215, wire_13214, wire_13175, wire_13174, wire_6835, wire_3702, wire_13269, wire_13251, wire_13250, wire_13220, wire_13211, wire_13210, wire_13171, wire_13170, wire_6833, wire_3662, wire_13271, wire_13249, wire_13248, wire_13212, wire_13209, wire_13208, wire_13169, wire_13168, wire_6831, wire_3662, wire_13273, wire_13247, wire_13246, wire_13207, wire_13206, wire_13204, wire_13167, wire_13166, wire_6829, wire_3662, wire_13275, wire_13243, wire_13242, wire_13203, wire_13202, wire_13196, wire_13163, wire_13162, wire_6827, wire_3706, wire_3662, wire_13277, wire_13241, wire_13240, wire_13201, wire_13200, wire_13188, wire_13161, wire_13160, wire_6825, wire_3706, wire_3662, wire_13279, wire_13239, wire_13238, wire_13199, wire_13198, wire_13180, wire_13159, wire_13158, wire_6823, wire_3706, wire_3662, wire_13281, wire_13235, wire_13234, wire_13195, wire_13194, wire_13172, wire_13155, wire_13154, wire_6821, wire_3706, wire_3658, wire_13283, wire_13233, wire_13232, wire_13193, wire_13192, wire_13164, wire_13153, wire_13152, wire_6819, wire_3706, wire_3658, wire_13285, wire_13231, wire_13230, wire_13191, wire_13190, wire_13156, wire_13151, wire_13150, wire_6817, wire_3706, wire_3658, wire_13287, wire_13227, wire_13226, wire_13187, wire_13186, wire_13148, wire_13147, wire_13146, wire_6815, wire_3702, wire_3658, wire_13289, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_13140, wire_6813, wire_3702, wire_3658, wire_13261, wire_13252, wire_13223, wire_13222, wire_13183, wire_13182, wire_13143, wire_13142, wire_6811, wire_3702, wire_3658};
    // CHNAXY TOTAL: 621
    assign wire_6691 = lut_tile_1_7_chanxy_out[0];
    assign wire_6693 = lut_tile_1_7_chanxy_out[1];
    assign wire_6695 = lut_tile_1_7_chanxy_out[2];
    assign wire_6697 = lut_tile_1_7_chanxy_out[3];
    assign wire_6699 = lut_tile_1_7_chanxy_out[4];
    assign wire_6701 = lut_tile_1_7_chanxy_out[5];
    assign wire_6703 = lut_tile_1_7_chanxy_out[6];
    assign wire_6705 = lut_tile_1_7_chanxy_out[7];
    assign wire_6707 = lut_tile_1_7_chanxy_out[8];
    assign wire_6709 = lut_tile_1_7_chanxy_out[9];
    assign wire_6711 = lut_tile_1_7_chanxy_out[10];
    assign wire_6713 = lut_tile_1_7_chanxy_out[11];
    assign wire_6715 = lut_tile_1_7_chanxy_out[12];
    assign wire_6717 = lut_tile_1_7_chanxy_out[13];
    assign wire_6719 = lut_tile_1_7_chanxy_out[14];
    assign wire_6780 = lut_tile_1_7_chanxy_out[15];
    assign wire_6782 = lut_tile_1_7_chanxy_out[16];
    assign wire_6784 = lut_tile_1_7_chanxy_out[17];
    assign wire_6786 = lut_tile_1_7_chanxy_out[18];
    assign wire_6788 = lut_tile_1_7_chanxy_out[19];
    assign wire_6790 = lut_tile_1_7_chanxy_out[20];
    assign wire_6792 = lut_tile_1_7_chanxy_out[21];
    assign wire_6794 = lut_tile_1_7_chanxy_out[22];
    assign wire_6796 = lut_tile_1_7_chanxy_out[23];
    assign wire_6798 = lut_tile_1_7_chanxy_out[24];
    assign wire_6800 = lut_tile_1_7_chanxy_out[25];
    assign wire_6802 = lut_tile_1_7_chanxy_out[26];
    assign wire_6804 = lut_tile_1_7_chanxy_out[27];
    assign wire_6806 = lut_tile_1_7_chanxy_out[28];
    assign wire_6808 = lut_tile_1_7_chanxy_out[29];
    assign wire_13140 = lut_tile_1_7_chanxy_out[30];
    assign wire_13141 = lut_tile_1_7_chanxy_out[31];
    assign wire_13142 = lut_tile_1_7_chanxy_out[32];
    assign wire_13144 = lut_tile_1_7_chanxy_out[33];
    assign wire_13146 = lut_tile_1_7_chanxy_out[34];
    assign wire_13148 = lut_tile_1_7_chanxy_out[35];
    assign wire_13149 = lut_tile_1_7_chanxy_out[36];
    assign wire_13150 = lut_tile_1_7_chanxy_out[37];
    assign wire_13152 = lut_tile_1_7_chanxy_out[38];
    assign wire_13154 = lut_tile_1_7_chanxy_out[39];
    assign wire_13156 = lut_tile_1_7_chanxy_out[40];
    assign wire_13157 = lut_tile_1_7_chanxy_out[41];
    assign wire_13158 = lut_tile_1_7_chanxy_out[42];
    assign wire_13160 = lut_tile_1_7_chanxy_out[43];
    assign wire_13162 = lut_tile_1_7_chanxy_out[44];
    assign wire_13164 = lut_tile_1_7_chanxy_out[45];
    assign wire_13165 = lut_tile_1_7_chanxy_out[46];
    assign wire_13166 = lut_tile_1_7_chanxy_out[47];
    assign wire_13168 = lut_tile_1_7_chanxy_out[48];
    assign wire_13170 = lut_tile_1_7_chanxy_out[49];
    assign wire_13172 = lut_tile_1_7_chanxy_out[50];
    assign wire_13173 = lut_tile_1_7_chanxy_out[51];
    assign wire_13174 = lut_tile_1_7_chanxy_out[52];
    assign wire_13176 = lut_tile_1_7_chanxy_out[53];
    assign wire_13178 = lut_tile_1_7_chanxy_out[54];
    assign wire_13180 = lut_tile_1_7_chanxy_out[55];
    assign wire_13181 = lut_tile_1_7_chanxy_out[56];
    assign wire_13182 = lut_tile_1_7_chanxy_out[57];
    assign wire_13184 = lut_tile_1_7_chanxy_out[58];
    assign wire_13186 = lut_tile_1_7_chanxy_out[59];
    assign wire_13188 = lut_tile_1_7_chanxy_out[60];
    assign wire_13189 = lut_tile_1_7_chanxy_out[61];
    assign wire_13190 = lut_tile_1_7_chanxy_out[62];
    assign wire_13192 = lut_tile_1_7_chanxy_out[63];
    assign wire_13194 = lut_tile_1_7_chanxy_out[64];
    assign wire_13196 = lut_tile_1_7_chanxy_out[65];
    assign wire_13197 = lut_tile_1_7_chanxy_out[66];
    assign wire_13198 = lut_tile_1_7_chanxy_out[67];
    assign wire_13200 = lut_tile_1_7_chanxy_out[68];
    assign wire_13202 = lut_tile_1_7_chanxy_out[69];
    assign wire_13204 = lut_tile_1_7_chanxy_out[70];
    assign wire_13205 = lut_tile_1_7_chanxy_out[71];
    assign wire_13206 = lut_tile_1_7_chanxy_out[72];
    assign wire_13208 = lut_tile_1_7_chanxy_out[73];
    assign wire_13210 = lut_tile_1_7_chanxy_out[74];
    assign wire_13212 = lut_tile_1_7_chanxy_out[75];
    assign wire_13213 = lut_tile_1_7_chanxy_out[76];
    assign wire_13214 = lut_tile_1_7_chanxy_out[77];
    assign wire_13216 = lut_tile_1_7_chanxy_out[78];
    assign wire_13218 = lut_tile_1_7_chanxy_out[79];
    assign wire_13220 = lut_tile_1_7_chanxy_out[80];
    assign wire_13221 = lut_tile_1_7_chanxy_out[81];
    assign wire_13222 = lut_tile_1_7_chanxy_out[82];
    assign wire_13224 = lut_tile_1_7_chanxy_out[83];
    assign wire_13226 = lut_tile_1_7_chanxy_out[84];
    assign wire_13228 = lut_tile_1_7_chanxy_out[85];
    assign wire_13229 = lut_tile_1_7_chanxy_out[86];
    assign wire_13230 = lut_tile_1_7_chanxy_out[87];
    assign wire_13232 = lut_tile_1_7_chanxy_out[88];
    assign wire_13234 = lut_tile_1_7_chanxy_out[89];
    assign wire_13236 = lut_tile_1_7_chanxy_out[90];
    assign wire_13237 = lut_tile_1_7_chanxy_out[91];
    assign wire_13238 = lut_tile_1_7_chanxy_out[92];
    assign wire_13240 = lut_tile_1_7_chanxy_out[93];
    assign wire_13242 = lut_tile_1_7_chanxy_out[94];
    assign wire_13244 = lut_tile_1_7_chanxy_out[95];
    assign wire_13245 = lut_tile_1_7_chanxy_out[96];
    assign wire_13246 = lut_tile_1_7_chanxy_out[97];
    assign wire_13248 = lut_tile_1_7_chanxy_out[98];
    assign wire_13250 = lut_tile_1_7_chanxy_out[99];
    assign wire_13252 = lut_tile_1_7_chanxy_out[100];
    assign wire_13253 = lut_tile_1_7_chanxy_out[101];
    assign wire_13254 = lut_tile_1_7_chanxy_out[102];
    assign wire_13256 = lut_tile_1_7_chanxy_out[103];
    assign wire_13258 = lut_tile_1_7_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_8_chanxy_in = {wire_6433, wire_6432, wire_6449, wire_6448, wire_13679, wire_6869, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6720, wire_4689, wire_6419, wire_6418, wire_6403, wire_6402, wire_6389, wire_6388, wire_6479, wire_6358, wire_13677, wire_6841, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6748, wire_4689, wire_6373, wire_6372, wire_6447, wire_6446, wire_6417, wire_6416, wire_6463, wire_6342, wire_13675, wire_6843, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6746, wire_4689, wire_6387, wire_6386, wire_6477, wire_6356, wire_6445, wire_6444, wire_6431, wire_6430, wire_13673, wire_6845, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6744, wire_4179, wire_6401, wire_6400, wire_6415, wire_6414, wire_6371, wire_6370, wire_6461, wire_6340, wire_13671, wire_6847, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6742, wire_4179, wire_6385, wire_6384, wire_6429, wire_6428, wire_6399, wire_6398, wire_6475, wire_6354, wire_13669, wire_6849, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6740, wire_4179, wire_6369, wire_6368, wire_6459, wire_6338, wire_6427, wire_6426, wire_6443, wire_6442, wire_13667, wire_6851, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6738, wire_4693, wire_4179, wire_6413, wire_6412, wire_6397, wire_6396, wire_6383, wire_6382, wire_6473, wire_6352, wire_13665, wire_6853, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6736, wire_4693, wire_4179, wire_6367, wire_6366, wire_6441, wire_6440, wire_6411, wire_6410, wire_6457, wire_6336, wire_13663, wire_6855, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6734, wire_4693, wire_4179, wire_6381, wire_6380, wire_6471, wire_6350, wire_6439, wire_6438, wire_4693, wire_6425, wire_6424, wire_4693, wire_13661, wire_6857, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6732, wire_4693, wire_4175, wire_6395, wire_6394, wire_4693, wire_6409, wire_6408, wire_4693, wire_6365, wire_6364, wire_4693, wire_6455, wire_6334, wire_4693, wire_13659, wire_6859, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6730, wire_4693, wire_4175, wire_6379, wire_6378, wire_4689, wire_6423, wire_6422, wire_4689, wire_6393, wire_6392, wire_4689, wire_6469, wire_6348, wire_4689, wire_13657, wire_6861, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6728, wire_4693, wire_4175, wire_6363, wire_6362, wire_4689, wire_6453, wire_6332, wire_4689, wire_6421, wire_6420, wire_4179, wire_6437, wire_6436, wire_4179, wire_13655, wire_6863, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6726, wire_4689, wire_4175, wire_6407, wire_6406, wire_4179, wire_6391, wire_6390, wire_4179, wire_6377, wire_6376, wire_4179, wire_6467, wire_6346, wire_4179, wire_13653, wire_6865, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6724, wire_4689, wire_4175, wire_6361, wire_6360, wire_4175, wire_6435, wire_6434, wire_4175, wire_6405, wire_6404, wire_4175, wire_6451, wire_6330, wire_4175, wire_13651, wire_6867, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6722, wire_4689, wire_4175, wire_6375, wire_6374, wire_4175, wire_6465, wire_6344, wire_4175, wire_13287, wire_13259, wire_13258, wire_13252, wire_13219, wire_13218, wire_13179, wire_13178, wire_6718, wire_4218, wire_13285, wire_13257, wire_13256, wire_13217, wire_13216, wire_13177, wire_13176, wire_13140, wire_6716, wire_4218, wire_13283, wire_13255, wire_13254, wire_13215, wire_13214, wire_13175, wire_13174, wire_13148, wire_6714, wire_4218, wire_13281, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_13156, wire_6712, wire_4178, wire_13279, wire_13249, wire_13248, wire_13209, wire_13208, wire_13169, wire_13168, wire_13164, wire_6710, wire_4178, wire_13277, wire_13247, wire_13246, wire_13207, wire_13206, wire_13172, wire_13167, wire_13166, wire_6708, wire_4178, wire_13275, wire_13243, wire_13242, wire_13203, wire_13202, wire_13180, wire_13163, wire_13162, wire_6706, wire_4222, wire_4178, wire_13273, wire_13241, wire_13240, wire_13201, wire_13200, wire_13188, wire_13161, wire_13160, wire_6704, wire_4222, wire_4178, wire_13271, wire_13239, wire_13238, wire_13199, wire_13198, wire_13196, wire_13159, wire_13158, wire_6702, wire_4222, wire_4178, wire_13269, wire_13235, wire_13234, wire_13204, wire_13195, wire_13194, wire_13155, wire_13154, wire_6700, wire_4222, wire_4174, wire_13267, wire_13233, wire_13232, wire_13212, wire_13193, wire_13192, wire_13153, wire_13152, wire_6698, wire_4222, wire_4174, wire_13265, wire_13231, wire_13230, wire_13220, wire_13191, wire_13190, wire_13151, wire_13150, wire_6696, wire_4222, wire_4174, wire_13263, wire_13228, wire_13227, wire_13226, wire_13187, wire_13186, wire_13147, wire_13146, wire_6694, wire_4218, wire_4174, wire_13261, wire_13236, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_6692, wire_4218, wire_4174, wire_13289, wire_13244, wire_13223, wire_13222, wire_13183, wire_13182, wire_13143, wire_13142, wire_6690, wire_4218, wire_4174, wire_13653, wire_13649, wire_13648, wire_13636, wire_13609, wire_13608, wire_13569, wire_13568, wire_6869, wire_4218, wire_13655, wire_13647, wire_13646, wire_13628, wire_13607, wire_13606, wire_13567, wire_13566, wire_6867, wire_4218, wire_13657, wire_13643, wire_13642, wire_13620, wire_13603, wire_13602, wire_13563, wire_13562, wire_6865, wire_4218, wire_13659, wire_13641, wire_13640, wire_13612, wire_13601, wire_13600, wire_13561, wire_13560, wire_6863, wire_4178, wire_13661, wire_13639, wire_13638, wire_13604, wire_13599, wire_13598, wire_13559, wire_13558, wire_6861, wire_4178, wire_13663, wire_13635, wire_13634, wire_13596, wire_13595, wire_13594, wire_13555, wire_13554, wire_6859, wire_4178, wire_13665, wire_13633, wire_13632, wire_13593, wire_13592, wire_13588, wire_13553, wire_13552, wire_6857, wire_4222, wire_4178, wire_13667, wire_13631, wire_13630, wire_13591, wire_13590, wire_13580, wire_13551, wire_13550, wire_6855, wire_4222, wire_4178, wire_13669, wire_13627, wire_13626, wire_13587, wire_13586, wire_13572, wire_13547, wire_13546, wire_6853, wire_4222, wire_4178, wire_13671, wire_13625, wire_13624, wire_13585, wire_13584, wire_13564, wire_13545, wire_13544, wire_6851, wire_4222, wire_4174, wire_13673, wire_13623, wire_13622, wire_13583, wire_13582, wire_13556, wire_13543, wire_13542, wire_6849, wire_4222, wire_4174, wire_13675, wire_13619, wire_13618, wire_13579, wire_13578, wire_13548, wire_13539, wire_13538, wire_6847, wire_4222, wire_4174, wire_13677, wire_13617, wire_13616, wire_13577, wire_13576, wire_13540, wire_13537, wire_13536, wire_6845, wire_4218, wire_4174, wire_13679, wire_13615, wire_13614, wire_13575, wire_13574, wire_13535, wire_13534, wire_13532, wire_6843, wire_4218, wire_4174, wire_13651, wire_13644, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_6841, wire_4218, wire_4174};
    // CHNAXY TOTAL: 621
    assign wire_6721 = lut_tile_1_8_chanxy_out[0];
    assign wire_6723 = lut_tile_1_8_chanxy_out[1];
    assign wire_6725 = lut_tile_1_8_chanxy_out[2];
    assign wire_6727 = lut_tile_1_8_chanxy_out[3];
    assign wire_6729 = lut_tile_1_8_chanxy_out[4];
    assign wire_6731 = lut_tile_1_8_chanxy_out[5];
    assign wire_6733 = lut_tile_1_8_chanxy_out[6];
    assign wire_6735 = lut_tile_1_8_chanxy_out[7];
    assign wire_6737 = lut_tile_1_8_chanxy_out[8];
    assign wire_6739 = lut_tile_1_8_chanxy_out[9];
    assign wire_6741 = lut_tile_1_8_chanxy_out[10];
    assign wire_6743 = lut_tile_1_8_chanxy_out[11];
    assign wire_6745 = lut_tile_1_8_chanxy_out[12];
    assign wire_6747 = lut_tile_1_8_chanxy_out[13];
    assign wire_6749 = lut_tile_1_8_chanxy_out[14];
    assign wire_6810 = lut_tile_1_8_chanxy_out[15];
    assign wire_6812 = lut_tile_1_8_chanxy_out[16];
    assign wire_6814 = lut_tile_1_8_chanxy_out[17];
    assign wire_6816 = lut_tile_1_8_chanxy_out[18];
    assign wire_6818 = lut_tile_1_8_chanxy_out[19];
    assign wire_6820 = lut_tile_1_8_chanxy_out[20];
    assign wire_6822 = lut_tile_1_8_chanxy_out[21];
    assign wire_6824 = lut_tile_1_8_chanxy_out[22];
    assign wire_6826 = lut_tile_1_8_chanxy_out[23];
    assign wire_6828 = lut_tile_1_8_chanxy_out[24];
    assign wire_6830 = lut_tile_1_8_chanxy_out[25];
    assign wire_6832 = lut_tile_1_8_chanxy_out[26];
    assign wire_6834 = lut_tile_1_8_chanxy_out[27];
    assign wire_6836 = lut_tile_1_8_chanxy_out[28];
    assign wire_6838 = lut_tile_1_8_chanxy_out[29];
    assign wire_13530 = lut_tile_1_8_chanxy_out[30];
    assign wire_13532 = lut_tile_1_8_chanxy_out[31];
    assign wire_13533 = lut_tile_1_8_chanxy_out[32];
    assign wire_13534 = lut_tile_1_8_chanxy_out[33];
    assign wire_13536 = lut_tile_1_8_chanxy_out[34];
    assign wire_13538 = lut_tile_1_8_chanxy_out[35];
    assign wire_13540 = lut_tile_1_8_chanxy_out[36];
    assign wire_13541 = lut_tile_1_8_chanxy_out[37];
    assign wire_13542 = lut_tile_1_8_chanxy_out[38];
    assign wire_13544 = lut_tile_1_8_chanxy_out[39];
    assign wire_13546 = lut_tile_1_8_chanxy_out[40];
    assign wire_13548 = lut_tile_1_8_chanxy_out[41];
    assign wire_13549 = lut_tile_1_8_chanxy_out[42];
    assign wire_13550 = lut_tile_1_8_chanxy_out[43];
    assign wire_13552 = lut_tile_1_8_chanxy_out[44];
    assign wire_13554 = lut_tile_1_8_chanxy_out[45];
    assign wire_13556 = lut_tile_1_8_chanxy_out[46];
    assign wire_13557 = lut_tile_1_8_chanxy_out[47];
    assign wire_13558 = lut_tile_1_8_chanxy_out[48];
    assign wire_13560 = lut_tile_1_8_chanxy_out[49];
    assign wire_13562 = lut_tile_1_8_chanxy_out[50];
    assign wire_13564 = lut_tile_1_8_chanxy_out[51];
    assign wire_13565 = lut_tile_1_8_chanxy_out[52];
    assign wire_13566 = lut_tile_1_8_chanxy_out[53];
    assign wire_13568 = lut_tile_1_8_chanxy_out[54];
    assign wire_13570 = lut_tile_1_8_chanxy_out[55];
    assign wire_13572 = lut_tile_1_8_chanxy_out[56];
    assign wire_13573 = lut_tile_1_8_chanxy_out[57];
    assign wire_13574 = lut_tile_1_8_chanxy_out[58];
    assign wire_13576 = lut_tile_1_8_chanxy_out[59];
    assign wire_13578 = lut_tile_1_8_chanxy_out[60];
    assign wire_13580 = lut_tile_1_8_chanxy_out[61];
    assign wire_13581 = lut_tile_1_8_chanxy_out[62];
    assign wire_13582 = lut_tile_1_8_chanxy_out[63];
    assign wire_13584 = lut_tile_1_8_chanxy_out[64];
    assign wire_13586 = lut_tile_1_8_chanxy_out[65];
    assign wire_13588 = lut_tile_1_8_chanxy_out[66];
    assign wire_13589 = lut_tile_1_8_chanxy_out[67];
    assign wire_13590 = lut_tile_1_8_chanxy_out[68];
    assign wire_13592 = lut_tile_1_8_chanxy_out[69];
    assign wire_13594 = lut_tile_1_8_chanxy_out[70];
    assign wire_13596 = lut_tile_1_8_chanxy_out[71];
    assign wire_13597 = lut_tile_1_8_chanxy_out[72];
    assign wire_13598 = lut_tile_1_8_chanxy_out[73];
    assign wire_13600 = lut_tile_1_8_chanxy_out[74];
    assign wire_13602 = lut_tile_1_8_chanxy_out[75];
    assign wire_13604 = lut_tile_1_8_chanxy_out[76];
    assign wire_13605 = lut_tile_1_8_chanxy_out[77];
    assign wire_13606 = lut_tile_1_8_chanxy_out[78];
    assign wire_13608 = lut_tile_1_8_chanxy_out[79];
    assign wire_13610 = lut_tile_1_8_chanxy_out[80];
    assign wire_13612 = lut_tile_1_8_chanxy_out[81];
    assign wire_13613 = lut_tile_1_8_chanxy_out[82];
    assign wire_13614 = lut_tile_1_8_chanxy_out[83];
    assign wire_13616 = lut_tile_1_8_chanxy_out[84];
    assign wire_13618 = lut_tile_1_8_chanxy_out[85];
    assign wire_13620 = lut_tile_1_8_chanxy_out[86];
    assign wire_13621 = lut_tile_1_8_chanxy_out[87];
    assign wire_13622 = lut_tile_1_8_chanxy_out[88];
    assign wire_13624 = lut_tile_1_8_chanxy_out[89];
    assign wire_13626 = lut_tile_1_8_chanxy_out[90];
    assign wire_13628 = lut_tile_1_8_chanxy_out[91];
    assign wire_13629 = lut_tile_1_8_chanxy_out[92];
    assign wire_13630 = lut_tile_1_8_chanxy_out[93];
    assign wire_13632 = lut_tile_1_8_chanxy_out[94];
    assign wire_13634 = lut_tile_1_8_chanxy_out[95];
    assign wire_13636 = lut_tile_1_8_chanxy_out[96];
    assign wire_13637 = lut_tile_1_8_chanxy_out[97];
    assign wire_13638 = lut_tile_1_8_chanxy_out[98];
    assign wire_13640 = lut_tile_1_8_chanxy_out[99];
    assign wire_13642 = lut_tile_1_8_chanxy_out[100];
    assign wire_13644 = lut_tile_1_8_chanxy_out[101];
    assign wire_13645 = lut_tile_1_8_chanxy_out[102];
    assign wire_13646 = lut_tile_1_8_chanxy_out[103];
    assign wire_13648 = lut_tile_1_8_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_9_chanxy_in = {wire_6433, wire_6432, wire_14069, wire_6899, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6750, wire_5205, wire_6449, wire_6448, wire_6419, wire_6418, wire_6403, wire_6402, wire_6509, wire_6388, wire_14067, wire_6871, wire_6869, wire_6868, wire_6859, wire_6858, wire_6849, wire_6848, wire_6778, wire_5205, wire_6479, wire_6478, wire_6493, wire_6372, wire_6447, wire_6446, wire_6417, wire_6416, wire_14065, wire_6873, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6776, wire_5205, wire_6463, wire_6462, wire_6507, wire_6386, wire_6477, wire_6476, wire_6445, wire_6444, wire_14063, wire_6875, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6774, wire_4695, wire_6431, wire_6430, wire_6401, wire_6400, wire_6415, wire_6414, wire_6491, wire_6370, wire_14061, wire_6877, wire_6867, wire_6866, wire_6857, wire_6856, wire_6847, wire_6846, wire_6772, wire_4695, wire_6461, wire_6460, wire_6505, wire_6384, wire_6429, wire_6428, wire_6399, wire_6398, wire_14059, wire_6879, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6770, wire_4695, wire_6475, wire_6474, wire_6489, wire_6368, wire_6459, wire_6458, wire_6427, wire_6426, wire_14057, wire_6881, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6768, wire_5209, wire_4695, wire_6443, wire_6442, wire_6413, wire_6412, wire_6397, wire_6396, wire_6503, wire_6382, wire_14055, wire_6883, wire_6865, wire_6864, wire_6855, wire_6854, wire_6845, wire_6844, wire_6766, wire_5209, wire_4695, wire_6473, wire_6472, wire_6487, wire_6366, wire_6441, wire_6440, wire_6411, wire_6410, wire_14053, wire_6885, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6764, wire_5209, wire_4695, wire_6457, wire_6456, wire_6501, wire_6380, wire_6471, wire_6470, wire_6439, wire_6438, wire_5209, wire_14051, wire_6887, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6762, wire_5209, wire_4691, wire_6425, wire_6424, wire_5209, wire_6395, wire_6394, wire_5209, wire_6409, wire_6408, wire_5209, wire_6485, wire_6364, wire_5209, wire_14049, wire_6889, wire_6863, wire_6862, wire_6853, wire_6852, wire_6843, wire_6842, wire_6760, wire_5209, wire_4691, wire_6455, wire_6454, wire_5209, wire_6499, wire_6378, wire_5205, wire_6423, wire_6422, wire_5205, wire_6393, wire_6392, wire_5205, wire_14047, wire_6891, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6758, wire_5209, wire_4691, wire_6469, wire_6468, wire_5205, wire_6483, wire_6362, wire_5205, wire_6453, wire_6452, wire_5205, wire_6421, wire_6420, wire_4695, wire_14045, wire_6893, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6756, wire_5205, wire_4691, wire_6437, wire_6436, wire_4695, wire_6407, wire_6406, wire_4695, wire_6391, wire_6390, wire_4695, wire_6497, wire_6376, wire_4695, wire_14043, wire_6895, wire_6861, wire_6860, wire_6851, wire_6850, wire_6841, wire_6840, wire_6754, wire_5205, wire_4691, wire_6467, wire_6466, wire_4695, wire_6481, wire_6360, wire_4691, wire_6435, wire_6434, wire_4691, wire_6405, wire_6404, wire_4691, wire_14041, wire_6897, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6752, wire_5205, wire_4691, wire_6451, wire_6450, wire_4691, wire_6495, wire_6374, wire_4691, wire_6465, wire_6464, wire_4691, wire_13677, wire_13649, wire_13648, wire_13644, wire_13609, wire_13608, wire_13569, wire_13568, wire_6748, wire_4734, wire_13675, wire_13647, wire_13646, wire_13607, wire_13606, wire_13567, wire_13566, wire_13532, wire_6746, wire_4734, wire_13673, wire_13643, wire_13642, wire_13603, wire_13602, wire_13563, wire_13562, wire_13540, wire_6744, wire_4734, wire_13671, wire_13641, wire_13640, wire_13601, wire_13600, wire_13561, wire_13560, wire_13548, wire_6742, wire_4694, wire_13669, wire_13639, wire_13638, wire_13599, wire_13598, wire_13559, wire_13558, wire_13556, wire_6740, wire_4694, wire_13667, wire_13635, wire_13634, wire_13595, wire_13594, wire_13564, wire_13555, wire_13554, wire_6738, wire_4694, wire_13665, wire_13633, wire_13632, wire_13593, wire_13592, wire_13572, wire_13553, wire_13552, wire_6736, wire_4738, wire_4694, wire_13663, wire_13631, wire_13630, wire_13591, wire_13590, wire_13580, wire_13551, wire_13550, wire_6734, wire_4738, wire_4694, wire_13661, wire_13627, wire_13626, wire_13588, wire_13587, wire_13586, wire_13547, wire_13546, wire_6732, wire_4738, wire_4694, wire_13659, wire_13625, wire_13624, wire_13596, wire_13585, wire_13584, wire_13545, wire_13544, wire_6730, wire_4738, wire_4690, wire_13657, wire_13623, wire_13622, wire_13604, wire_13583, wire_13582, wire_13543, wire_13542, wire_6728, wire_4738, wire_4690, wire_13655, wire_13619, wire_13618, wire_13612, wire_13579, wire_13578, wire_13539, wire_13538, wire_6726, wire_4738, wire_4690, wire_13653, wire_13620, wire_13617, wire_13616, wire_13577, wire_13576, wire_13537, wire_13536, wire_6724, wire_4734, wire_4690, wire_13651, wire_13628, wire_13615, wire_13614, wire_13575, wire_13574, wire_13535, wire_13534, wire_6722, wire_4734, wire_4690, wire_13679, wire_13636, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_6720, wire_4734, wire_4690, wire_14043, wire_14039, wire_14038, wire_14028, wire_13999, wire_13998, wire_13959, wire_13958, wire_6899, wire_4734, wire_14045, wire_14035, wire_14034, wire_14020, wire_13995, wire_13994, wire_13955, wire_13954, wire_6897, wire_4734, wire_14047, wire_14033, wire_14032, wire_14012, wire_13993, wire_13992, wire_13953, wire_13952, wire_6895, wire_4734, wire_14049, wire_14031, wire_14030, wire_14004, wire_13991, wire_13990, wire_13951, wire_13950, wire_6893, wire_4694, wire_14051, wire_14027, wire_14026, wire_13996, wire_13987, wire_13986, wire_13947, wire_13946, wire_6891, wire_4694, wire_14053, wire_14025, wire_14024, wire_13988, wire_13985, wire_13984, wire_13945, wire_13944, wire_6889, wire_4694, wire_14055, wire_14023, wire_14022, wire_13983, wire_13982, wire_13980, wire_13943, wire_13942, wire_6887, wire_4738, wire_4694, wire_14057, wire_14019, wire_14018, wire_13979, wire_13978, wire_13972, wire_13939, wire_13938, wire_6885, wire_4738, wire_4694, wire_14059, wire_14017, wire_14016, wire_13977, wire_13976, wire_13964, wire_13937, wire_13936, wire_6883, wire_4738, wire_4694, wire_14061, wire_14015, wire_14014, wire_13975, wire_13974, wire_13956, wire_13935, wire_13934, wire_6881, wire_4738, wire_4690, wire_14063, wire_14011, wire_14010, wire_13971, wire_13970, wire_13948, wire_13931, wire_13930, wire_6879, wire_4738, wire_4690, wire_14065, wire_14009, wire_14008, wire_13969, wire_13968, wire_13940, wire_13929, wire_13928, wire_6877, wire_4738, wire_4690, wire_14067, wire_14007, wire_14006, wire_13967, wire_13966, wire_13932, wire_13927, wire_13926, wire_6875, wire_4734, wire_4690, wire_14069, wire_14003, wire_14002, wire_13963, wire_13962, wire_13924, wire_13923, wire_13922, wire_6873, wire_4734, wire_4690, wire_14041, wire_14036, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_6871, wire_4734, wire_4690};
    // CHNAXY TOTAL: 621
    assign wire_6751 = lut_tile_1_9_chanxy_out[0];
    assign wire_6753 = lut_tile_1_9_chanxy_out[1];
    assign wire_6755 = lut_tile_1_9_chanxy_out[2];
    assign wire_6757 = lut_tile_1_9_chanxy_out[3];
    assign wire_6759 = lut_tile_1_9_chanxy_out[4];
    assign wire_6761 = lut_tile_1_9_chanxy_out[5];
    assign wire_6763 = lut_tile_1_9_chanxy_out[6];
    assign wire_6765 = lut_tile_1_9_chanxy_out[7];
    assign wire_6767 = lut_tile_1_9_chanxy_out[8];
    assign wire_6769 = lut_tile_1_9_chanxy_out[9];
    assign wire_6771 = lut_tile_1_9_chanxy_out[10];
    assign wire_6773 = lut_tile_1_9_chanxy_out[11];
    assign wire_6775 = lut_tile_1_9_chanxy_out[12];
    assign wire_6777 = lut_tile_1_9_chanxy_out[13];
    assign wire_6779 = lut_tile_1_9_chanxy_out[14];
    assign wire_6840 = lut_tile_1_9_chanxy_out[15];
    assign wire_6842 = lut_tile_1_9_chanxy_out[16];
    assign wire_6844 = lut_tile_1_9_chanxy_out[17];
    assign wire_6846 = lut_tile_1_9_chanxy_out[18];
    assign wire_6848 = lut_tile_1_9_chanxy_out[19];
    assign wire_6850 = lut_tile_1_9_chanxy_out[20];
    assign wire_6852 = lut_tile_1_9_chanxy_out[21];
    assign wire_6854 = lut_tile_1_9_chanxy_out[22];
    assign wire_6856 = lut_tile_1_9_chanxy_out[23];
    assign wire_6858 = lut_tile_1_9_chanxy_out[24];
    assign wire_6860 = lut_tile_1_9_chanxy_out[25];
    assign wire_6862 = lut_tile_1_9_chanxy_out[26];
    assign wire_6864 = lut_tile_1_9_chanxy_out[27];
    assign wire_6866 = lut_tile_1_9_chanxy_out[28];
    assign wire_6868 = lut_tile_1_9_chanxy_out[29];
    assign wire_13920 = lut_tile_1_9_chanxy_out[30];
    assign wire_13922 = lut_tile_1_9_chanxy_out[31];
    assign wire_13924 = lut_tile_1_9_chanxy_out[32];
    assign wire_13925 = lut_tile_1_9_chanxy_out[33];
    assign wire_13926 = lut_tile_1_9_chanxy_out[34];
    assign wire_13928 = lut_tile_1_9_chanxy_out[35];
    assign wire_13930 = lut_tile_1_9_chanxy_out[36];
    assign wire_13932 = lut_tile_1_9_chanxy_out[37];
    assign wire_13933 = lut_tile_1_9_chanxy_out[38];
    assign wire_13934 = lut_tile_1_9_chanxy_out[39];
    assign wire_13936 = lut_tile_1_9_chanxy_out[40];
    assign wire_13938 = lut_tile_1_9_chanxy_out[41];
    assign wire_13940 = lut_tile_1_9_chanxy_out[42];
    assign wire_13941 = lut_tile_1_9_chanxy_out[43];
    assign wire_13942 = lut_tile_1_9_chanxy_out[44];
    assign wire_13944 = lut_tile_1_9_chanxy_out[45];
    assign wire_13946 = lut_tile_1_9_chanxy_out[46];
    assign wire_13948 = lut_tile_1_9_chanxy_out[47];
    assign wire_13949 = lut_tile_1_9_chanxy_out[48];
    assign wire_13950 = lut_tile_1_9_chanxy_out[49];
    assign wire_13952 = lut_tile_1_9_chanxy_out[50];
    assign wire_13954 = lut_tile_1_9_chanxy_out[51];
    assign wire_13956 = lut_tile_1_9_chanxy_out[52];
    assign wire_13957 = lut_tile_1_9_chanxy_out[53];
    assign wire_13958 = lut_tile_1_9_chanxy_out[54];
    assign wire_13960 = lut_tile_1_9_chanxy_out[55];
    assign wire_13962 = lut_tile_1_9_chanxy_out[56];
    assign wire_13964 = lut_tile_1_9_chanxy_out[57];
    assign wire_13965 = lut_tile_1_9_chanxy_out[58];
    assign wire_13966 = lut_tile_1_9_chanxy_out[59];
    assign wire_13968 = lut_tile_1_9_chanxy_out[60];
    assign wire_13970 = lut_tile_1_9_chanxy_out[61];
    assign wire_13972 = lut_tile_1_9_chanxy_out[62];
    assign wire_13973 = lut_tile_1_9_chanxy_out[63];
    assign wire_13974 = lut_tile_1_9_chanxy_out[64];
    assign wire_13976 = lut_tile_1_9_chanxy_out[65];
    assign wire_13978 = lut_tile_1_9_chanxy_out[66];
    assign wire_13980 = lut_tile_1_9_chanxy_out[67];
    assign wire_13981 = lut_tile_1_9_chanxy_out[68];
    assign wire_13982 = lut_tile_1_9_chanxy_out[69];
    assign wire_13984 = lut_tile_1_9_chanxy_out[70];
    assign wire_13986 = lut_tile_1_9_chanxy_out[71];
    assign wire_13988 = lut_tile_1_9_chanxy_out[72];
    assign wire_13989 = lut_tile_1_9_chanxy_out[73];
    assign wire_13990 = lut_tile_1_9_chanxy_out[74];
    assign wire_13992 = lut_tile_1_9_chanxy_out[75];
    assign wire_13994 = lut_tile_1_9_chanxy_out[76];
    assign wire_13996 = lut_tile_1_9_chanxy_out[77];
    assign wire_13997 = lut_tile_1_9_chanxy_out[78];
    assign wire_13998 = lut_tile_1_9_chanxy_out[79];
    assign wire_14000 = lut_tile_1_9_chanxy_out[80];
    assign wire_14002 = lut_tile_1_9_chanxy_out[81];
    assign wire_14004 = lut_tile_1_9_chanxy_out[82];
    assign wire_14005 = lut_tile_1_9_chanxy_out[83];
    assign wire_14006 = lut_tile_1_9_chanxy_out[84];
    assign wire_14008 = lut_tile_1_9_chanxy_out[85];
    assign wire_14010 = lut_tile_1_9_chanxy_out[86];
    assign wire_14012 = lut_tile_1_9_chanxy_out[87];
    assign wire_14013 = lut_tile_1_9_chanxy_out[88];
    assign wire_14014 = lut_tile_1_9_chanxy_out[89];
    assign wire_14016 = lut_tile_1_9_chanxy_out[90];
    assign wire_14018 = lut_tile_1_9_chanxy_out[91];
    assign wire_14020 = lut_tile_1_9_chanxy_out[92];
    assign wire_14021 = lut_tile_1_9_chanxy_out[93];
    assign wire_14022 = lut_tile_1_9_chanxy_out[94];
    assign wire_14024 = lut_tile_1_9_chanxy_out[95];
    assign wire_14026 = lut_tile_1_9_chanxy_out[96];
    assign wire_14028 = lut_tile_1_9_chanxy_out[97];
    assign wire_14029 = lut_tile_1_9_chanxy_out[98];
    assign wire_14030 = lut_tile_1_9_chanxy_out[99];
    assign wire_14032 = lut_tile_1_9_chanxy_out[100];
    assign wire_14034 = lut_tile_1_9_chanxy_out[101];
    assign wire_14036 = lut_tile_1_9_chanxy_out[102];
    assign wire_14037 = lut_tile_1_9_chanxy_out[103];
    assign wire_14038 = lut_tile_1_9_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_1_10_chanxy_in = {wire_14459, wire_6876, wire_6854, wire_6832, wire_6808, wire_5686, wire_5680, wire_5671, wire_5665, wire_6480, wire_5686, wire_6390, wire_5686, wire_6420, wire_5686, wire_6452, wire_5686, wire_14457, wire_6898, wire_6846, wire_6824, wire_6800, wire_5686, wire_5680, wire_5671, wire_5665, wire_6482, wire_5686, wire_6392, wire_5686, wire_6422, wire_5683, wire_6454, wire_5683, wire_14455, wire_6890, wire_6868, wire_6816, wire_6792, wire_5686, wire_5680, wire_5671, wire_5665, wire_6484, wire_5683, wire_6394, wire_5683, wire_6424, wire_5683, wire_6456, wire_5683, wire_14453, wire_6882, wire_6860, wire_6838, wire_6784, wire_5686, wire_5677, wire_5671, wire_5211, wire_6486, wire_5680, wire_6396, wire_5680, wire_6426, wire_5680, wire_6458, wire_5680, wire_14451, wire_6874, wire_6852, wire_6830, wire_6806, wire_5686, wire_5677, wire_5671, wire_5211, wire_6488, wire_5680, wire_6398, wire_5680, wire_6428, wire_5677, wire_6460, wire_5677, wire_14449, wire_6896, wire_6844, wire_6822, wire_6798, wire_5686, wire_5677, wire_5671, wire_5211, wire_6490, wire_5677, wire_6400, wire_5677, wire_6430, wire_5677, wire_6462, wire_5677, wire_14447, wire_6888, wire_6866, wire_6814, wire_6790, wire_5683, wire_5677, wire_5668, wire_5211, wire_6492, wire_5674, wire_6402, wire_5674, wire_6432, wire_5674, wire_6464, wire_5674, wire_14445, wire_6880, wire_6858, wire_6836, wire_6782, wire_5683, wire_5677, wire_5668, wire_5211, wire_6494, wire_5674, wire_6404, wire_5674, wire_6434, wire_5671, wire_6466, wire_5671, wire_14443, wire_6872, wire_6850, wire_6828, wire_6804, wire_5683, wire_5677, wire_5668, wire_5211, wire_6496, wire_5671, wire_6406, wire_5671, wire_6436, wire_5671, wire_6468, wire_5671, wire_14441, wire_6894, wire_6842, wire_6820, wire_6796, wire_5683, wire_5674, wire_5668, wire_5207, wire_6498, wire_5668, wire_6408, wire_5668, wire_6438, wire_5668, wire_6470, wire_5668, wire_14439, wire_6886, wire_6864, wire_6812, wire_6788, wire_5683, wire_5674, wire_5668, wire_5207, wire_6500, wire_5668, wire_6410, wire_5668, wire_6440, wire_5665, wire_6472, wire_5665, wire_14437, wire_6878, wire_6856, wire_6834, wire_6780, wire_5683, wire_5674, wire_5668, wire_5207, wire_6502, wire_5665, wire_6412, wire_5665, wire_6442, wire_5665, wire_6474, wire_5665, wire_14435, wire_6870, wire_6848, wire_6826, wire_6802, wire_5680, wire_5674, wire_5665, wire_5207, wire_6504, wire_5211, wire_6414, wire_5211, wire_6444, wire_5211, wire_6476, wire_5211, wire_14433, wire_6892, wire_6840, wire_6818, wire_6794, wire_5680, wire_5674, wire_5665, wire_5207, wire_6506, wire_5211, wire_6416, wire_5211, wire_6446, wire_5207, wire_6478, wire_5207, wire_14431, wire_6884, wire_6862, wire_6810, wire_6786, wire_5680, wire_5674, wire_5665, wire_5207, wire_6508, wire_5207, wire_6418, wire_5207, wire_6448, wire_5207, wire_6450, wire_5207, wire_14427, wire_14426, wire_14067, wire_14039, wire_14038, wire_14036, wire_13999, wire_13998, wire_13959, wire_13958, wire_6778, wire_5250, wire_14363, wire_14362, wire_14065, wire_14035, wire_14034, wire_13995, wire_13994, wire_13955, wire_13954, wire_13924, wire_6776, wire_5250, wire_14417, wire_14416, wire_14063, wire_14033, wire_14032, wire_13993, wire_13992, wire_13953, wire_13952, wire_13932, wire_6774, wire_5250, wire_14355, wire_14354, wire_14061, wire_14031, wire_14030, wire_13991, wire_13990, wire_13951, wire_13950, wire_13940, wire_6772, wire_5210, wire_14411, wire_14410, wire_14059, wire_14027, wire_14026, wire_13987, wire_13986, wire_13948, wire_13947, wire_13946, wire_6770, wire_5210, wire_14345, wire_14344, wire_14057, wire_14025, wire_14024, wire_13985, wire_13984, wire_13956, wire_13945, wire_13944, wire_6768, wire_5210, wire_14403, wire_14402, wire_14055, wire_14023, wire_14022, wire_13983, wire_13982, wire_13964, wire_13943, wire_13942, wire_6766, wire_5254, wire_5210, wire_14339, wire_14338, wire_14053, wire_14019, wire_14018, wire_13979, wire_13978, wire_13972, wire_13939, wire_13938, wire_6764, wire_5254, wire_5210, wire_14393, wire_14392, wire_14051, wire_14017, wire_14016, wire_13980, wire_13977, wire_13976, wire_13937, wire_13936, wire_6762, wire_5254, wire_5210, wire_14331, wire_14330, wire_5254, wire_14049, wire_14015, wire_14014, wire_13988, wire_13975, wire_13974, wire_13935, wire_13934, wire_6760, wire_5254, wire_5206, wire_14387, wire_14386, wire_5254, wire_14047, wire_14011, wire_14010, wire_13996, wire_13971, wire_13970, wire_13931, wire_13930, wire_6758, wire_5254, wire_5206, wire_14321, wire_14320, wire_5250, wire_14045, wire_14009, wire_14008, wire_14004, wire_13969, wire_13968, wire_13929, wire_13928, wire_6756, wire_5254, wire_5206, wire_14379, wire_14378, wire_5210, wire_14043, wire_14012, wire_14007, wire_14006, wire_13967, wire_13966, wire_13927, wire_13926, wire_6754, wire_5250, wire_5206, wire_14315, wire_14314, wire_5210, wire_14041, wire_14020, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_6752, wire_5250, wire_5206, wire_14369, wire_14368, wire_5206, wire_14069, wire_14028, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_6750, wire_5250, wire_5206, wire_14443, wire_14364, wire_14457, wire_14420, wire_14415, wire_14414, wire_14455, wire_14412, wire_14439, wire_14348, wire_14343, wire_14342, wire_14437, wire_14340, wire_14451, wire_14396, wire_14391, wire_14390, wire_14449, wire_14388, wire_5254, wire_14433, wire_14324, wire_5250, wire_14319, wire_14318, wire_5250, wire_14431, wire_14316, wire_5210, wire_14445, wire_14372, wire_5206, wire_14367, wire_14366, wire_5206, wire_14425, wire_14424, wire_14419, wire_14418, wire_14359, wire_14358, wire_14353, wire_14352, wire_14347, wire_14346, wire_14407, wire_14406, wire_14401, wire_14400, wire_14395, wire_14394, wire_14335, wire_14334, wire_14329, wire_14328, wire_5254, wire_14323, wire_14322, wire_5250, wire_14383, wire_14382, wire_5250, wire_14377, wire_14376, wire_5210, wire_14371, wire_14370, wire_5206, wire_14311, wire_14310, wire_5206, wire_14459, wire_14428, wire_14423, wire_14422, wire_14361, wire_14360, wire_14441, wire_14356, wire_14351, wire_14350, wire_14409, wire_14408, wire_14453, wire_14404, wire_14399, wire_14398, wire_14337, wire_14336, wire_14435, wire_14332, wire_5254, wire_14327, wire_14326, wire_5254, wire_14385, wire_14384, wire_5250, wire_14447, wire_14380, wire_5210, wire_14375, wire_14374, wire_5210, wire_14313, wire_14312, wire_5206};
    // CHNAXY TOTAL: 558
    assign wire_6781 = lut_tile_1_10_chanxy_out[0];
    assign wire_6783 = lut_tile_1_10_chanxy_out[1];
    assign wire_6785 = lut_tile_1_10_chanxy_out[2];
    assign wire_6787 = lut_tile_1_10_chanxy_out[3];
    assign wire_6789 = lut_tile_1_10_chanxy_out[4];
    assign wire_6791 = lut_tile_1_10_chanxy_out[5];
    assign wire_6793 = lut_tile_1_10_chanxy_out[6];
    assign wire_6795 = lut_tile_1_10_chanxy_out[7];
    assign wire_6797 = lut_tile_1_10_chanxy_out[8];
    assign wire_6799 = lut_tile_1_10_chanxy_out[9];
    assign wire_6801 = lut_tile_1_10_chanxy_out[10];
    assign wire_6803 = lut_tile_1_10_chanxy_out[11];
    assign wire_6805 = lut_tile_1_10_chanxy_out[12];
    assign wire_6807 = lut_tile_1_10_chanxy_out[13];
    assign wire_6809 = lut_tile_1_10_chanxy_out[14];
    assign wire_6811 = lut_tile_1_10_chanxy_out[15];
    assign wire_6813 = lut_tile_1_10_chanxy_out[16];
    assign wire_6815 = lut_tile_1_10_chanxy_out[17];
    assign wire_6817 = lut_tile_1_10_chanxy_out[18];
    assign wire_6819 = lut_tile_1_10_chanxy_out[19];
    assign wire_6821 = lut_tile_1_10_chanxy_out[20];
    assign wire_6823 = lut_tile_1_10_chanxy_out[21];
    assign wire_6825 = lut_tile_1_10_chanxy_out[22];
    assign wire_6827 = lut_tile_1_10_chanxy_out[23];
    assign wire_6829 = lut_tile_1_10_chanxy_out[24];
    assign wire_6831 = lut_tile_1_10_chanxy_out[25];
    assign wire_6833 = lut_tile_1_10_chanxy_out[26];
    assign wire_6835 = lut_tile_1_10_chanxy_out[27];
    assign wire_6837 = lut_tile_1_10_chanxy_out[28];
    assign wire_6839 = lut_tile_1_10_chanxy_out[29];
    assign wire_6841 = lut_tile_1_10_chanxy_out[30];
    assign wire_6843 = lut_tile_1_10_chanxy_out[31];
    assign wire_6845 = lut_tile_1_10_chanxy_out[32];
    assign wire_6847 = lut_tile_1_10_chanxy_out[33];
    assign wire_6849 = lut_tile_1_10_chanxy_out[34];
    assign wire_6851 = lut_tile_1_10_chanxy_out[35];
    assign wire_6853 = lut_tile_1_10_chanxy_out[36];
    assign wire_6855 = lut_tile_1_10_chanxy_out[37];
    assign wire_6857 = lut_tile_1_10_chanxy_out[38];
    assign wire_6859 = lut_tile_1_10_chanxy_out[39];
    assign wire_6861 = lut_tile_1_10_chanxy_out[40];
    assign wire_6863 = lut_tile_1_10_chanxy_out[41];
    assign wire_6865 = lut_tile_1_10_chanxy_out[42];
    assign wire_6867 = lut_tile_1_10_chanxy_out[43];
    assign wire_6869 = lut_tile_1_10_chanxy_out[44];
    assign wire_6870 = lut_tile_1_10_chanxy_out[45];
    assign wire_6871 = lut_tile_1_10_chanxy_out[46];
    assign wire_6872 = lut_tile_1_10_chanxy_out[47];
    assign wire_6873 = lut_tile_1_10_chanxy_out[48];
    assign wire_6874 = lut_tile_1_10_chanxy_out[49];
    assign wire_6875 = lut_tile_1_10_chanxy_out[50];
    assign wire_6876 = lut_tile_1_10_chanxy_out[51];
    assign wire_6877 = lut_tile_1_10_chanxy_out[52];
    assign wire_6878 = lut_tile_1_10_chanxy_out[53];
    assign wire_6879 = lut_tile_1_10_chanxy_out[54];
    assign wire_6880 = lut_tile_1_10_chanxy_out[55];
    assign wire_6881 = lut_tile_1_10_chanxy_out[56];
    assign wire_6882 = lut_tile_1_10_chanxy_out[57];
    assign wire_6883 = lut_tile_1_10_chanxy_out[58];
    assign wire_6884 = lut_tile_1_10_chanxy_out[59];
    assign wire_6885 = lut_tile_1_10_chanxy_out[60];
    assign wire_6886 = lut_tile_1_10_chanxy_out[61];
    assign wire_6887 = lut_tile_1_10_chanxy_out[62];
    assign wire_6888 = lut_tile_1_10_chanxy_out[63];
    assign wire_6889 = lut_tile_1_10_chanxy_out[64];
    assign wire_6890 = lut_tile_1_10_chanxy_out[65];
    assign wire_6891 = lut_tile_1_10_chanxy_out[66];
    assign wire_6892 = lut_tile_1_10_chanxy_out[67];
    assign wire_6893 = lut_tile_1_10_chanxy_out[68];
    assign wire_6894 = lut_tile_1_10_chanxy_out[69];
    assign wire_6895 = lut_tile_1_10_chanxy_out[70];
    assign wire_6896 = lut_tile_1_10_chanxy_out[71];
    assign wire_6897 = lut_tile_1_10_chanxy_out[72];
    assign wire_6898 = lut_tile_1_10_chanxy_out[73];
    assign wire_6899 = lut_tile_1_10_chanxy_out[74];
    assign wire_14310 = lut_tile_1_10_chanxy_out[75];
    assign wire_14312 = lut_tile_1_10_chanxy_out[76];
    assign wire_14314 = lut_tile_1_10_chanxy_out[77];
    assign wire_14316 = lut_tile_1_10_chanxy_out[78];
    assign wire_14317 = lut_tile_1_10_chanxy_out[79];
    assign wire_14318 = lut_tile_1_10_chanxy_out[80];
    assign wire_14320 = lut_tile_1_10_chanxy_out[81];
    assign wire_14322 = lut_tile_1_10_chanxy_out[82];
    assign wire_14324 = lut_tile_1_10_chanxy_out[83];
    assign wire_14325 = lut_tile_1_10_chanxy_out[84];
    assign wire_14326 = lut_tile_1_10_chanxy_out[85];
    assign wire_14328 = lut_tile_1_10_chanxy_out[86];
    assign wire_14330 = lut_tile_1_10_chanxy_out[87];
    assign wire_14332 = lut_tile_1_10_chanxy_out[88];
    assign wire_14333 = lut_tile_1_10_chanxy_out[89];
    assign wire_14334 = lut_tile_1_10_chanxy_out[90];
    assign wire_14336 = lut_tile_1_10_chanxy_out[91];
    assign wire_14338 = lut_tile_1_10_chanxy_out[92];
    assign wire_14340 = lut_tile_1_10_chanxy_out[93];
    assign wire_14341 = lut_tile_1_10_chanxy_out[94];
    assign wire_14342 = lut_tile_1_10_chanxy_out[95];
    assign wire_14344 = lut_tile_1_10_chanxy_out[96];
    assign wire_14346 = lut_tile_1_10_chanxy_out[97];
    assign wire_14348 = lut_tile_1_10_chanxy_out[98];
    assign wire_14349 = lut_tile_1_10_chanxy_out[99];
    assign wire_14350 = lut_tile_1_10_chanxy_out[100];
    assign wire_14352 = lut_tile_1_10_chanxy_out[101];
    assign wire_14354 = lut_tile_1_10_chanxy_out[102];
    assign wire_14356 = lut_tile_1_10_chanxy_out[103];
    assign wire_14357 = lut_tile_1_10_chanxy_out[104];
    assign wire_14358 = lut_tile_1_10_chanxy_out[105];
    assign wire_14360 = lut_tile_1_10_chanxy_out[106];
    assign wire_14362 = lut_tile_1_10_chanxy_out[107];
    assign wire_14364 = lut_tile_1_10_chanxy_out[108];
    assign wire_14365 = lut_tile_1_10_chanxy_out[109];
    assign wire_14366 = lut_tile_1_10_chanxy_out[110];
    assign wire_14368 = lut_tile_1_10_chanxy_out[111];
    assign wire_14370 = lut_tile_1_10_chanxy_out[112];
    assign wire_14372 = lut_tile_1_10_chanxy_out[113];
    assign wire_14373 = lut_tile_1_10_chanxy_out[114];
    assign wire_14374 = lut_tile_1_10_chanxy_out[115];
    assign wire_14376 = lut_tile_1_10_chanxy_out[116];
    assign wire_14378 = lut_tile_1_10_chanxy_out[117];
    assign wire_14380 = lut_tile_1_10_chanxy_out[118];
    assign wire_14381 = lut_tile_1_10_chanxy_out[119];
    assign wire_14382 = lut_tile_1_10_chanxy_out[120];
    assign wire_14384 = lut_tile_1_10_chanxy_out[121];
    assign wire_14386 = lut_tile_1_10_chanxy_out[122];
    assign wire_14388 = lut_tile_1_10_chanxy_out[123];
    assign wire_14389 = lut_tile_1_10_chanxy_out[124];
    assign wire_14390 = lut_tile_1_10_chanxy_out[125];
    assign wire_14392 = lut_tile_1_10_chanxy_out[126];
    assign wire_14394 = lut_tile_1_10_chanxy_out[127];
    assign wire_14396 = lut_tile_1_10_chanxy_out[128];
    assign wire_14397 = lut_tile_1_10_chanxy_out[129];
    assign wire_14398 = lut_tile_1_10_chanxy_out[130];
    assign wire_14400 = lut_tile_1_10_chanxy_out[131];
    assign wire_14402 = lut_tile_1_10_chanxy_out[132];
    assign wire_14404 = lut_tile_1_10_chanxy_out[133];
    assign wire_14405 = lut_tile_1_10_chanxy_out[134];
    assign wire_14406 = lut_tile_1_10_chanxy_out[135];
    assign wire_14408 = lut_tile_1_10_chanxy_out[136];
    assign wire_14410 = lut_tile_1_10_chanxy_out[137];
    assign wire_14412 = lut_tile_1_10_chanxy_out[138];
    assign wire_14413 = lut_tile_1_10_chanxy_out[139];
    assign wire_14414 = lut_tile_1_10_chanxy_out[140];
    assign wire_14416 = lut_tile_1_10_chanxy_out[141];
    assign wire_14418 = lut_tile_1_10_chanxy_out[142];
    assign wire_14420 = lut_tile_1_10_chanxy_out[143];
    assign wire_14421 = lut_tile_1_10_chanxy_out[144];
    assign wire_14422 = lut_tile_1_10_chanxy_out[145];
    assign wire_14424 = lut_tile_1_10_chanxy_out[146];
    assign wire_14426 = lut_tile_1_10_chanxy_out[147];
    assign wire_14428 = lut_tile_1_10_chanxy_out[148];
    assign wire_14429 = lut_tile_1_10_chanxy_out[149];
   // CHANXY OUT
    assign lut_tile_2_1_chanxy_in = {wire_10916, wire_6631, wire_6629, wire_6628, wire_6589, wire_6588, wire_6549, wire_6548, wire_6522, wire_1119, wire_10908, wire_6659, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_6530, wire_1119, wire_10900, wire_6657, wire_6623, wire_6622, wire_6583, wire_6582, wire_6543, wire_6542, wire_6538, wire_1119, wire_10892, wire_6655, wire_6621, wire_6620, wire_6581, wire_6580, wire_6546, wire_6541, wire_6540, wire_609, wire_10884, wire_6653, wire_6617, wire_6616, wire_6577, wire_6576, wire_6554, wire_6537, wire_6536, wire_609, wire_10876, wire_6651, wire_6615, wire_6614, wire_6575, wire_6574, wire_6562, wire_6535, wire_6534, wire_609, wire_10868, wire_6649, wire_6613, wire_6612, wire_6573, wire_6572, wire_6570, wire_6533, wire_6532, wire_1123, wire_609, wire_10860, wire_6647, wire_6609, wire_6608, wire_6578, wire_6569, wire_6568, wire_6529, wire_6528, wire_1123, wire_609, wire_10852, wire_6645, wire_6607, wire_6606, wire_6586, wire_6567, wire_6566, wire_6527, wire_6526, wire_1123, wire_609, wire_10844, wire_6643, wire_6605, wire_6604, wire_6594, wire_6565, wire_6564, wire_6525, wire_6524, wire_1123, wire_605, wire_10836, wire_6641, wire_6602, wire_6601, wire_6600, wire_6561, wire_6560, wire_6521, wire_6520, wire_1123, wire_605, wire_10828, wire_6639, wire_6610, wire_6599, wire_6598, wire_6559, wire_6558, wire_6519, wire_6518, wire_1123, wire_605, wire_10820, wire_6637, wire_6618, wire_6597, wire_6596, wire_6557, wire_6556, wire_6517, wire_6516, wire_1119, wire_605, wire_10812, wire_6635, wire_6626, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512, wire_1119, wire_605, wire_10804, wire_6633, wire_6591, wire_6590, wire_6551, wire_6550, wire_6514, wire_6511, wire_6510, wire_1119, wire_605, wire_10979, wire_7049, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_6906, wire_1119, wire_10977, wire_7021, wire_7018, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_1119, wire_10975, wire_7023, wire_7013, wire_7012, wire_7010, wire_6973, wire_6972, wire_6933, wire_6932, wire_1119, wire_10973, wire_7025, wire_7009, wire_7008, wire_7002, wire_6969, wire_6968, wire_6929, wire_6928, wire_609, wire_10971, wire_7027, wire_7007, wire_7006, wire_6994, wire_6967, wire_6966, wire_6927, wire_6926, wire_609, wire_10969, wire_7029, wire_7005, wire_7004, wire_6986, wire_6965, wire_6964, wire_6925, wire_6924, wire_609, wire_10967, wire_7031, wire_7001, wire_7000, wire_6978, wire_6961, wire_6960, wire_6921, wire_6920, wire_1123, wire_609, wire_10965, wire_7033, wire_6999, wire_6998, wire_6970, wire_6959, wire_6958, wire_6919, wire_6918, wire_1123, wire_609, wire_10963, wire_7035, wire_6997, wire_6996, wire_6962, wire_6957, wire_6956, wire_6917, wire_6916, wire_1123, wire_609, wire_10961, wire_7037, wire_6993, wire_6992, wire_6954, wire_6953, wire_6952, wire_6913, wire_6912, wire_1123, wire_605, wire_10959, wire_7039, wire_6991, wire_6990, wire_6951, wire_6950, wire_6946, wire_6911, wire_6910, wire_1123, wire_605, wire_10957, wire_7041, wire_6989, wire_6988, wire_6949, wire_6948, wire_6938, wire_6909, wire_6908, wire_1123, wire_605, wire_10955, wire_7043, wire_6985, wire_6984, wire_6945, wire_6944, wire_6930, wire_6905, wire_6904, wire_1119, wire_605, wire_10953, wire_7045, wire_6983, wire_6982, wire_6943, wire_6942, wire_6922, wire_6903, wire_6902, wire_1119, wire_605, wire_10951, wire_7047, wire_6981, wire_6980, wire_6941, wire_6940, wire_6914, wire_6901, wire_6900, wire_1119, wire_605, wire_10953, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10910, wire_7049, wire_648, wire_10465, wire_10464, wire_10529, wire_10528, wire_10589, wire_10526, wire_10573, wire_10462, wire_10955, wire_10915, wire_10914, wire_10902, wire_10875, wire_10874, wire_10835, wire_10834, wire_7047, wire_648, wire_10559, wire_10558, wire_10523, wire_10522, wire_10543, wire_10542, wire_10521, wire_10520, wire_10957, wire_10913, wire_10912, wire_10894, wire_10873, wire_10872, wire_10833, wire_10832, wire_7045, wire_648, wire_10587, wire_10518, wire_10459, wire_10458, wire_10557, wire_10556, wire_10515, wire_10514, wire_10959, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10886, wire_7043, wire_608, wire_10513, wire_10512, wire_10457, wire_10456, wire_10571, wire_10454, wire_10585, wire_10510, wire_10961, wire_10907, wire_10906, wire_10878, wire_10867, wire_10866, wire_10827, wire_10826, wire_7041, wire_608, wire_10541, wire_10540, wire_10451, wire_10450, wire_10555, wire_10554, wire_10449, wire_10448, wire_10963, wire_10905, wire_10904, wire_10870, wire_10865, wire_10864, wire_10825, wire_10824, wire_7039, wire_608, wire_10569, wire_10446, wire_10507, wire_10506, wire_10539, wire_10538, wire_10443, wire_10442, wire_10965, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10862, wire_7037, wire_652, wire_608, wire_10441, wire_10440, wire_10505, wire_10504, wire_10583, wire_10502, wire_10567, wire_10438, wire_10967, wire_10899, wire_10898, wire_10859, wire_10858, wire_10854, wire_10819, wire_10818, wire_7035, wire_652, wire_608, wire_10553, wire_10552, wire_10499, wire_10498, wire_10537, wire_10536, wire_10497, wire_10496, wire_10969, wire_10897, wire_10896, wire_10857, wire_10856, wire_10846, wire_10817, wire_10816, wire_7033, wire_652, wire_608, wire_10581, wire_10494, wire_10435, wire_10434, wire_10551, wire_10550, wire_10491, wire_10490, wire_10971, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10838, wire_7031, wire_652, wire_604, wire_10489, wire_10488, wire_652, wire_10433, wire_10432, wire_652, wire_10565, wire_10430, wire_652, wire_10579, wire_10486, wire_652, wire_10973, wire_10891, wire_10890, wire_10851, wire_10850, wire_10830, wire_10811, wire_10810, wire_7029, wire_652, wire_604, wire_10535, wire_10534, wire_652, wire_10427, wire_10426, wire_652, wire_10549, wire_10548, wire_648, wire_10425, wire_10424, wire_648, wire_10975, wire_10889, wire_10888, wire_10849, wire_10848, wire_10822, wire_10809, wire_10808, wire_7027, wire_652, wire_604, wire_10563, wire_10422, wire_648, wire_10483, wire_10482, wire_648, wire_10533, wire_10532, wire_648, wire_10419, wire_10418, wire_648, wire_10977, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10814, wire_7025, wire_648, wire_604, wire_10417, wire_10416, wire_608, wire_10481, wire_10480, wire_608, wire_10577, wire_10478, wire_608, wire_10561, wire_10414, wire_608, wire_10979, wire_10883, wire_10882, wire_10843, wire_10842, wire_10806, wire_10803, wire_10802, wire_7023, wire_648, wire_604, wire_10547, wire_10546, wire_608, wire_10475, wire_10474, wire_608, wire_10531, wire_10530, wire_604, wire_10473, wire_10472, wire_604, wire_10951, wire_10918, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_7021, wire_648, wire_604, wire_10575, wire_10470, wire_604, wire_10411, wire_10410, wire_604, wire_10545, wire_10544, wire_604, wire_10467, wire_10466, wire_604};
    // CHNAXY TOTAL: 621
    assign wire_6900 = lut_tile_2_1_chanxy_out[0];
    assign wire_6902 = lut_tile_2_1_chanxy_out[1];
    assign wire_6904 = lut_tile_2_1_chanxy_out[2];
    assign wire_6906 = lut_tile_2_1_chanxy_out[3];
    assign wire_6907 = lut_tile_2_1_chanxy_out[4];
    assign wire_6908 = lut_tile_2_1_chanxy_out[5];
    assign wire_6910 = lut_tile_2_1_chanxy_out[6];
    assign wire_6912 = lut_tile_2_1_chanxy_out[7];
    assign wire_6914 = lut_tile_2_1_chanxy_out[8];
    assign wire_6915 = lut_tile_2_1_chanxy_out[9];
    assign wire_6916 = lut_tile_2_1_chanxy_out[10];
    assign wire_6918 = lut_tile_2_1_chanxy_out[11];
    assign wire_6920 = lut_tile_2_1_chanxy_out[12];
    assign wire_6922 = lut_tile_2_1_chanxy_out[13];
    assign wire_6923 = lut_tile_2_1_chanxy_out[14];
    assign wire_6924 = lut_tile_2_1_chanxy_out[15];
    assign wire_6926 = lut_tile_2_1_chanxy_out[16];
    assign wire_6928 = lut_tile_2_1_chanxy_out[17];
    assign wire_6930 = lut_tile_2_1_chanxy_out[18];
    assign wire_6931 = lut_tile_2_1_chanxy_out[19];
    assign wire_6932 = lut_tile_2_1_chanxy_out[20];
    assign wire_6934 = lut_tile_2_1_chanxy_out[21];
    assign wire_6936 = lut_tile_2_1_chanxy_out[22];
    assign wire_6938 = lut_tile_2_1_chanxy_out[23];
    assign wire_6939 = lut_tile_2_1_chanxy_out[24];
    assign wire_6940 = lut_tile_2_1_chanxy_out[25];
    assign wire_6942 = lut_tile_2_1_chanxy_out[26];
    assign wire_6944 = lut_tile_2_1_chanxy_out[27];
    assign wire_6946 = lut_tile_2_1_chanxy_out[28];
    assign wire_6947 = lut_tile_2_1_chanxy_out[29];
    assign wire_6948 = lut_tile_2_1_chanxy_out[30];
    assign wire_6950 = lut_tile_2_1_chanxy_out[31];
    assign wire_6952 = lut_tile_2_1_chanxy_out[32];
    assign wire_6954 = lut_tile_2_1_chanxy_out[33];
    assign wire_6955 = lut_tile_2_1_chanxy_out[34];
    assign wire_6956 = lut_tile_2_1_chanxy_out[35];
    assign wire_6958 = lut_tile_2_1_chanxy_out[36];
    assign wire_6960 = lut_tile_2_1_chanxy_out[37];
    assign wire_6962 = lut_tile_2_1_chanxy_out[38];
    assign wire_6963 = lut_tile_2_1_chanxy_out[39];
    assign wire_6964 = lut_tile_2_1_chanxy_out[40];
    assign wire_6966 = lut_tile_2_1_chanxy_out[41];
    assign wire_6968 = lut_tile_2_1_chanxy_out[42];
    assign wire_6970 = lut_tile_2_1_chanxy_out[43];
    assign wire_6971 = lut_tile_2_1_chanxy_out[44];
    assign wire_6972 = lut_tile_2_1_chanxy_out[45];
    assign wire_6974 = lut_tile_2_1_chanxy_out[46];
    assign wire_6976 = lut_tile_2_1_chanxy_out[47];
    assign wire_6978 = lut_tile_2_1_chanxy_out[48];
    assign wire_6979 = lut_tile_2_1_chanxy_out[49];
    assign wire_6980 = lut_tile_2_1_chanxy_out[50];
    assign wire_6982 = lut_tile_2_1_chanxy_out[51];
    assign wire_6984 = lut_tile_2_1_chanxy_out[52];
    assign wire_6986 = lut_tile_2_1_chanxy_out[53];
    assign wire_6987 = lut_tile_2_1_chanxy_out[54];
    assign wire_6988 = lut_tile_2_1_chanxy_out[55];
    assign wire_6990 = lut_tile_2_1_chanxy_out[56];
    assign wire_6992 = lut_tile_2_1_chanxy_out[57];
    assign wire_6994 = lut_tile_2_1_chanxy_out[58];
    assign wire_6995 = lut_tile_2_1_chanxy_out[59];
    assign wire_6996 = lut_tile_2_1_chanxy_out[60];
    assign wire_6998 = lut_tile_2_1_chanxy_out[61];
    assign wire_7000 = lut_tile_2_1_chanxy_out[62];
    assign wire_7002 = lut_tile_2_1_chanxy_out[63];
    assign wire_7003 = lut_tile_2_1_chanxy_out[64];
    assign wire_7004 = lut_tile_2_1_chanxy_out[65];
    assign wire_7006 = lut_tile_2_1_chanxy_out[66];
    assign wire_7008 = lut_tile_2_1_chanxy_out[67];
    assign wire_7010 = lut_tile_2_1_chanxy_out[68];
    assign wire_7011 = lut_tile_2_1_chanxy_out[69];
    assign wire_7012 = lut_tile_2_1_chanxy_out[70];
    assign wire_7014 = lut_tile_2_1_chanxy_out[71];
    assign wire_7016 = lut_tile_2_1_chanxy_out[72];
    assign wire_7018 = lut_tile_2_1_chanxy_out[73];
    assign wire_7019 = lut_tile_2_1_chanxy_out[74];
    assign wire_10807 = lut_tile_2_1_chanxy_out[75];
    assign wire_10815 = lut_tile_2_1_chanxy_out[76];
    assign wire_10823 = lut_tile_2_1_chanxy_out[77];
    assign wire_10831 = lut_tile_2_1_chanxy_out[78];
    assign wire_10839 = lut_tile_2_1_chanxy_out[79];
    assign wire_10847 = lut_tile_2_1_chanxy_out[80];
    assign wire_10855 = lut_tile_2_1_chanxy_out[81];
    assign wire_10863 = lut_tile_2_1_chanxy_out[82];
    assign wire_10871 = lut_tile_2_1_chanxy_out[83];
    assign wire_10879 = lut_tile_2_1_chanxy_out[84];
    assign wire_10887 = lut_tile_2_1_chanxy_out[85];
    assign wire_10895 = lut_tile_2_1_chanxy_out[86];
    assign wire_10903 = lut_tile_2_1_chanxy_out[87];
    assign wire_10911 = lut_tile_2_1_chanxy_out[88];
    assign wire_10919 = lut_tile_2_1_chanxy_out[89];
    assign wire_10920 = lut_tile_2_1_chanxy_out[90];
    assign wire_10922 = lut_tile_2_1_chanxy_out[91];
    assign wire_10924 = lut_tile_2_1_chanxy_out[92];
    assign wire_10926 = lut_tile_2_1_chanxy_out[93];
    assign wire_10928 = lut_tile_2_1_chanxy_out[94];
    assign wire_10930 = lut_tile_2_1_chanxy_out[95];
    assign wire_10932 = lut_tile_2_1_chanxy_out[96];
    assign wire_10934 = lut_tile_2_1_chanxy_out[97];
    assign wire_10936 = lut_tile_2_1_chanxy_out[98];
    assign wire_10938 = lut_tile_2_1_chanxy_out[99];
    assign wire_10940 = lut_tile_2_1_chanxy_out[100];
    assign wire_10942 = lut_tile_2_1_chanxy_out[101];
    assign wire_10944 = lut_tile_2_1_chanxy_out[102];
    assign wire_10946 = lut_tile_2_1_chanxy_out[103];
    assign wire_10948 = lut_tile_2_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_2_2_chanxy_in = {wire_11308, wire_6661, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6524, wire_1635, wire_11300, wire_6689, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_6532, wire_1635, wire_11292, wire_6687, wire_6623, wire_6622, wire_6583, wire_6582, wire_6543, wire_6542, wire_6540, wire_1635, wire_11284, wire_6685, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6548, wire_1125, wire_11276, wire_6683, wire_6617, wire_6616, wire_6577, wire_6576, wire_6556, wire_6537, wire_6536, wire_1125, wire_11268, wire_6681, wire_6615, wire_6614, wire_6575, wire_6574, wire_6564, wire_6535, wire_6534, wire_1125, wire_11260, wire_6679, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6572, wire_1639, wire_1125, wire_11252, wire_6677, wire_6609, wire_6608, wire_6580, wire_6569, wire_6568, wire_6529, wire_6528, wire_1639, wire_1125, wire_11244, wire_6675, wire_6607, wire_6606, wire_6588, wire_6567, wire_6566, wire_6527, wire_6526, wire_1639, wire_1125, wire_11236, wire_6673, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6596, wire_1639, wire_1121, wire_11228, wire_6671, wire_6604, wire_6601, wire_6600, wire_6561, wire_6560, wire_6521, wire_6520, wire_1639, wire_1121, wire_11220, wire_6669, wire_6612, wire_6599, wire_6598, wire_6559, wire_6558, wire_6519, wire_6518, wire_1639, wire_1121, wire_11212, wire_6667, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6620, wire_1635, wire_1121, wire_11204, wire_6665, wire_6628, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512, wire_1635, wire_1121, wire_11196, wire_6663, wire_6591, wire_6590, wire_6551, wire_6550, wire_6516, wire_6511, wire_6510, wire_1635, wire_1121, wire_11369, wire_7079, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6900, wire_1635, wire_11367, wire_7051, wire_7017, wire_7016, wire_7012, wire_6977, wire_6976, wire_6937, wire_6936, wire_1635, wire_11365, wire_7053, wire_7015, wire_7014, wire_7004, wire_6975, wire_6974, wire_6935, wire_6934, wire_1635, wire_11363, wire_7055, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6996, wire_1125, wire_11361, wire_7057, wire_7009, wire_7008, wire_6988, wire_6969, wire_6968, wire_6929, wire_6928, wire_1125, wire_11359, wire_7059, wire_7007, wire_7006, wire_6980, wire_6967, wire_6966, wire_6927, wire_6926, wire_1125, wire_11357, wire_7061, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6972, wire_1639, wire_1125, wire_11355, wire_7063, wire_7001, wire_7000, wire_6964, wire_6961, wire_6960, wire_6921, wire_6920, wire_1639, wire_1125, wire_11353, wire_7065, wire_6999, wire_6998, wire_6959, wire_6958, wire_6956, wire_6919, wire_6918, wire_1639, wire_1125, wire_11351, wire_7067, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6948, wire_1639, wire_1121, wire_11349, wire_7069, wire_6993, wire_6992, wire_6953, wire_6952, wire_6940, wire_6913, wire_6912, wire_1639, wire_1121, wire_11347, wire_7071, wire_6991, wire_6990, wire_6951, wire_6950, wire_6932, wire_6911, wire_6910, wire_1639, wire_1121, wire_11345, wire_7073, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_6924, wire_1635, wire_1121, wire_11343, wire_7075, wire_6985, wire_6984, wire_6945, wire_6944, wire_6916, wire_6905, wire_6904, wire_1635, wire_1121, wire_11341, wire_7077, wire_6983, wire_6982, wire_6943, wire_6942, wire_6908, wire_6903, wire_6902, wire_1635, wire_1121, wire_10977, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10918, wire_7018, wire_1164, wire_10975, wire_10915, wire_10914, wire_10875, wire_10874, wire_10835, wire_10834, wire_10806, wire_7010, wire_1164, wire_10973, wire_10913, wire_10912, wire_10873, wire_10872, wire_10833, wire_10832, wire_10814, wire_7002, wire_1164, wire_10971, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10822, wire_6994, wire_1124, wire_10969, wire_10907, wire_10906, wire_10867, wire_10866, wire_10830, wire_10827, wire_10826, wire_6986, wire_1124, wire_10967, wire_10905, wire_10904, wire_10865, wire_10864, wire_10838, wire_10825, wire_10824, wire_6978, wire_1124, wire_10965, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10846, wire_6970, wire_1168, wire_1124, wire_10963, wire_10899, wire_10898, wire_10859, wire_10858, wire_10854, wire_10819, wire_10818, wire_6962, wire_1168, wire_1124, wire_10961, wire_10897, wire_10896, wire_10862, wire_10857, wire_10856, wire_10817, wire_10816, wire_6954, wire_1168, wire_1124, wire_10959, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10870, wire_6946, wire_1168, wire_1120, wire_10957, wire_10891, wire_10890, wire_10878, wire_10851, wire_10850, wire_10811, wire_10810, wire_6938, wire_1168, wire_1120, wire_10955, wire_10889, wire_10888, wire_10886, wire_10849, wire_10848, wire_10809, wire_10808, wire_6930, wire_1168, wire_1120, wire_10953, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10894, wire_6922, wire_1164, wire_1120, wire_10951, wire_10902, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_6914, wire_1164, wire_1120, wire_10979, wire_10910, wire_10881, wire_10880, wire_10841, wire_10840, wire_10801, wire_10800, wire_6906, wire_1164, wire_1120, wire_11343, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11294, wire_7079, wire_1164, wire_11345, wire_11307, wire_11306, wire_11286, wire_11267, wire_11266, wire_11227, wire_11226, wire_7077, wire_1164, wire_11347, wire_11305, wire_11304, wire_11278, wire_11265, wire_11264, wire_11225, wire_11224, wire_7075, wire_1164, wire_11349, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11270, wire_7073, wire_1124, wire_11351, wire_11299, wire_11298, wire_11262, wire_11259, wire_11258, wire_11219, wire_11218, wire_7071, wire_1124, wire_11353, wire_11297, wire_11296, wire_11257, wire_11256, wire_11254, wire_11217, wire_11216, wire_7069, wire_1124, wire_11355, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11246, wire_7067, wire_1168, wire_1124, wire_11357, wire_11291, wire_11290, wire_11251, wire_11250, wire_11238, wire_11211, wire_11210, wire_7065, wire_1168, wire_1124, wire_11359, wire_11289, wire_11288, wire_11249, wire_11248, wire_11230, wire_11209, wire_11208, wire_7063, wire_1168, wire_1124, wire_11361, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11222, wire_7061, wire_1168, wire_1120, wire_11363, wire_11283, wire_11282, wire_11243, wire_11242, wire_11214, wire_11203, wire_11202, wire_7059, wire_1168, wire_1120, wire_11365, wire_11281, wire_11280, wire_11241, wire_11240, wire_11206, wire_11201, wire_11200, wire_7057, wire_1168, wire_1120, wire_11367, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11198, wire_7055, wire_1164, wire_1120, wire_11369, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_11190, wire_7053, wire_1164, wire_1120, wire_11341, wire_11302, wire_11273, wire_11272, wire_11233, wire_11232, wire_11193, wire_11192, wire_7051, wire_1164, wire_1120};
    // CHNAXY TOTAL: 636
    assign wire_6901 = lut_tile_2_2_chanxy_out[0];
    assign wire_6909 = lut_tile_2_2_chanxy_out[1];
    assign wire_6917 = lut_tile_2_2_chanxy_out[2];
    assign wire_6925 = lut_tile_2_2_chanxy_out[3];
    assign wire_6933 = lut_tile_2_2_chanxy_out[4];
    assign wire_6941 = lut_tile_2_2_chanxy_out[5];
    assign wire_6949 = lut_tile_2_2_chanxy_out[6];
    assign wire_6957 = lut_tile_2_2_chanxy_out[7];
    assign wire_6965 = lut_tile_2_2_chanxy_out[8];
    assign wire_6973 = lut_tile_2_2_chanxy_out[9];
    assign wire_6981 = lut_tile_2_2_chanxy_out[10];
    assign wire_6989 = lut_tile_2_2_chanxy_out[11];
    assign wire_6997 = lut_tile_2_2_chanxy_out[12];
    assign wire_7005 = lut_tile_2_2_chanxy_out[13];
    assign wire_7013 = lut_tile_2_2_chanxy_out[14];
    assign wire_7020 = lut_tile_2_2_chanxy_out[15];
    assign wire_7022 = lut_tile_2_2_chanxy_out[16];
    assign wire_7024 = lut_tile_2_2_chanxy_out[17];
    assign wire_7026 = lut_tile_2_2_chanxy_out[18];
    assign wire_7028 = lut_tile_2_2_chanxy_out[19];
    assign wire_7030 = lut_tile_2_2_chanxy_out[20];
    assign wire_7032 = lut_tile_2_2_chanxy_out[21];
    assign wire_7034 = lut_tile_2_2_chanxy_out[22];
    assign wire_7036 = lut_tile_2_2_chanxy_out[23];
    assign wire_7038 = lut_tile_2_2_chanxy_out[24];
    assign wire_7040 = lut_tile_2_2_chanxy_out[25];
    assign wire_7042 = lut_tile_2_2_chanxy_out[26];
    assign wire_7044 = lut_tile_2_2_chanxy_out[27];
    assign wire_7046 = lut_tile_2_2_chanxy_out[28];
    assign wire_7048 = lut_tile_2_2_chanxy_out[29];
    assign wire_11191 = lut_tile_2_2_chanxy_out[30];
    assign wire_11199 = lut_tile_2_2_chanxy_out[31];
    assign wire_11207 = lut_tile_2_2_chanxy_out[32];
    assign wire_11215 = lut_tile_2_2_chanxy_out[33];
    assign wire_11223 = lut_tile_2_2_chanxy_out[34];
    assign wire_11231 = lut_tile_2_2_chanxy_out[35];
    assign wire_11239 = lut_tile_2_2_chanxy_out[36];
    assign wire_11247 = lut_tile_2_2_chanxy_out[37];
    assign wire_11255 = lut_tile_2_2_chanxy_out[38];
    assign wire_11263 = lut_tile_2_2_chanxy_out[39];
    assign wire_11271 = lut_tile_2_2_chanxy_out[40];
    assign wire_11279 = lut_tile_2_2_chanxy_out[41];
    assign wire_11287 = lut_tile_2_2_chanxy_out[42];
    assign wire_11295 = lut_tile_2_2_chanxy_out[43];
    assign wire_11303 = lut_tile_2_2_chanxy_out[44];
    assign wire_11310 = lut_tile_2_2_chanxy_out[45];
    assign wire_11312 = lut_tile_2_2_chanxy_out[46];
    assign wire_11314 = lut_tile_2_2_chanxy_out[47];
    assign wire_11316 = lut_tile_2_2_chanxy_out[48];
    assign wire_11318 = lut_tile_2_2_chanxy_out[49];
    assign wire_11320 = lut_tile_2_2_chanxy_out[50];
    assign wire_11322 = lut_tile_2_2_chanxy_out[51];
    assign wire_11324 = lut_tile_2_2_chanxy_out[52];
    assign wire_11326 = lut_tile_2_2_chanxy_out[53];
    assign wire_11328 = lut_tile_2_2_chanxy_out[54];
    assign wire_11330 = lut_tile_2_2_chanxy_out[55];
    assign wire_11332 = lut_tile_2_2_chanxy_out[56];
    assign wire_11334 = lut_tile_2_2_chanxy_out[57];
    assign wire_11336 = lut_tile_2_2_chanxy_out[58];
    assign wire_11338 = lut_tile_2_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_3_chanxy_in = {wire_11692, wire_6691, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6518, wire_2151, wire_11684, wire_6719, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6526, wire_2151, wire_11676, wire_6717, wire_6625, wire_6624, wire_6585, wire_6584, wire_6545, wire_6544, wire_6534, wire_2151, wire_11668, wire_6715, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6542, wire_1641, wire_11660, wire_6713, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6550, wire_1641, wire_11652, wire_6711, wire_6617, wire_6616, wire_6577, wire_6576, wire_6558, wire_6537, wire_6536, wire_1641, wire_11644, wire_6709, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6566, wire_2155, wire_1641, wire_11636, wire_6707, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6574, wire_2155, wire_1641, wire_11628, wire_6705, wire_6609, wire_6608, wire_6582, wire_6569, wire_6568, wire_6529, wire_6528, wire_2155, wire_1641, wire_11620, wire_6703, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6590, wire_2155, wire_1637, wire_11612, wire_6701, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6598, wire_2155, wire_1637, wire_11604, wire_6699, wire_6606, wire_6601, wire_6600, wire_6561, wire_6560, wire_6521, wire_6520, wire_2155, wire_1637, wire_11596, wire_6697, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6614, wire_2151, wire_1637, wire_11588, wire_6695, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6622, wire_2151, wire_1637, wire_11580, wire_6693, wire_6593, wire_6592, wire_6553, wire_6552, wire_6513, wire_6512, wire_6510, wire_2151, wire_1637, wire_11759, wire_7109, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6902, wire_2151, wire_11757, wire_7081, wire_7017, wire_7016, wire_7014, wire_6977, wire_6976, wire_6937, wire_6936, wire_2151, wire_11755, wire_7083, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_7006, wire_2151, wire_11753, wire_7085, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6998, wire_1641, wire_11751, wire_7087, wire_7009, wire_7008, wire_6990, wire_6969, wire_6968, wire_6929, wire_6928, wire_1641, wire_11749, wire_7089, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6982, wire_1641, wire_11747, wire_7091, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6974, wire_2155, wire_1641, wire_11745, wire_7093, wire_7001, wire_7000, wire_6966, wire_6961, wire_6960, wire_6921, wire_6920, wire_2155, wire_1641, wire_11743, wire_7095, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_6958, wire_2155, wire_1641, wire_11741, wire_7097, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6950, wire_2155, wire_1637, wire_11739, wire_7099, wire_6993, wire_6992, wire_6953, wire_6952, wire_6942, wire_6913, wire_6912, wire_2155, wire_1637, wire_11737, wire_7101, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_6934, wire_2155, wire_1637, wire_11735, wire_7103, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_6926, wire_2151, wire_1637, wire_11733, wire_7105, wire_6985, wire_6984, wire_6945, wire_6944, wire_6918, wire_6905, wire_6904, wire_2151, wire_1637, wire_11731, wire_7107, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_6910, wire_2151, wire_1637, wire_11367, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11302, wire_7012, wire_1680, wire_11365, wire_11307, wire_11306, wire_11267, wire_11266, wire_11227, wire_11226, wire_11190, wire_7004, wire_1680, wire_11363, wire_11305, wire_11304, wire_11265, wire_11264, wire_11225, wire_11224, wire_11198, wire_6996, wire_1680, wire_11361, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11206, wire_6988, wire_1640, wire_11359, wire_11299, wire_11298, wire_11259, wire_11258, wire_11219, wire_11218, wire_11214, wire_6980, wire_1640, wire_11357, wire_11297, wire_11296, wire_11257, wire_11256, wire_11222, wire_11217, wire_11216, wire_6972, wire_1640, wire_11355, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11230, wire_6964, wire_1684, wire_1640, wire_11353, wire_11291, wire_11290, wire_11251, wire_11250, wire_11238, wire_11211, wire_11210, wire_6956, wire_1684, wire_1640, wire_11351, wire_11289, wire_11288, wire_11249, wire_11248, wire_11246, wire_11209, wire_11208, wire_6948, wire_1684, wire_1640, wire_11349, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11254, wire_6940, wire_1684, wire_1636, wire_11347, wire_11283, wire_11282, wire_11262, wire_11243, wire_11242, wire_11203, wire_11202, wire_6932, wire_1684, wire_1636, wire_11345, wire_11281, wire_11280, wire_11270, wire_11241, wire_11240, wire_11201, wire_11200, wire_6924, wire_1684, wire_1636, wire_11343, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11278, wire_6916, wire_1680, wire_1636, wire_11341, wire_11286, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_6908, wire_1680, wire_1636, wire_11369, wire_11294, wire_11273, wire_11272, wire_11233, wire_11232, wire_11193, wire_11192, wire_6900, wire_1680, wire_1636, wire_11733, wire_11699, wire_11698, wire_11686, wire_11659, wire_11658, wire_11619, wire_11618, wire_7109, wire_1680, wire_11735, wire_11697, wire_11696, wire_11678, wire_11657, wire_11656, wire_11617, wire_11616, wire_7107, wire_1680, wire_11737, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11670, wire_7105, wire_1680, wire_11739, wire_11691, wire_11690, wire_11662, wire_11651, wire_11650, wire_11611, wire_11610, wire_7103, wire_1640, wire_11741, wire_11689, wire_11688, wire_11654, wire_11649, wire_11648, wire_11609, wire_11608, wire_7101, wire_1640, wire_11743, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11646, wire_7099, wire_1640, wire_11745, wire_11683, wire_11682, wire_11643, wire_11642, wire_11638, wire_11603, wire_11602, wire_7097, wire_1684, wire_1640, wire_11747, wire_11681, wire_11680, wire_11641, wire_11640, wire_11630, wire_11601, wire_11600, wire_7095, wire_1684, wire_1640, wire_11749, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11622, wire_7093, wire_1684, wire_1640, wire_11751, wire_11675, wire_11674, wire_11635, wire_11634, wire_11614, wire_11595, wire_11594, wire_7091, wire_1684, wire_1636, wire_11753, wire_11673, wire_11672, wire_11633, wire_11632, wire_11606, wire_11593, wire_11592, wire_7089, wire_1684, wire_1636, wire_11755, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11598, wire_7087, wire_1684, wire_1636, wire_11757, wire_11667, wire_11666, wire_11627, wire_11626, wire_11590, wire_11587, wire_11586, wire_7085, wire_1680, wire_1636, wire_11759, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_11582, wire_7083, wire_1680, wire_1636, wire_11731, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11694, wire_7081, wire_1680, wire_1636};
    // CHNAXY TOTAL: 636
    assign wire_6903 = lut_tile_2_3_chanxy_out[0];
    assign wire_6911 = lut_tile_2_3_chanxy_out[1];
    assign wire_6919 = lut_tile_2_3_chanxy_out[2];
    assign wire_6927 = lut_tile_2_3_chanxy_out[3];
    assign wire_6935 = lut_tile_2_3_chanxy_out[4];
    assign wire_6943 = lut_tile_2_3_chanxy_out[5];
    assign wire_6951 = lut_tile_2_3_chanxy_out[6];
    assign wire_6959 = lut_tile_2_3_chanxy_out[7];
    assign wire_6967 = lut_tile_2_3_chanxy_out[8];
    assign wire_6975 = lut_tile_2_3_chanxy_out[9];
    assign wire_6983 = lut_tile_2_3_chanxy_out[10];
    assign wire_6991 = lut_tile_2_3_chanxy_out[11];
    assign wire_6999 = lut_tile_2_3_chanxy_out[12];
    assign wire_7007 = lut_tile_2_3_chanxy_out[13];
    assign wire_7015 = lut_tile_2_3_chanxy_out[14];
    assign wire_7050 = lut_tile_2_3_chanxy_out[15];
    assign wire_7052 = lut_tile_2_3_chanxy_out[16];
    assign wire_7054 = lut_tile_2_3_chanxy_out[17];
    assign wire_7056 = lut_tile_2_3_chanxy_out[18];
    assign wire_7058 = lut_tile_2_3_chanxy_out[19];
    assign wire_7060 = lut_tile_2_3_chanxy_out[20];
    assign wire_7062 = lut_tile_2_3_chanxy_out[21];
    assign wire_7064 = lut_tile_2_3_chanxy_out[22];
    assign wire_7066 = lut_tile_2_3_chanxy_out[23];
    assign wire_7068 = lut_tile_2_3_chanxy_out[24];
    assign wire_7070 = lut_tile_2_3_chanxy_out[25];
    assign wire_7072 = lut_tile_2_3_chanxy_out[26];
    assign wire_7074 = lut_tile_2_3_chanxy_out[27];
    assign wire_7076 = lut_tile_2_3_chanxy_out[28];
    assign wire_7078 = lut_tile_2_3_chanxy_out[29];
    assign wire_11583 = lut_tile_2_3_chanxy_out[30];
    assign wire_11591 = lut_tile_2_3_chanxy_out[31];
    assign wire_11599 = lut_tile_2_3_chanxy_out[32];
    assign wire_11607 = lut_tile_2_3_chanxy_out[33];
    assign wire_11615 = lut_tile_2_3_chanxy_out[34];
    assign wire_11623 = lut_tile_2_3_chanxy_out[35];
    assign wire_11631 = lut_tile_2_3_chanxy_out[36];
    assign wire_11639 = lut_tile_2_3_chanxy_out[37];
    assign wire_11647 = lut_tile_2_3_chanxy_out[38];
    assign wire_11655 = lut_tile_2_3_chanxy_out[39];
    assign wire_11663 = lut_tile_2_3_chanxy_out[40];
    assign wire_11671 = lut_tile_2_3_chanxy_out[41];
    assign wire_11679 = lut_tile_2_3_chanxy_out[42];
    assign wire_11687 = lut_tile_2_3_chanxy_out[43];
    assign wire_11695 = lut_tile_2_3_chanxy_out[44];
    assign wire_11700 = lut_tile_2_3_chanxy_out[45];
    assign wire_11702 = lut_tile_2_3_chanxy_out[46];
    assign wire_11704 = lut_tile_2_3_chanxy_out[47];
    assign wire_11706 = lut_tile_2_3_chanxy_out[48];
    assign wire_11708 = lut_tile_2_3_chanxy_out[49];
    assign wire_11710 = lut_tile_2_3_chanxy_out[50];
    assign wire_11712 = lut_tile_2_3_chanxy_out[51];
    assign wire_11714 = lut_tile_2_3_chanxy_out[52];
    assign wire_11716 = lut_tile_2_3_chanxy_out[53];
    assign wire_11718 = lut_tile_2_3_chanxy_out[54];
    assign wire_11720 = lut_tile_2_3_chanxy_out[55];
    assign wire_11722 = lut_tile_2_3_chanxy_out[56];
    assign wire_11724 = lut_tile_2_3_chanxy_out[57];
    assign wire_11726 = lut_tile_2_3_chanxy_out[58];
    assign wire_11728 = lut_tile_2_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_4_chanxy_in = {wire_12084, wire_6721, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6520, wire_2667, wire_12076, wire_6749, wire_6659, wire_6658, wire_6649, wire_6648, wire_6639, wire_6638, wire_6528, wire_2667, wire_12068, wire_6747, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6536, wire_2667, wire_12060, wire_6745, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6544, wire_2157, wire_12052, wire_6743, wire_6657, wire_6656, wire_6647, wire_6646, wire_6637, wire_6636, wire_6552, wire_2157, wire_12044, wire_6741, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6560, wire_2157, wire_12036, wire_6739, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6568, wire_2671, wire_2157, wire_12028, wire_6737, wire_6655, wire_6654, wire_6645, wire_6644, wire_6635, wire_6634, wire_6576, wire_2671, wire_2157, wire_12020, wire_6735, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6584, wire_2671, wire_2157, wire_12012, wire_6733, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6592, wire_2671, wire_2153, wire_12004, wire_6731, wire_6653, wire_6652, wire_6643, wire_6642, wire_6633, wire_6632, wire_6600, wire_2671, wire_2153, wire_11996, wire_6729, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6608, wire_2671, wire_2153, wire_11988, wire_6727, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6616, wire_2667, wire_2153, wire_11980, wire_6725, wire_6651, wire_6650, wire_6641, wire_6640, wire_6631, wire_6630, wire_6624, wire_2667, wire_2153, wire_11972, wire_6723, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6512, wire_2667, wire_2153, wire_12149, wire_7139, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6904, wire_2667, wire_12147, wire_7111, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7016, wire_2667, wire_12145, wire_7113, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_7008, wire_2667, wire_12143, wire_7115, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_7000, wire_2157, wire_12141, wire_7117, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_6992, wire_2157, wire_12139, wire_7119, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6984, wire_2157, wire_12137, wire_7121, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6976, wire_2671, wire_2157, wire_12135, wire_7123, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_6968, wire_2671, wire_2157, wire_12133, wire_7125, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_6960, wire_2671, wire_2157, wire_12131, wire_7127, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6952, wire_2671, wire_2153, wire_12129, wire_7129, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_6944, wire_2671, wire_2153, wire_12127, wire_7131, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_6936, wire_2671, wire_2153, wire_12125, wire_7133, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_6928, wire_2667, wire_2153, wire_12123, wire_7135, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_6920, wire_2667, wire_2153, wire_12121, wire_7137, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_6912, wire_2667, wire_2153, wire_11757, wire_11699, wire_11698, wire_11694, wire_11659, wire_11658, wire_11619, wire_11618, wire_7014, wire_2196, wire_11755, wire_11697, wire_11696, wire_11657, wire_11656, wire_11617, wire_11616, wire_11582, wire_7006, wire_2196, wire_11753, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11590, wire_6998, wire_2196, wire_11751, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_11598, wire_6990, wire_2156, wire_11749, wire_11689, wire_11688, wire_11649, wire_11648, wire_11609, wire_11608, wire_11606, wire_6982, wire_2156, wire_11747, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11614, wire_6974, wire_2156, wire_11745, wire_11683, wire_11682, wire_11643, wire_11642, wire_11622, wire_11603, wire_11602, wire_6966, wire_2200, wire_2156, wire_11743, wire_11681, wire_11680, wire_11641, wire_11640, wire_11630, wire_11601, wire_11600, wire_6958, wire_2200, wire_2156, wire_11741, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11638, wire_6950, wire_2200, wire_2156, wire_11739, wire_11675, wire_11674, wire_11646, wire_11635, wire_11634, wire_11595, wire_11594, wire_6942, wire_2200, wire_2152, wire_11737, wire_11673, wire_11672, wire_11654, wire_11633, wire_11632, wire_11593, wire_11592, wire_6934, wire_2200, wire_2152, wire_11735, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11662, wire_6926, wire_2200, wire_2152, wire_11733, wire_11670, wire_11667, wire_11666, wire_11627, wire_11626, wire_11587, wire_11586, wire_6918, wire_2196, wire_2152, wire_11731, wire_11678, wire_11665, wire_11664, wire_11625, wire_11624, wire_11585, wire_11584, wire_6910, wire_2196, wire_2152, wire_11759, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11686, wire_6902, wire_2196, wire_2152, wire_12123, wire_12089, wire_12088, wire_12078, wire_12049, wire_12048, wire_12009, wire_12008, wire_7139, wire_2196, wire_12125, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_12070, wire_7137, wire_2196, wire_12127, wire_12083, wire_12082, wire_12062, wire_12043, wire_12042, wire_12003, wire_12002, wire_7135, wire_2196, wire_12129, wire_12081, wire_12080, wire_12054, wire_12041, wire_12040, wire_12001, wire_12000, wire_7133, wire_2156, wire_12131, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12046, wire_7131, wire_2156, wire_12133, wire_12075, wire_12074, wire_12038, wire_12035, wire_12034, wire_11995, wire_11994, wire_7129, wire_2156, wire_12135, wire_12073, wire_12072, wire_12033, wire_12032, wire_12030, wire_11993, wire_11992, wire_7127, wire_2200, wire_2156, wire_12137, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12022, wire_7125, wire_2200, wire_2156, wire_12139, wire_12067, wire_12066, wire_12027, wire_12026, wire_12014, wire_11987, wire_11986, wire_7123, wire_2200, wire_2156, wire_12141, wire_12065, wire_12064, wire_12025, wire_12024, wire_12006, wire_11985, wire_11984, wire_7121, wire_2200, wire_2152, wire_12143, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_11998, wire_7119, wire_2200, wire_2152, wire_12145, wire_12059, wire_12058, wire_12019, wire_12018, wire_11990, wire_11979, wire_11978, wire_7117, wire_2200, wire_2152, wire_12147, wire_12057, wire_12056, wire_12017, wire_12016, wire_11982, wire_11977, wire_11976, wire_7115, wire_2196, wire_2152, wire_12149, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_11974, wire_7113, wire_2196, wire_2152, wire_12121, wire_12086, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7111, wire_2196, wire_2152};
    // CHNAXY TOTAL: 636
    assign wire_6905 = lut_tile_2_4_chanxy_out[0];
    assign wire_6913 = lut_tile_2_4_chanxy_out[1];
    assign wire_6921 = lut_tile_2_4_chanxy_out[2];
    assign wire_6929 = lut_tile_2_4_chanxy_out[3];
    assign wire_6937 = lut_tile_2_4_chanxy_out[4];
    assign wire_6945 = lut_tile_2_4_chanxy_out[5];
    assign wire_6953 = lut_tile_2_4_chanxy_out[6];
    assign wire_6961 = lut_tile_2_4_chanxy_out[7];
    assign wire_6969 = lut_tile_2_4_chanxy_out[8];
    assign wire_6977 = lut_tile_2_4_chanxy_out[9];
    assign wire_6985 = lut_tile_2_4_chanxy_out[10];
    assign wire_6993 = lut_tile_2_4_chanxy_out[11];
    assign wire_7001 = lut_tile_2_4_chanxy_out[12];
    assign wire_7009 = lut_tile_2_4_chanxy_out[13];
    assign wire_7017 = lut_tile_2_4_chanxy_out[14];
    assign wire_7080 = lut_tile_2_4_chanxy_out[15];
    assign wire_7082 = lut_tile_2_4_chanxy_out[16];
    assign wire_7084 = lut_tile_2_4_chanxy_out[17];
    assign wire_7086 = lut_tile_2_4_chanxy_out[18];
    assign wire_7088 = lut_tile_2_4_chanxy_out[19];
    assign wire_7090 = lut_tile_2_4_chanxy_out[20];
    assign wire_7092 = lut_tile_2_4_chanxy_out[21];
    assign wire_7094 = lut_tile_2_4_chanxy_out[22];
    assign wire_7096 = lut_tile_2_4_chanxy_out[23];
    assign wire_7098 = lut_tile_2_4_chanxy_out[24];
    assign wire_7100 = lut_tile_2_4_chanxy_out[25];
    assign wire_7102 = lut_tile_2_4_chanxy_out[26];
    assign wire_7104 = lut_tile_2_4_chanxy_out[27];
    assign wire_7106 = lut_tile_2_4_chanxy_out[28];
    assign wire_7108 = lut_tile_2_4_chanxy_out[29];
    assign wire_11975 = lut_tile_2_4_chanxy_out[30];
    assign wire_11983 = lut_tile_2_4_chanxy_out[31];
    assign wire_11991 = lut_tile_2_4_chanxy_out[32];
    assign wire_11999 = lut_tile_2_4_chanxy_out[33];
    assign wire_12007 = lut_tile_2_4_chanxy_out[34];
    assign wire_12015 = lut_tile_2_4_chanxy_out[35];
    assign wire_12023 = lut_tile_2_4_chanxy_out[36];
    assign wire_12031 = lut_tile_2_4_chanxy_out[37];
    assign wire_12039 = lut_tile_2_4_chanxy_out[38];
    assign wire_12047 = lut_tile_2_4_chanxy_out[39];
    assign wire_12055 = lut_tile_2_4_chanxy_out[40];
    assign wire_12063 = lut_tile_2_4_chanxy_out[41];
    assign wire_12071 = lut_tile_2_4_chanxy_out[42];
    assign wire_12079 = lut_tile_2_4_chanxy_out[43];
    assign wire_12087 = lut_tile_2_4_chanxy_out[44];
    assign wire_12090 = lut_tile_2_4_chanxy_out[45];
    assign wire_12092 = lut_tile_2_4_chanxy_out[46];
    assign wire_12094 = lut_tile_2_4_chanxy_out[47];
    assign wire_12096 = lut_tile_2_4_chanxy_out[48];
    assign wire_12098 = lut_tile_2_4_chanxy_out[49];
    assign wire_12100 = lut_tile_2_4_chanxy_out[50];
    assign wire_12102 = lut_tile_2_4_chanxy_out[51];
    assign wire_12104 = lut_tile_2_4_chanxy_out[52];
    assign wire_12106 = lut_tile_2_4_chanxy_out[53];
    assign wire_12108 = lut_tile_2_4_chanxy_out[54];
    assign wire_12110 = lut_tile_2_4_chanxy_out[55];
    assign wire_12112 = lut_tile_2_4_chanxy_out[56];
    assign wire_12114 = lut_tile_2_4_chanxy_out[57];
    assign wire_12116 = lut_tile_2_4_chanxy_out[58];
    assign wire_12118 = lut_tile_2_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_5_chanxy_in = {wire_12476, wire_6751, wire_6689, wire_6688, wire_6679, wire_6678, wire_6669, wire_6668, wire_6632, wire_3183, wire_12468, wire_6779, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6634, wire_3183, wire_12460, wire_6777, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6636, wire_3183, wire_12452, wire_6775, wire_6687, wire_6686, wire_6677, wire_6676, wire_6667, wire_6666, wire_6638, wire_2673, wire_12444, wire_6773, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6640, wire_2673, wire_12436, wire_6771, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6642, wire_2673, wire_12428, wire_6769, wire_6685, wire_6684, wire_6675, wire_6674, wire_6665, wire_6664, wire_6644, wire_3187, wire_2673, wire_12420, wire_6767, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6646, wire_3187, wire_2673, wire_12412, wire_6765, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6648, wire_3187, wire_2673, wire_12404, wire_6763, wire_6683, wire_6682, wire_6673, wire_6672, wire_6663, wire_6662, wire_6650, wire_3187, wire_2669, wire_12396, wire_6761, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6652, wire_3187, wire_2669, wire_12388, wire_6759, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6654, wire_3187, wire_2669, wire_12380, wire_6757, wire_6681, wire_6680, wire_6671, wire_6670, wire_6661, wire_6660, wire_6656, wire_3183, wire_2669, wire_12372, wire_6755, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6658, wire_3183, wire_2669, wire_12364, wire_6753, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6630, wire_3183, wire_2669, wire_12539, wire_7169, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7020, wire_3183, wire_12537, wire_7141, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7048, wire_3183, wire_12535, wire_7143, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_7046, wire_3183, wire_12533, wire_7145, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7044, wire_2673, wire_12531, wire_7147, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7042, wire_2673, wire_12529, wire_7149, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_7040, wire_2673, wire_12527, wire_7151, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7038, wire_3187, wire_2673, wire_12525, wire_7153, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7036, wire_3187, wire_2673, wire_12523, wire_7155, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_7034, wire_3187, wire_2673, wire_12521, wire_7157, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7032, wire_3187, wire_2669, wire_12519, wire_7159, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7030, wire_3187, wire_2669, wire_12517, wire_7161, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_7028, wire_3187, wire_2669, wire_12515, wire_7163, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7026, wire_3183, wire_2669, wire_12513, wire_7165, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7024, wire_3183, wire_2669, wire_12511, wire_7167, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_7022, wire_3183, wire_2669, wire_12147, wire_12089, wire_12088, wire_12086, wire_12049, wire_12048, wire_12009, wire_12008, wire_7016, wire_2712, wire_12145, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_11974, wire_7008, wire_2712, wire_12143, wire_12083, wire_12082, wire_12043, wire_12042, wire_12003, wire_12002, wire_11982, wire_7000, wire_2712, wire_12141, wire_12081, wire_12080, wire_12041, wire_12040, wire_12001, wire_12000, wire_11990, wire_6992, wire_2672, wire_12139, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_11998, wire_6984, wire_2672, wire_12137, wire_12075, wire_12074, wire_12035, wire_12034, wire_12006, wire_11995, wire_11994, wire_6976, wire_2672, wire_12135, wire_12073, wire_12072, wire_12033, wire_12032, wire_12014, wire_11993, wire_11992, wire_6968, wire_2716, wire_2672, wire_12133, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12022, wire_6960, wire_2716, wire_2672, wire_12131, wire_12067, wire_12066, wire_12030, wire_12027, wire_12026, wire_11987, wire_11986, wire_6952, wire_2716, wire_2672, wire_12129, wire_12065, wire_12064, wire_12038, wire_12025, wire_12024, wire_11985, wire_11984, wire_6944, wire_2716, wire_2668, wire_12127, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12046, wire_6936, wire_2716, wire_2668, wire_12125, wire_12059, wire_12058, wire_12054, wire_12019, wire_12018, wire_11979, wire_11978, wire_6928, wire_2716, wire_2668, wire_12123, wire_12062, wire_12057, wire_12056, wire_12017, wire_12016, wire_11977, wire_11976, wire_6920, wire_2712, wire_2668, wire_12121, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12070, wire_6912, wire_2712, wire_2668, wire_12149, wire_12078, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_6904, wire_2712, wire_2668, wire_12513, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12470, wire_7169, wire_2712, wire_12515, wire_12475, wire_12474, wire_12462, wire_12435, wire_12434, wire_12395, wire_12394, wire_7167, wire_2712, wire_12517, wire_12473, wire_12472, wire_12454, wire_12433, wire_12432, wire_12393, wire_12392, wire_7165, wire_2712, wire_12519, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12446, wire_7163, wire_2672, wire_12521, wire_12467, wire_12466, wire_12438, wire_12427, wire_12426, wire_12387, wire_12386, wire_7161, wire_2672, wire_12523, wire_12465, wire_12464, wire_12430, wire_12425, wire_12424, wire_12385, wire_12384, wire_7159, wire_2672, wire_12525, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12422, wire_7157, wire_2716, wire_2672, wire_12527, wire_12459, wire_12458, wire_12419, wire_12418, wire_12414, wire_12379, wire_12378, wire_7155, wire_2716, wire_2672, wire_12529, wire_12457, wire_12456, wire_12417, wire_12416, wire_12406, wire_12377, wire_12376, wire_7153, wire_2716, wire_2672, wire_12531, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12398, wire_7151, wire_2716, wire_2668, wire_12533, wire_12451, wire_12450, wire_12411, wire_12410, wire_12390, wire_12371, wire_12370, wire_7149, wire_2716, wire_2668, wire_12535, wire_12449, wire_12448, wire_12409, wire_12408, wire_12382, wire_12369, wire_12368, wire_7147, wire_2716, wire_2668, wire_12537, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12374, wire_7145, wire_2712, wire_2668, wire_12539, wire_12443, wire_12442, wire_12403, wire_12402, wire_12366, wire_12363, wire_12362, wire_7143, wire_2712, wire_2668, wire_12511, wire_12478, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_7141, wire_2712, wire_2668};
    // CHNAXY TOTAL: 636
    assign wire_7021 = lut_tile_2_5_chanxy_out[0];
    assign wire_7023 = lut_tile_2_5_chanxy_out[1];
    assign wire_7025 = lut_tile_2_5_chanxy_out[2];
    assign wire_7027 = lut_tile_2_5_chanxy_out[3];
    assign wire_7029 = lut_tile_2_5_chanxy_out[4];
    assign wire_7031 = lut_tile_2_5_chanxy_out[5];
    assign wire_7033 = lut_tile_2_5_chanxy_out[6];
    assign wire_7035 = lut_tile_2_5_chanxy_out[7];
    assign wire_7037 = lut_tile_2_5_chanxy_out[8];
    assign wire_7039 = lut_tile_2_5_chanxy_out[9];
    assign wire_7041 = lut_tile_2_5_chanxy_out[10];
    assign wire_7043 = lut_tile_2_5_chanxy_out[11];
    assign wire_7045 = lut_tile_2_5_chanxy_out[12];
    assign wire_7047 = lut_tile_2_5_chanxy_out[13];
    assign wire_7049 = lut_tile_2_5_chanxy_out[14];
    assign wire_7110 = lut_tile_2_5_chanxy_out[15];
    assign wire_7112 = lut_tile_2_5_chanxy_out[16];
    assign wire_7114 = lut_tile_2_5_chanxy_out[17];
    assign wire_7116 = lut_tile_2_5_chanxy_out[18];
    assign wire_7118 = lut_tile_2_5_chanxy_out[19];
    assign wire_7120 = lut_tile_2_5_chanxy_out[20];
    assign wire_7122 = lut_tile_2_5_chanxy_out[21];
    assign wire_7124 = lut_tile_2_5_chanxy_out[22];
    assign wire_7126 = lut_tile_2_5_chanxy_out[23];
    assign wire_7128 = lut_tile_2_5_chanxy_out[24];
    assign wire_7130 = lut_tile_2_5_chanxy_out[25];
    assign wire_7132 = lut_tile_2_5_chanxy_out[26];
    assign wire_7134 = lut_tile_2_5_chanxy_out[27];
    assign wire_7136 = lut_tile_2_5_chanxy_out[28];
    assign wire_7138 = lut_tile_2_5_chanxy_out[29];
    assign wire_12367 = lut_tile_2_5_chanxy_out[30];
    assign wire_12375 = lut_tile_2_5_chanxy_out[31];
    assign wire_12383 = lut_tile_2_5_chanxy_out[32];
    assign wire_12391 = lut_tile_2_5_chanxy_out[33];
    assign wire_12399 = lut_tile_2_5_chanxy_out[34];
    assign wire_12407 = lut_tile_2_5_chanxy_out[35];
    assign wire_12415 = lut_tile_2_5_chanxy_out[36];
    assign wire_12423 = lut_tile_2_5_chanxy_out[37];
    assign wire_12431 = lut_tile_2_5_chanxy_out[38];
    assign wire_12439 = lut_tile_2_5_chanxy_out[39];
    assign wire_12447 = lut_tile_2_5_chanxy_out[40];
    assign wire_12455 = lut_tile_2_5_chanxy_out[41];
    assign wire_12463 = lut_tile_2_5_chanxy_out[42];
    assign wire_12471 = lut_tile_2_5_chanxy_out[43];
    assign wire_12479 = lut_tile_2_5_chanxy_out[44];
    assign wire_12480 = lut_tile_2_5_chanxy_out[45];
    assign wire_12482 = lut_tile_2_5_chanxy_out[46];
    assign wire_12484 = lut_tile_2_5_chanxy_out[47];
    assign wire_12486 = lut_tile_2_5_chanxy_out[48];
    assign wire_12488 = lut_tile_2_5_chanxy_out[49];
    assign wire_12490 = lut_tile_2_5_chanxy_out[50];
    assign wire_12492 = lut_tile_2_5_chanxy_out[51];
    assign wire_12494 = lut_tile_2_5_chanxy_out[52];
    assign wire_12496 = lut_tile_2_5_chanxy_out[53];
    assign wire_12498 = lut_tile_2_5_chanxy_out[54];
    assign wire_12500 = lut_tile_2_5_chanxy_out[55];
    assign wire_12502 = lut_tile_2_5_chanxy_out[56];
    assign wire_12504 = lut_tile_2_5_chanxy_out[57];
    assign wire_12506 = lut_tile_2_5_chanxy_out[58];
    assign wire_12508 = lut_tile_2_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_6_chanxy_in = {wire_12868, wire_6781, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6662, wire_3699, wire_12860, wire_6809, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6664, wire_3699, wire_12852, wire_6807, wire_6719, wire_6718, wire_6709, wire_6708, wire_6699, wire_6698, wire_6666, wire_3699, wire_12844, wire_6805, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6668, wire_3189, wire_12836, wire_6803, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6670, wire_3189, wire_12828, wire_6801, wire_6717, wire_6716, wire_6707, wire_6706, wire_6697, wire_6696, wire_6672, wire_3189, wire_12820, wire_6799, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6674, wire_3703, wire_3189, wire_12812, wire_6797, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6676, wire_3703, wire_3189, wire_12804, wire_6795, wire_6715, wire_6714, wire_6705, wire_6704, wire_6695, wire_6694, wire_6678, wire_3703, wire_3189, wire_12796, wire_6793, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6680, wire_3703, wire_3185, wire_12788, wire_6791, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6682, wire_3703, wire_3185, wire_12780, wire_6789, wire_6713, wire_6712, wire_6703, wire_6702, wire_6693, wire_6692, wire_6684, wire_3703, wire_3185, wire_12772, wire_6787, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6686, wire_3699, wire_3185, wire_12764, wire_6785, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6688, wire_3699, wire_3185, wire_12756, wire_6783, wire_6711, wire_6710, wire_6701, wire_6700, wire_6691, wire_6690, wire_6660, wire_3699, wire_3185, wire_12929, wire_7199, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7050, wire_3699, wire_12927, wire_7171, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7078, wire_3699, wire_12925, wire_7173, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7076, wire_3699, wire_12923, wire_7175, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7074, wire_3189, wire_12921, wire_7177, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7072, wire_3189, wire_12919, wire_7179, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7070, wire_3189, wire_12917, wire_7181, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7068, wire_3703, wire_3189, wire_12915, wire_7183, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7066, wire_3703, wire_3189, wire_12913, wire_7185, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7064, wire_3703, wire_3189, wire_12911, wire_7187, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7062, wire_3703, wire_3185, wire_12909, wire_7189, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7060, wire_3703, wire_3185, wire_12907, wire_7191, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7058, wire_3703, wire_3185, wire_12905, wire_7193, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7056, wire_3699, wire_3185, wire_12903, wire_7195, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7054, wire_3699, wire_3185, wire_12901, wire_7197, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7052, wire_3699, wire_3185, wire_12537, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12478, wire_7048, wire_3228, wire_12535, wire_12475, wire_12474, wire_12435, wire_12434, wire_12395, wire_12394, wire_12366, wire_7046, wire_3228, wire_12533, wire_12473, wire_12472, wire_12433, wire_12432, wire_12393, wire_12392, wire_12374, wire_7044, wire_3228, wire_12531, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12382, wire_7042, wire_3188, wire_12529, wire_12467, wire_12466, wire_12427, wire_12426, wire_12390, wire_12387, wire_12386, wire_7040, wire_3188, wire_12527, wire_12465, wire_12464, wire_12425, wire_12424, wire_12398, wire_12385, wire_12384, wire_7038, wire_3188, wire_12525, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12406, wire_7036, wire_3232, wire_3188, wire_12523, wire_12459, wire_12458, wire_12419, wire_12418, wire_12414, wire_12379, wire_12378, wire_7034, wire_3232, wire_3188, wire_12521, wire_12457, wire_12456, wire_12422, wire_12417, wire_12416, wire_12377, wire_12376, wire_7032, wire_3232, wire_3188, wire_12519, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12430, wire_7030, wire_3232, wire_3184, wire_12517, wire_12451, wire_12450, wire_12438, wire_12411, wire_12410, wire_12371, wire_12370, wire_7028, wire_3232, wire_3184, wire_12515, wire_12449, wire_12448, wire_12446, wire_12409, wire_12408, wire_12369, wire_12368, wire_7026, wire_3232, wire_3184, wire_12513, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12454, wire_7024, wire_3228, wire_3184, wire_12511, wire_12462, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_7022, wire_3228, wire_3184, wire_12539, wire_12470, wire_12441, wire_12440, wire_12401, wire_12400, wire_12361, wire_12360, wire_7020, wire_3228, wire_3184, wire_12903, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12854, wire_7199, wire_3228, wire_12905, wire_12867, wire_12866, wire_12846, wire_12827, wire_12826, wire_12787, wire_12786, wire_7197, wire_3228, wire_12907, wire_12865, wire_12864, wire_12838, wire_12825, wire_12824, wire_12785, wire_12784, wire_7195, wire_3228, wire_12909, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12830, wire_7193, wire_3188, wire_12911, wire_12859, wire_12858, wire_12822, wire_12819, wire_12818, wire_12779, wire_12778, wire_7191, wire_3188, wire_12913, wire_12857, wire_12856, wire_12817, wire_12816, wire_12814, wire_12777, wire_12776, wire_7189, wire_3188, wire_12915, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12806, wire_7187, wire_3232, wire_3188, wire_12917, wire_12851, wire_12850, wire_12811, wire_12810, wire_12798, wire_12771, wire_12770, wire_7185, wire_3232, wire_3188, wire_12919, wire_12849, wire_12848, wire_12809, wire_12808, wire_12790, wire_12769, wire_12768, wire_7183, wire_3232, wire_3188, wire_12921, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12782, wire_7181, wire_3232, wire_3184, wire_12923, wire_12843, wire_12842, wire_12803, wire_12802, wire_12774, wire_12763, wire_12762, wire_7179, wire_3232, wire_3184, wire_12925, wire_12841, wire_12840, wire_12801, wire_12800, wire_12766, wire_12761, wire_12760, wire_7177, wire_3232, wire_3184, wire_12927, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12758, wire_7175, wire_3228, wire_3184, wire_12929, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_12750, wire_7173, wire_3228, wire_3184, wire_12901, wire_12862, wire_12833, wire_12832, wire_12793, wire_12792, wire_12753, wire_12752, wire_7171, wire_3228, wire_3184};
    // CHNAXY TOTAL: 636
    assign wire_7051 = lut_tile_2_6_chanxy_out[0];
    assign wire_7053 = lut_tile_2_6_chanxy_out[1];
    assign wire_7055 = lut_tile_2_6_chanxy_out[2];
    assign wire_7057 = lut_tile_2_6_chanxy_out[3];
    assign wire_7059 = lut_tile_2_6_chanxy_out[4];
    assign wire_7061 = lut_tile_2_6_chanxy_out[5];
    assign wire_7063 = lut_tile_2_6_chanxy_out[6];
    assign wire_7065 = lut_tile_2_6_chanxy_out[7];
    assign wire_7067 = lut_tile_2_6_chanxy_out[8];
    assign wire_7069 = lut_tile_2_6_chanxy_out[9];
    assign wire_7071 = lut_tile_2_6_chanxy_out[10];
    assign wire_7073 = lut_tile_2_6_chanxy_out[11];
    assign wire_7075 = lut_tile_2_6_chanxy_out[12];
    assign wire_7077 = lut_tile_2_6_chanxy_out[13];
    assign wire_7079 = lut_tile_2_6_chanxy_out[14];
    assign wire_7140 = lut_tile_2_6_chanxy_out[15];
    assign wire_7142 = lut_tile_2_6_chanxy_out[16];
    assign wire_7144 = lut_tile_2_6_chanxy_out[17];
    assign wire_7146 = lut_tile_2_6_chanxy_out[18];
    assign wire_7148 = lut_tile_2_6_chanxy_out[19];
    assign wire_7150 = lut_tile_2_6_chanxy_out[20];
    assign wire_7152 = lut_tile_2_6_chanxy_out[21];
    assign wire_7154 = lut_tile_2_6_chanxy_out[22];
    assign wire_7156 = lut_tile_2_6_chanxy_out[23];
    assign wire_7158 = lut_tile_2_6_chanxy_out[24];
    assign wire_7160 = lut_tile_2_6_chanxy_out[25];
    assign wire_7162 = lut_tile_2_6_chanxy_out[26];
    assign wire_7164 = lut_tile_2_6_chanxy_out[27];
    assign wire_7166 = lut_tile_2_6_chanxy_out[28];
    assign wire_7168 = lut_tile_2_6_chanxy_out[29];
    assign wire_12751 = lut_tile_2_6_chanxy_out[30];
    assign wire_12759 = lut_tile_2_6_chanxy_out[31];
    assign wire_12767 = lut_tile_2_6_chanxy_out[32];
    assign wire_12775 = lut_tile_2_6_chanxy_out[33];
    assign wire_12783 = lut_tile_2_6_chanxy_out[34];
    assign wire_12791 = lut_tile_2_6_chanxy_out[35];
    assign wire_12799 = lut_tile_2_6_chanxy_out[36];
    assign wire_12807 = lut_tile_2_6_chanxy_out[37];
    assign wire_12815 = lut_tile_2_6_chanxy_out[38];
    assign wire_12823 = lut_tile_2_6_chanxy_out[39];
    assign wire_12831 = lut_tile_2_6_chanxy_out[40];
    assign wire_12839 = lut_tile_2_6_chanxy_out[41];
    assign wire_12847 = lut_tile_2_6_chanxy_out[42];
    assign wire_12855 = lut_tile_2_6_chanxy_out[43];
    assign wire_12863 = lut_tile_2_6_chanxy_out[44];
    assign wire_12870 = lut_tile_2_6_chanxy_out[45];
    assign wire_12872 = lut_tile_2_6_chanxy_out[46];
    assign wire_12874 = lut_tile_2_6_chanxy_out[47];
    assign wire_12876 = lut_tile_2_6_chanxy_out[48];
    assign wire_12878 = lut_tile_2_6_chanxy_out[49];
    assign wire_12880 = lut_tile_2_6_chanxy_out[50];
    assign wire_12882 = lut_tile_2_6_chanxy_out[51];
    assign wire_12884 = lut_tile_2_6_chanxy_out[52];
    assign wire_12886 = lut_tile_2_6_chanxy_out[53];
    assign wire_12888 = lut_tile_2_6_chanxy_out[54];
    assign wire_12890 = lut_tile_2_6_chanxy_out[55];
    assign wire_12892 = lut_tile_2_6_chanxy_out[56];
    assign wire_12894 = lut_tile_2_6_chanxy_out[57];
    assign wire_12896 = lut_tile_2_6_chanxy_out[58];
    assign wire_12898 = lut_tile_2_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_7_chanxy_in = {wire_13252, wire_6811, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6692, wire_4215, wire_13244, wire_6839, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6694, wire_4215, wire_13236, wire_6837, wire_6749, wire_6748, wire_6739, wire_6738, wire_6729, wire_6728, wire_6696, wire_4215, wire_13228, wire_6835, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6698, wire_3705, wire_13220, wire_6833, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6700, wire_3705, wire_13212, wire_6831, wire_6747, wire_6746, wire_6737, wire_6736, wire_6727, wire_6726, wire_6702, wire_3705, wire_13204, wire_6829, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6704, wire_4219, wire_3705, wire_13196, wire_6827, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6706, wire_4219, wire_3705, wire_13188, wire_6825, wire_6745, wire_6744, wire_6735, wire_6734, wire_6725, wire_6724, wire_6708, wire_4219, wire_3705, wire_13180, wire_6823, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6710, wire_4219, wire_3701, wire_13172, wire_6821, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6712, wire_4219, wire_3701, wire_13164, wire_6819, wire_6743, wire_6742, wire_6733, wire_6732, wire_6723, wire_6722, wire_6714, wire_4219, wire_3701, wire_13156, wire_6817, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6716, wire_4215, wire_3701, wire_13148, wire_6815, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6718, wire_4215, wire_3701, wire_13140, wire_6813, wire_6741, wire_6740, wire_6731, wire_6730, wire_6721, wire_6720, wire_6690, wire_4215, wire_3701, wire_13319, wire_7229, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7080, wire_4215, wire_13317, wire_7201, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7108, wire_4215, wire_13315, wire_7203, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7106, wire_4215, wire_13313, wire_7205, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7104, wire_3705, wire_13311, wire_7207, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7102, wire_3705, wire_13309, wire_7209, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7100, wire_3705, wire_13307, wire_7211, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7098, wire_4219, wire_3705, wire_13305, wire_7213, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7096, wire_4219, wire_3705, wire_13303, wire_7215, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7094, wire_4219, wire_3705, wire_13301, wire_7217, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7092, wire_4219, wire_3701, wire_13299, wire_7219, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7090, wire_4219, wire_3701, wire_13297, wire_7221, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7088, wire_4219, wire_3701, wire_13295, wire_7223, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7086, wire_4215, wire_3701, wire_13293, wire_7225, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7084, wire_4215, wire_3701, wire_13291, wire_7227, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7082, wire_4215, wire_3701, wire_12927, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12862, wire_7078, wire_3744, wire_12925, wire_12867, wire_12866, wire_12827, wire_12826, wire_12787, wire_12786, wire_12750, wire_7076, wire_3744, wire_12923, wire_12865, wire_12864, wire_12825, wire_12824, wire_12785, wire_12784, wire_12758, wire_7074, wire_3744, wire_12921, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12766, wire_7072, wire_3704, wire_12919, wire_12859, wire_12858, wire_12819, wire_12818, wire_12779, wire_12778, wire_12774, wire_7070, wire_3704, wire_12917, wire_12857, wire_12856, wire_12817, wire_12816, wire_12782, wire_12777, wire_12776, wire_7068, wire_3704, wire_12915, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12790, wire_7066, wire_3748, wire_3704, wire_12913, wire_12851, wire_12850, wire_12811, wire_12810, wire_12798, wire_12771, wire_12770, wire_7064, wire_3748, wire_3704, wire_12911, wire_12849, wire_12848, wire_12809, wire_12808, wire_12806, wire_12769, wire_12768, wire_7062, wire_3748, wire_3704, wire_12909, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12814, wire_7060, wire_3748, wire_3700, wire_12907, wire_12843, wire_12842, wire_12822, wire_12803, wire_12802, wire_12763, wire_12762, wire_7058, wire_3748, wire_3700, wire_12905, wire_12841, wire_12840, wire_12830, wire_12801, wire_12800, wire_12761, wire_12760, wire_7056, wire_3748, wire_3700, wire_12903, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12838, wire_7054, wire_3744, wire_3700, wire_12901, wire_12846, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_7052, wire_3744, wire_3700, wire_12929, wire_12854, wire_12833, wire_12832, wire_12793, wire_12792, wire_12753, wire_12752, wire_7050, wire_3744, wire_3700, wire_13293, wire_13259, wire_13258, wire_13246, wire_13219, wire_13218, wire_13179, wire_13178, wire_7229, wire_3744, wire_13295, wire_13257, wire_13256, wire_13238, wire_13217, wire_13216, wire_13177, wire_13176, wire_7227, wire_3744, wire_13297, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13230, wire_7225, wire_3744, wire_13299, wire_13251, wire_13250, wire_13222, wire_13211, wire_13210, wire_13171, wire_13170, wire_7223, wire_3704, wire_13301, wire_13249, wire_13248, wire_13214, wire_13209, wire_13208, wire_13169, wire_13168, wire_7221, wire_3704, wire_13303, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13206, wire_7219, wire_3704, wire_13305, wire_13243, wire_13242, wire_13203, wire_13202, wire_13198, wire_13163, wire_13162, wire_7217, wire_3748, wire_3704, wire_13307, wire_13241, wire_13240, wire_13201, wire_13200, wire_13190, wire_13161, wire_13160, wire_7215, wire_3748, wire_3704, wire_13309, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13182, wire_7213, wire_3748, wire_3704, wire_13311, wire_13235, wire_13234, wire_13195, wire_13194, wire_13174, wire_13155, wire_13154, wire_7211, wire_3748, wire_3700, wire_13313, wire_13233, wire_13232, wire_13193, wire_13192, wire_13166, wire_13153, wire_13152, wire_7209, wire_3748, wire_3700, wire_13315, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13158, wire_7207, wire_3748, wire_3700, wire_13317, wire_13227, wire_13226, wire_13187, wire_13186, wire_13150, wire_13147, wire_13146, wire_7205, wire_3744, wire_3700, wire_13319, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_13142, wire_7203, wire_3744, wire_3700, wire_13291, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13254, wire_7201, wire_3744, wire_3700};
    // CHNAXY TOTAL: 636
    assign wire_7081 = lut_tile_2_7_chanxy_out[0];
    assign wire_7083 = lut_tile_2_7_chanxy_out[1];
    assign wire_7085 = lut_tile_2_7_chanxy_out[2];
    assign wire_7087 = lut_tile_2_7_chanxy_out[3];
    assign wire_7089 = lut_tile_2_7_chanxy_out[4];
    assign wire_7091 = lut_tile_2_7_chanxy_out[5];
    assign wire_7093 = lut_tile_2_7_chanxy_out[6];
    assign wire_7095 = lut_tile_2_7_chanxy_out[7];
    assign wire_7097 = lut_tile_2_7_chanxy_out[8];
    assign wire_7099 = lut_tile_2_7_chanxy_out[9];
    assign wire_7101 = lut_tile_2_7_chanxy_out[10];
    assign wire_7103 = lut_tile_2_7_chanxy_out[11];
    assign wire_7105 = lut_tile_2_7_chanxy_out[12];
    assign wire_7107 = lut_tile_2_7_chanxy_out[13];
    assign wire_7109 = lut_tile_2_7_chanxy_out[14];
    assign wire_7170 = lut_tile_2_7_chanxy_out[15];
    assign wire_7172 = lut_tile_2_7_chanxy_out[16];
    assign wire_7174 = lut_tile_2_7_chanxy_out[17];
    assign wire_7176 = lut_tile_2_7_chanxy_out[18];
    assign wire_7178 = lut_tile_2_7_chanxy_out[19];
    assign wire_7180 = lut_tile_2_7_chanxy_out[20];
    assign wire_7182 = lut_tile_2_7_chanxy_out[21];
    assign wire_7184 = lut_tile_2_7_chanxy_out[22];
    assign wire_7186 = lut_tile_2_7_chanxy_out[23];
    assign wire_7188 = lut_tile_2_7_chanxy_out[24];
    assign wire_7190 = lut_tile_2_7_chanxy_out[25];
    assign wire_7192 = lut_tile_2_7_chanxy_out[26];
    assign wire_7194 = lut_tile_2_7_chanxy_out[27];
    assign wire_7196 = lut_tile_2_7_chanxy_out[28];
    assign wire_7198 = lut_tile_2_7_chanxy_out[29];
    assign wire_13143 = lut_tile_2_7_chanxy_out[30];
    assign wire_13151 = lut_tile_2_7_chanxy_out[31];
    assign wire_13159 = lut_tile_2_7_chanxy_out[32];
    assign wire_13167 = lut_tile_2_7_chanxy_out[33];
    assign wire_13175 = lut_tile_2_7_chanxy_out[34];
    assign wire_13183 = lut_tile_2_7_chanxy_out[35];
    assign wire_13191 = lut_tile_2_7_chanxy_out[36];
    assign wire_13199 = lut_tile_2_7_chanxy_out[37];
    assign wire_13207 = lut_tile_2_7_chanxy_out[38];
    assign wire_13215 = lut_tile_2_7_chanxy_out[39];
    assign wire_13223 = lut_tile_2_7_chanxy_out[40];
    assign wire_13231 = lut_tile_2_7_chanxy_out[41];
    assign wire_13239 = lut_tile_2_7_chanxy_out[42];
    assign wire_13247 = lut_tile_2_7_chanxy_out[43];
    assign wire_13255 = lut_tile_2_7_chanxy_out[44];
    assign wire_13260 = lut_tile_2_7_chanxy_out[45];
    assign wire_13262 = lut_tile_2_7_chanxy_out[46];
    assign wire_13264 = lut_tile_2_7_chanxy_out[47];
    assign wire_13266 = lut_tile_2_7_chanxy_out[48];
    assign wire_13268 = lut_tile_2_7_chanxy_out[49];
    assign wire_13270 = lut_tile_2_7_chanxy_out[50];
    assign wire_13272 = lut_tile_2_7_chanxy_out[51];
    assign wire_13274 = lut_tile_2_7_chanxy_out[52];
    assign wire_13276 = lut_tile_2_7_chanxy_out[53];
    assign wire_13278 = lut_tile_2_7_chanxy_out[54];
    assign wire_13280 = lut_tile_2_7_chanxy_out[55];
    assign wire_13282 = lut_tile_2_7_chanxy_out[56];
    assign wire_13284 = lut_tile_2_7_chanxy_out[57];
    assign wire_13286 = lut_tile_2_7_chanxy_out[58];
    assign wire_13288 = lut_tile_2_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_8_chanxy_in = {wire_13644, wire_6841, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6722, wire_4731, wire_13636, wire_6869, wire_6779, wire_6778, wire_6769, wire_6768, wire_6759, wire_6758, wire_6724, wire_4731, wire_13628, wire_6867, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6726, wire_4731, wire_13620, wire_6865, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6728, wire_4221, wire_13612, wire_6863, wire_6777, wire_6776, wire_6767, wire_6766, wire_6757, wire_6756, wire_6730, wire_4221, wire_13604, wire_6861, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6732, wire_4221, wire_13596, wire_6859, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6734, wire_4735, wire_4221, wire_13588, wire_6857, wire_6775, wire_6774, wire_6765, wire_6764, wire_6755, wire_6754, wire_6736, wire_4735, wire_4221, wire_13580, wire_6855, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6738, wire_4735, wire_4221, wire_13572, wire_6853, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6740, wire_4735, wire_4217, wire_13564, wire_6851, wire_6773, wire_6772, wire_6763, wire_6762, wire_6753, wire_6752, wire_6742, wire_4735, wire_4217, wire_13556, wire_6849, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6744, wire_4735, wire_4217, wire_13548, wire_6847, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6746, wire_4731, wire_4217, wire_13540, wire_6845, wire_6771, wire_6770, wire_6761, wire_6760, wire_6751, wire_6750, wire_6748, wire_4731, wire_4217, wire_13532, wire_6843, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6720, wire_4731, wire_4217, wire_13709, wire_7259, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7110, wire_4731, wire_13707, wire_7231, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7138, wire_4731, wire_13705, wire_7233, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7136, wire_4731, wire_13703, wire_7235, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7134, wire_4221, wire_13701, wire_7237, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7132, wire_4221, wire_13699, wire_7239, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7130, wire_4221, wire_13697, wire_7241, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7128, wire_4735, wire_4221, wire_13695, wire_7243, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7126, wire_4735, wire_4221, wire_13693, wire_7245, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7124, wire_4735, wire_4221, wire_13691, wire_7247, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7122, wire_4735, wire_4217, wire_13689, wire_7249, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7120, wire_4735, wire_4217, wire_13687, wire_7251, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7118, wire_4735, wire_4217, wire_13685, wire_7253, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7116, wire_4731, wire_4217, wire_13683, wire_7255, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7114, wire_4731, wire_4217, wire_13681, wire_7257, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7112, wire_4731, wire_4217, wire_13317, wire_13259, wire_13258, wire_13254, wire_13219, wire_13218, wire_13179, wire_13178, wire_7108, wire_4260, wire_13315, wire_13257, wire_13256, wire_13217, wire_13216, wire_13177, wire_13176, wire_13142, wire_7106, wire_4260, wire_13313, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13150, wire_7104, wire_4260, wire_13311, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_13158, wire_7102, wire_4220, wire_13309, wire_13249, wire_13248, wire_13209, wire_13208, wire_13169, wire_13168, wire_13166, wire_7100, wire_4220, wire_13307, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13174, wire_7098, wire_4220, wire_13305, wire_13243, wire_13242, wire_13203, wire_13202, wire_13182, wire_13163, wire_13162, wire_7096, wire_4264, wire_4220, wire_13303, wire_13241, wire_13240, wire_13201, wire_13200, wire_13190, wire_13161, wire_13160, wire_7094, wire_4264, wire_4220, wire_13301, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13198, wire_7092, wire_4264, wire_4220, wire_13299, wire_13235, wire_13234, wire_13206, wire_13195, wire_13194, wire_13155, wire_13154, wire_7090, wire_4264, wire_4216, wire_13297, wire_13233, wire_13232, wire_13214, wire_13193, wire_13192, wire_13153, wire_13152, wire_7088, wire_4264, wire_4216, wire_13295, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13222, wire_7086, wire_4264, wire_4216, wire_13293, wire_13230, wire_13227, wire_13226, wire_13187, wire_13186, wire_13147, wire_13146, wire_7084, wire_4260, wire_4216, wire_13291, wire_13238, wire_13225, wire_13224, wire_13185, wire_13184, wire_13145, wire_13144, wire_7082, wire_4260, wire_4216, wire_13319, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13246, wire_7080, wire_4260, wire_4216, wire_13683, wire_13649, wire_13648, wire_13638, wire_13609, wire_13608, wire_13569, wire_13568, wire_7259, wire_4260, wire_13685, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13630, wire_7257, wire_4260, wire_13687, wire_13643, wire_13642, wire_13622, wire_13603, wire_13602, wire_13563, wire_13562, wire_7255, wire_4260, wire_13689, wire_13641, wire_13640, wire_13614, wire_13601, wire_13600, wire_13561, wire_13560, wire_7253, wire_4220, wire_13691, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13606, wire_7251, wire_4220, wire_13693, wire_13635, wire_13634, wire_13598, wire_13595, wire_13594, wire_13555, wire_13554, wire_7249, wire_4220, wire_13695, wire_13633, wire_13632, wire_13593, wire_13592, wire_13590, wire_13553, wire_13552, wire_7247, wire_4264, wire_4220, wire_13697, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13582, wire_7245, wire_4264, wire_4220, wire_13699, wire_13627, wire_13626, wire_13587, wire_13586, wire_13574, wire_13547, wire_13546, wire_7243, wire_4264, wire_4220, wire_13701, wire_13625, wire_13624, wire_13585, wire_13584, wire_13566, wire_13545, wire_13544, wire_7241, wire_4264, wire_4216, wire_13703, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13558, wire_7239, wire_4264, wire_4216, wire_13705, wire_13619, wire_13618, wire_13579, wire_13578, wire_13550, wire_13539, wire_13538, wire_7237, wire_4264, wire_4216, wire_13707, wire_13617, wire_13616, wire_13577, wire_13576, wire_13542, wire_13537, wire_13536, wire_7235, wire_4260, wire_4216, wire_13709, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13534, wire_7233, wire_4260, wire_4216, wire_13681, wire_13646, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7231, wire_4260, wire_4216};
    // CHNAXY TOTAL: 636
    assign wire_7111 = lut_tile_2_8_chanxy_out[0];
    assign wire_7113 = lut_tile_2_8_chanxy_out[1];
    assign wire_7115 = lut_tile_2_8_chanxy_out[2];
    assign wire_7117 = lut_tile_2_8_chanxy_out[3];
    assign wire_7119 = lut_tile_2_8_chanxy_out[4];
    assign wire_7121 = lut_tile_2_8_chanxy_out[5];
    assign wire_7123 = lut_tile_2_8_chanxy_out[6];
    assign wire_7125 = lut_tile_2_8_chanxy_out[7];
    assign wire_7127 = lut_tile_2_8_chanxy_out[8];
    assign wire_7129 = lut_tile_2_8_chanxy_out[9];
    assign wire_7131 = lut_tile_2_8_chanxy_out[10];
    assign wire_7133 = lut_tile_2_8_chanxy_out[11];
    assign wire_7135 = lut_tile_2_8_chanxy_out[12];
    assign wire_7137 = lut_tile_2_8_chanxy_out[13];
    assign wire_7139 = lut_tile_2_8_chanxy_out[14];
    assign wire_7200 = lut_tile_2_8_chanxy_out[15];
    assign wire_7202 = lut_tile_2_8_chanxy_out[16];
    assign wire_7204 = lut_tile_2_8_chanxy_out[17];
    assign wire_7206 = lut_tile_2_8_chanxy_out[18];
    assign wire_7208 = lut_tile_2_8_chanxy_out[19];
    assign wire_7210 = lut_tile_2_8_chanxy_out[20];
    assign wire_7212 = lut_tile_2_8_chanxy_out[21];
    assign wire_7214 = lut_tile_2_8_chanxy_out[22];
    assign wire_7216 = lut_tile_2_8_chanxy_out[23];
    assign wire_7218 = lut_tile_2_8_chanxy_out[24];
    assign wire_7220 = lut_tile_2_8_chanxy_out[25];
    assign wire_7222 = lut_tile_2_8_chanxy_out[26];
    assign wire_7224 = lut_tile_2_8_chanxy_out[27];
    assign wire_7226 = lut_tile_2_8_chanxy_out[28];
    assign wire_7228 = lut_tile_2_8_chanxy_out[29];
    assign wire_13535 = lut_tile_2_8_chanxy_out[30];
    assign wire_13543 = lut_tile_2_8_chanxy_out[31];
    assign wire_13551 = lut_tile_2_8_chanxy_out[32];
    assign wire_13559 = lut_tile_2_8_chanxy_out[33];
    assign wire_13567 = lut_tile_2_8_chanxy_out[34];
    assign wire_13575 = lut_tile_2_8_chanxy_out[35];
    assign wire_13583 = lut_tile_2_8_chanxy_out[36];
    assign wire_13591 = lut_tile_2_8_chanxy_out[37];
    assign wire_13599 = lut_tile_2_8_chanxy_out[38];
    assign wire_13607 = lut_tile_2_8_chanxy_out[39];
    assign wire_13615 = lut_tile_2_8_chanxy_out[40];
    assign wire_13623 = lut_tile_2_8_chanxy_out[41];
    assign wire_13631 = lut_tile_2_8_chanxy_out[42];
    assign wire_13639 = lut_tile_2_8_chanxy_out[43];
    assign wire_13647 = lut_tile_2_8_chanxy_out[44];
    assign wire_13650 = lut_tile_2_8_chanxy_out[45];
    assign wire_13652 = lut_tile_2_8_chanxy_out[46];
    assign wire_13654 = lut_tile_2_8_chanxy_out[47];
    assign wire_13656 = lut_tile_2_8_chanxy_out[48];
    assign wire_13658 = lut_tile_2_8_chanxy_out[49];
    assign wire_13660 = lut_tile_2_8_chanxy_out[50];
    assign wire_13662 = lut_tile_2_8_chanxy_out[51];
    assign wire_13664 = lut_tile_2_8_chanxy_out[52];
    assign wire_13666 = lut_tile_2_8_chanxy_out[53];
    assign wire_13668 = lut_tile_2_8_chanxy_out[54];
    assign wire_13670 = lut_tile_2_8_chanxy_out[55];
    assign wire_13672 = lut_tile_2_8_chanxy_out[56];
    assign wire_13674 = lut_tile_2_8_chanxy_out[57];
    assign wire_13676 = lut_tile_2_8_chanxy_out[58];
    assign wire_13678 = lut_tile_2_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_9_chanxy_in = {wire_14036, wire_6871, wire_6809, wire_6808, wire_6799, wire_6798, wire_6789, wire_6788, wire_6752, wire_5247, wire_14028, wire_6899, wire_6869, wire_6868, wire_6859, wire_6858, wire_6849, wire_6848, wire_6754, wire_5247, wire_14020, wire_6897, wire_6839, wire_6838, wire_6829, wire_6828, wire_6819, wire_6818, wire_6756, wire_5247, wire_14012, wire_6895, wire_6807, wire_6806, wire_6797, wire_6796, wire_6787, wire_6786, wire_6758, wire_4737, wire_14004, wire_6893, wire_6867, wire_6866, wire_6857, wire_6856, wire_6847, wire_6846, wire_6760, wire_4737, wire_13996, wire_6891, wire_6837, wire_6836, wire_6827, wire_6826, wire_6817, wire_6816, wire_6762, wire_4737, wire_13988, wire_6889, wire_6805, wire_6804, wire_6795, wire_6794, wire_6785, wire_6784, wire_6764, wire_5251, wire_4737, wire_13980, wire_6887, wire_6865, wire_6864, wire_6855, wire_6854, wire_6845, wire_6844, wire_6766, wire_5251, wire_4737, wire_13972, wire_6885, wire_6835, wire_6834, wire_6825, wire_6824, wire_6815, wire_6814, wire_6768, wire_5251, wire_4737, wire_13964, wire_6883, wire_6803, wire_6802, wire_6793, wire_6792, wire_6783, wire_6782, wire_6770, wire_5251, wire_4733, wire_13956, wire_6881, wire_6863, wire_6862, wire_6853, wire_6852, wire_6843, wire_6842, wire_6772, wire_5251, wire_4733, wire_13948, wire_6879, wire_6833, wire_6832, wire_6823, wire_6822, wire_6813, wire_6812, wire_6774, wire_5251, wire_4733, wire_13940, wire_6877, wire_6801, wire_6800, wire_6791, wire_6790, wire_6781, wire_6780, wire_6776, wire_5247, wire_4733, wire_13932, wire_6875, wire_6861, wire_6860, wire_6851, wire_6850, wire_6841, wire_6840, wire_6778, wire_5247, wire_4733, wire_13924, wire_6873, wire_6831, wire_6830, wire_6821, wire_6820, wire_6811, wire_6810, wire_6750, wire_5247, wire_4733, wire_14099, wire_7289, wire_7259, wire_7258, wire_7249, wire_7248, wire_7239, wire_7238, wire_7140, wire_5247, wire_14097, wire_7261, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7168, wire_5247, wire_14095, wire_7263, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7166, wire_5247, wire_14093, wire_7265, wire_7257, wire_7256, wire_7247, wire_7246, wire_7237, wire_7236, wire_7164, wire_4737, wire_14091, wire_7267, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7162, wire_4737, wire_14089, wire_7269, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7160, wire_4737, wire_14087, wire_7271, wire_7255, wire_7254, wire_7245, wire_7244, wire_7235, wire_7234, wire_7158, wire_5251, wire_4737, wire_14085, wire_7273, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7156, wire_5251, wire_4737, wire_14083, wire_7275, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7154, wire_5251, wire_4737, wire_14081, wire_7277, wire_7253, wire_7252, wire_7243, wire_7242, wire_7233, wire_7232, wire_7152, wire_5251, wire_4733, wire_14079, wire_7279, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7150, wire_5251, wire_4733, wire_14077, wire_7281, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7148, wire_5251, wire_4733, wire_14075, wire_7283, wire_7251, wire_7250, wire_7241, wire_7240, wire_7231, wire_7230, wire_7146, wire_5247, wire_4733, wire_14073, wire_7285, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7144, wire_5247, wire_4733, wire_14071, wire_7287, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7142, wire_5247, wire_4733, wire_13707, wire_13649, wire_13648, wire_13646, wire_13609, wire_13608, wire_13569, wire_13568, wire_7138, wire_4776, wire_13705, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13534, wire_7136, wire_4776, wire_13703, wire_13643, wire_13642, wire_13603, wire_13602, wire_13563, wire_13562, wire_13542, wire_7134, wire_4776, wire_13701, wire_13641, wire_13640, wire_13601, wire_13600, wire_13561, wire_13560, wire_13550, wire_7132, wire_4736, wire_13699, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13558, wire_7130, wire_4736, wire_13697, wire_13635, wire_13634, wire_13595, wire_13594, wire_13566, wire_13555, wire_13554, wire_7128, wire_4736, wire_13695, wire_13633, wire_13632, wire_13593, wire_13592, wire_13574, wire_13553, wire_13552, wire_7126, wire_4780, wire_4736, wire_13693, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13582, wire_7124, wire_4780, wire_4736, wire_13691, wire_13627, wire_13626, wire_13590, wire_13587, wire_13586, wire_13547, wire_13546, wire_7122, wire_4780, wire_4736, wire_13689, wire_13625, wire_13624, wire_13598, wire_13585, wire_13584, wire_13545, wire_13544, wire_7120, wire_4780, wire_4732, wire_13687, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13606, wire_7118, wire_4780, wire_4732, wire_13685, wire_13619, wire_13618, wire_13614, wire_13579, wire_13578, wire_13539, wire_13538, wire_7116, wire_4780, wire_4732, wire_13683, wire_13622, wire_13617, wire_13616, wire_13577, wire_13576, wire_13537, wire_13536, wire_7114, wire_4776, wire_4732, wire_13681, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13630, wire_7112, wire_4776, wire_4732, wire_13709, wire_13638, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7110, wire_4776, wire_4732, wire_14073, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14030, wire_7289, wire_4776, wire_14075, wire_14035, wire_14034, wire_14022, wire_13995, wire_13994, wire_13955, wire_13954, wire_7287, wire_4776, wire_14077, wire_14033, wire_14032, wire_14014, wire_13993, wire_13992, wire_13953, wire_13952, wire_7285, wire_4776, wire_14079, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_14006, wire_7283, wire_4736, wire_14081, wire_14027, wire_14026, wire_13998, wire_13987, wire_13986, wire_13947, wire_13946, wire_7281, wire_4736, wire_14083, wire_14025, wire_14024, wire_13990, wire_13985, wire_13984, wire_13945, wire_13944, wire_7279, wire_4736, wire_14085, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13982, wire_7277, wire_4780, wire_4736, wire_14087, wire_14019, wire_14018, wire_13979, wire_13978, wire_13974, wire_13939, wire_13938, wire_7275, wire_4780, wire_4736, wire_14089, wire_14017, wire_14016, wire_13977, wire_13976, wire_13966, wire_13937, wire_13936, wire_7273, wire_4780, wire_4736, wire_14091, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13958, wire_7271, wire_4780, wire_4732, wire_14093, wire_14011, wire_14010, wire_13971, wire_13970, wire_13950, wire_13931, wire_13930, wire_7269, wire_4780, wire_4732, wire_14095, wire_14009, wire_14008, wire_13969, wire_13968, wire_13942, wire_13929, wire_13928, wire_7267, wire_4780, wire_4732, wire_14097, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_13934, wire_7265, wire_4776, wire_4732, wire_14099, wire_14003, wire_14002, wire_13963, wire_13962, wire_13926, wire_13923, wire_13922, wire_7263, wire_4776, wire_4732, wire_14071, wire_14038, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_7261, wire_4776, wire_4732};
    // CHNAXY TOTAL: 636
    assign wire_7141 = lut_tile_2_9_chanxy_out[0];
    assign wire_7143 = lut_tile_2_9_chanxy_out[1];
    assign wire_7145 = lut_tile_2_9_chanxy_out[2];
    assign wire_7147 = lut_tile_2_9_chanxy_out[3];
    assign wire_7149 = lut_tile_2_9_chanxy_out[4];
    assign wire_7151 = lut_tile_2_9_chanxy_out[5];
    assign wire_7153 = lut_tile_2_9_chanxy_out[6];
    assign wire_7155 = lut_tile_2_9_chanxy_out[7];
    assign wire_7157 = lut_tile_2_9_chanxy_out[8];
    assign wire_7159 = lut_tile_2_9_chanxy_out[9];
    assign wire_7161 = lut_tile_2_9_chanxy_out[10];
    assign wire_7163 = lut_tile_2_9_chanxy_out[11];
    assign wire_7165 = lut_tile_2_9_chanxy_out[12];
    assign wire_7167 = lut_tile_2_9_chanxy_out[13];
    assign wire_7169 = lut_tile_2_9_chanxy_out[14];
    assign wire_7230 = lut_tile_2_9_chanxy_out[15];
    assign wire_7232 = lut_tile_2_9_chanxy_out[16];
    assign wire_7234 = lut_tile_2_9_chanxy_out[17];
    assign wire_7236 = lut_tile_2_9_chanxy_out[18];
    assign wire_7238 = lut_tile_2_9_chanxy_out[19];
    assign wire_7240 = lut_tile_2_9_chanxy_out[20];
    assign wire_7242 = lut_tile_2_9_chanxy_out[21];
    assign wire_7244 = lut_tile_2_9_chanxy_out[22];
    assign wire_7246 = lut_tile_2_9_chanxy_out[23];
    assign wire_7248 = lut_tile_2_9_chanxy_out[24];
    assign wire_7250 = lut_tile_2_9_chanxy_out[25];
    assign wire_7252 = lut_tile_2_9_chanxy_out[26];
    assign wire_7254 = lut_tile_2_9_chanxy_out[27];
    assign wire_7256 = lut_tile_2_9_chanxy_out[28];
    assign wire_7258 = lut_tile_2_9_chanxy_out[29];
    assign wire_13927 = lut_tile_2_9_chanxy_out[30];
    assign wire_13935 = lut_tile_2_9_chanxy_out[31];
    assign wire_13943 = lut_tile_2_9_chanxy_out[32];
    assign wire_13951 = lut_tile_2_9_chanxy_out[33];
    assign wire_13959 = lut_tile_2_9_chanxy_out[34];
    assign wire_13967 = lut_tile_2_9_chanxy_out[35];
    assign wire_13975 = lut_tile_2_9_chanxy_out[36];
    assign wire_13983 = lut_tile_2_9_chanxy_out[37];
    assign wire_13991 = lut_tile_2_9_chanxy_out[38];
    assign wire_13999 = lut_tile_2_9_chanxy_out[39];
    assign wire_14007 = lut_tile_2_9_chanxy_out[40];
    assign wire_14015 = lut_tile_2_9_chanxy_out[41];
    assign wire_14023 = lut_tile_2_9_chanxy_out[42];
    assign wire_14031 = lut_tile_2_9_chanxy_out[43];
    assign wire_14039 = lut_tile_2_9_chanxy_out[44];
    assign wire_14040 = lut_tile_2_9_chanxy_out[45];
    assign wire_14042 = lut_tile_2_9_chanxy_out[46];
    assign wire_14044 = lut_tile_2_9_chanxy_out[47];
    assign wire_14046 = lut_tile_2_9_chanxy_out[48];
    assign wire_14048 = lut_tile_2_9_chanxy_out[49];
    assign wire_14050 = lut_tile_2_9_chanxy_out[50];
    assign wire_14052 = lut_tile_2_9_chanxy_out[51];
    assign wire_14054 = lut_tile_2_9_chanxy_out[52];
    assign wire_14056 = lut_tile_2_9_chanxy_out[53];
    assign wire_14058 = lut_tile_2_9_chanxy_out[54];
    assign wire_14060 = lut_tile_2_9_chanxy_out[55];
    assign wire_14062 = lut_tile_2_9_chanxy_out[56];
    assign wire_14064 = lut_tile_2_9_chanxy_out[57];
    assign wire_14066 = lut_tile_2_9_chanxy_out[58];
    assign wire_14068 = lut_tile_2_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_2_10_chanxy_in = {wire_14428, wire_6876, wire_6854, wire_6832, wire_6808, wire_5734, wire_5728, wire_5719, wire_5713, wire_14420, wire_6898, wire_6846, wire_6824, wire_6800, wire_5734, wire_5728, wire_5719, wire_5713, wire_14412, wire_6890, wire_6868, wire_6816, wire_6792, wire_5734, wire_5728, wire_5719, wire_5713, wire_14404, wire_6882, wire_6860, wire_6838, wire_6784, wire_5734, wire_5725, wire_5719, wire_5253, wire_14396, wire_6874, wire_6852, wire_6830, wire_6806, wire_5734, wire_5725, wire_5719, wire_5253, wire_14388, wire_6896, wire_6844, wire_6822, wire_6798, wire_5734, wire_5725, wire_5719, wire_5253, wire_14380, wire_6888, wire_6866, wire_6814, wire_6790, wire_5731, wire_5725, wire_5716, wire_5253, wire_14372, wire_6880, wire_6858, wire_6836, wire_6782, wire_5731, wire_5725, wire_5716, wire_5253, wire_14364, wire_6872, wire_6850, wire_6828, wire_6804, wire_5731, wire_5725, wire_5716, wire_5253, wire_14356, wire_6894, wire_6842, wire_6820, wire_6796, wire_5731, wire_5722, wire_5716, wire_5249, wire_14348, wire_6886, wire_6864, wire_6812, wire_6788, wire_5731, wire_5722, wire_5716, wire_5249, wire_14340, wire_6878, wire_6856, wire_6834, wire_6780, wire_5731, wire_5722, wire_5716, wire_5249, wire_14332, wire_6870, wire_6848, wire_6826, wire_6802, wire_5728, wire_5722, wire_5713, wire_5249, wire_14324, wire_6892, wire_6840, wire_6818, wire_6794, wire_5728, wire_5722, wire_5713, wire_5249, wire_14316, wire_6884, wire_6862, wire_6810, wire_6786, wire_5728, wire_5722, wire_5713, wire_5249, wire_14489, wire_7288, wire_7236, wire_7214, wire_7192, wire_5734, wire_5728, wire_5719, wire_5713, wire_14487, wire_7280, wire_7258, wire_7206, wire_7184, wire_5734, wire_5728, wire_5719, wire_5713, wire_14485, wire_7272, wire_7250, wire_7228, wire_7176, wire_5734, wire_5728, wire_5719, wire_5713, wire_14483, wire_7264, wire_7242, wire_7220, wire_7198, wire_5734, wire_5725, wire_5719, wire_5253, wire_14481, wire_7286, wire_7234, wire_7212, wire_7190, wire_5734, wire_5725, wire_5719, wire_5253, wire_14479, wire_7278, wire_7256, wire_7204, wire_7182, wire_5734, wire_5725, wire_5719, wire_5253, wire_14477, wire_7270, wire_7248, wire_7226, wire_7174, wire_5731, wire_5725, wire_5716, wire_5253, wire_14475, wire_7262, wire_7240, wire_7218, wire_7196, wire_5731, wire_5725, wire_5716, wire_5253, wire_14473, wire_7284, wire_7232, wire_7210, wire_7188, wire_5731, wire_5725, wire_5716, wire_5253, wire_14471, wire_7276, wire_7254, wire_7202, wire_7180, wire_5731, wire_5722, wire_5716, wire_5249, wire_14469, wire_7268, wire_7246, wire_7224, wire_7172, wire_5731, wire_5722, wire_5716, wire_5249, wire_14467, wire_7260, wire_7238, wire_7216, wire_7194, wire_5731, wire_5722, wire_5716, wire_5249, wire_14465, wire_7282, wire_7230, wire_7208, wire_7186, wire_5728, wire_5722, wire_5713, wire_5249, wire_14463, wire_7274, wire_7252, wire_7200, wire_7178, wire_5728, wire_5722, wire_5713, wire_5249, wire_14461, wire_7266, wire_7244, wire_7222, wire_7170, wire_5728, wire_5722, wire_5713, wire_5249, wire_14459, wire_14458, wire_14097, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14038, wire_7168, wire_5292, wire_14489, wire_14422, wire_14095, wire_14035, wire_14034, wire_13995, wire_13994, wire_13955, wire_13954, wire_13926, wire_7166, wire_5292, wire_14361, wire_14360, wire_14093, wire_14033, wire_14032, wire_13993, wire_13992, wire_13953, wire_13952, wire_13934, wire_7164, wire_5292, wire_14441, wire_14440, wire_14091, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_13942, wire_7162, wire_5252, wire_14471, wire_14350, wire_14089, wire_14027, wire_14026, wire_13987, wire_13986, wire_13950, wire_13947, wire_13946, wire_7160, wire_5252, wire_14409, wire_14408, wire_14087, wire_14025, wire_14024, wire_13985, wire_13984, wire_13958, wire_13945, wire_13944, wire_7158, wire_5252, wire_14453, wire_14452, wire_14085, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13966, wire_7156, wire_5296, wire_5252, wire_14483, wire_14398, wire_14083, wire_14019, wire_14018, wire_13979, wire_13978, wire_13974, wire_13939, wire_13938, wire_7154, wire_5296, wire_5252, wire_14337, wire_14336, wire_14081, wire_14017, wire_14016, wire_13982, wire_13977, wire_13976, wire_13937, wire_13936, wire_7152, wire_5296, wire_5252, wire_14435, wire_14434, wire_5296, wire_14079, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13990, wire_7150, wire_5296, wire_5248, wire_14465, wire_14326, wire_5296, wire_14077, wire_14011, wire_14010, wire_13998, wire_13971, wire_13970, wire_13931, wire_13930, wire_7148, wire_5296, wire_5248, wire_14385, wire_14384, wire_5292, wire_14075, wire_14009, wire_14008, wire_14006, wire_13969, wire_13968, wire_13929, wire_13928, wire_7146, wire_5296, wire_5248, wire_14447, wire_14446, wire_5252, wire_14073, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_14014, wire_7144, wire_5292, wire_5248, wire_14477, wire_14374, wire_5252, wire_14071, wire_14022, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_7142, wire_5292, wire_5248, wire_14313, wire_14312, wire_5248, wire_14099, wire_14030, wire_14001, wire_14000, wire_13961, wire_13960, wire_13921, wire_13920, wire_7140, wire_5292, wire_5248, wire_14427, wire_14426, wire_14363, wire_14362, wire_14417, wire_14416, wire_14355, wire_14354, wire_14411, wire_14410, wire_14345, wire_14344, wire_14403, wire_14402, wire_14339, wire_14338, wire_14393, wire_14392, wire_14331, wire_14330, wire_5296, wire_14387, wire_14386, wire_5296, wire_14321, wire_14320, wire_5292, wire_14379, wire_14378, wire_5252, wire_14315, wire_14314, wire_5252, wire_14369, wire_14368, wire_5248, wire_14443, wire_14442, wire_14457, wire_14456, wire_14487, wire_14414, wire_14455, wire_14454, wire_14439, wire_14438, wire_14469, wire_14342, wire_14437, wire_14436, wire_14451, wire_14450, wire_14481, wire_14390, wire_14449, wire_14448, wire_5296, wire_14433, wire_14432, wire_5292, wire_14463, wire_14318, wire_5292, wire_14431, wire_14430, wire_5252, wire_14445, wire_14444, wire_5248, wire_14475, wire_14366, wire_5248, wire_14425, wire_14424, wire_14419, wire_14418, wire_14473, wire_14358, wire_14353, wire_14352, wire_14347, wire_14346, wire_14485, wire_14406, wire_14401, wire_14400, wire_14395, wire_14394, wire_14467, wire_14334, wire_14329, wire_14328, wire_5296, wire_14323, wire_14322, wire_5292, wire_14479, wire_14382, wire_5292, wire_14377, wire_14376, wire_5252, wire_14371, wire_14370, wire_5248, wire_14461, wire_14310, wire_5248};
    // CHNAXY TOTAL: 573
    assign wire_7171 = lut_tile_2_10_chanxy_out[0];
    assign wire_7173 = lut_tile_2_10_chanxy_out[1];
    assign wire_7175 = lut_tile_2_10_chanxy_out[2];
    assign wire_7177 = lut_tile_2_10_chanxy_out[3];
    assign wire_7179 = lut_tile_2_10_chanxy_out[4];
    assign wire_7181 = lut_tile_2_10_chanxy_out[5];
    assign wire_7183 = lut_tile_2_10_chanxy_out[6];
    assign wire_7185 = lut_tile_2_10_chanxy_out[7];
    assign wire_7187 = lut_tile_2_10_chanxy_out[8];
    assign wire_7189 = lut_tile_2_10_chanxy_out[9];
    assign wire_7191 = lut_tile_2_10_chanxy_out[10];
    assign wire_7193 = lut_tile_2_10_chanxy_out[11];
    assign wire_7195 = lut_tile_2_10_chanxy_out[12];
    assign wire_7197 = lut_tile_2_10_chanxy_out[13];
    assign wire_7199 = lut_tile_2_10_chanxy_out[14];
    assign wire_7201 = lut_tile_2_10_chanxy_out[15];
    assign wire_7203 = lut_tile_2_10_chanxy_out[16];
    assign wire_7205 = lut_tile_2_10_chanxy_out[17];
    assign wire_7207 = lut_tile_2_10_chanxy_out[18];
    assign wire_7209 = lut_tile_2_10_chanxy_out[19];
    assign wire_7211 = lut_tile_2_10_chanxy_out[20];
    assign wire_7213 = lut_tile_2_10_chanxy_out[21];
    assign wire_7215 = lut_tile_2_10_chanxy_out[22];
    assign wire_7217 = lut_tile_2_10_chanxy_out[23];
    assign wire_7219 = lut_tile_2_10_chanxy_out[24];
    assign wire_7221 = lut_tile_2_10_chanxy_out[25];
    assign wire_7223 = lut_tile_2_10_chanxy_out[26];
    assign wire_7225 = lut_tile_2_10_chanxy_out[27];
    assign wire_7227 = lut_tile_2_10_chanxy_out[28];
    assign wire_7229 = lut_tile_2_10_chanxy_out[29];
    assign wire_7231 = lut_tile_2_10_chanxy_out[30];
    assign wire_7233 = lut_tile_2_10_chanxy_out[31];
    assign wire_7235 = lut_tile_2_10_chanxy_out[32];
    assign wire_7237 = lut_tile_2_10_chanxy_out[33];
    assign wire_7239 = lut_tile_2_10_chanxy_out[34];
    assign wire_7241 = lut_tile_2_10_chanxy_out[35];
    assign wire_7243 = lut_tile_2_10_chanxy_out[36];
    assign wire_7245 = lut_tile_2_10_chanxy_out[37];
    assign wire_7247 = lut_tile_2_10_chanxy_out[38];
    assign wire_7249 = lut_tile_2_10_chanxy_out[39];
    assign wire_7251 = lut_tile_2_10_chanxy_out[40];
    assign wire_7253 = lut_tile_2_10_chanxy_out[41];
    assign wire_7255 = lut_tile_2_10_chanxy_out[42];
    assign wire_7257 = lut_tile_2_10_chanxy_out[43];
    assign wire_7259 = lut_tile_2_10_chanxy_out[44];
    assign wire_7260 = lut_tile_2_10_chanxy_out[45];
    assign wire_7261 = lut_tile_2_10_chanxy_out[46];
    assign wire_7262 = lut_tile_2_10_chanxy_out[47];
    assign wire_7263 = lut_tile_2_10_chanxy_out[48];
    assign wire_7264 = lut_tile_2_10_chanxy_out[49];
    assign wire_7265 = lut_tile_2_10_chanxy_out[50];
    assign wire_7266 = lut_tile_2_10_chanxy_out[51];
    assign wire_7267 = lut_tile_2_10_chanxy_out[52];
    assign wire_7268 = lut_tile_2_10_chanxy_out[53];
    assign wire_7269 = lut_tile_2_10_chanxy_out[54];
    assign wire_7270 = lut_tile_2_10_chanxy_out[55];
    assign wire_7271 = lut_tile_2_10_chanxy_out[56];
    assign wire_7272 = lut_tile_2_10_chanxy_out[57];
    assign wire_7273 = lut_tile_2_10_chanxy_out[58];
    assign wire_7274 = lut_tile_2_10_chanxy_out[59];
    assign wire_7275 = lut_tile_2_10_chanxy_out[60];
    assign wire_7276 = lut_tile_2_10_chanxy_out[61];
    assign wire_7277 = lut_tile_2_10_chanxy_out[62];
    assign wire_7278 = lut_tile_2_10_chanxy_out[63];
    assign wire_7279 = lut_tile_2_10_chanxy_out[64];
    assign wire_7280 = lut_tile_2_10_chanxy_out[65];
    assign wire_7281 = lut_tile_2_10_chanxy_out[66];
    assign wire_7282 = lut_tile_2_10_chanxy_out[67];
    assign wire_7283 = lut_tile_2_10_chanxy_out[68];
    assign wire_7284 = lut_tile_2_10_chanxy_out[69];
    assign wire_7285 = lut_tile_2_10_chanxy_out[70];
    assign wire_7286 = lut_tile_2_10_chanxy_out[71];
    assign wire_7287 = lut_tile_2_10_chanxy_out[72];
    assign wire_7288 = lut_tile_2_10_chanxy_out[73];
    assign wire_7289 = lut_tile_2_10_chanxy_out[74];
    assign wire_14311 = lut_tile_2_10_chanxy_out[75];
    assign wire_14319 = lut_tile_2_10_chanxy_out[76];
    assign wire_14327 = lut_tile_2_10_chanxy_out[77];
    assign wire_14335 = lut_tile_2_10_chanxy_out[78];
    assign wire_14343 = lut_tile_2_10_chanxy_out[79];
    assign wire_14351 = lut_tile_2_10_chanxy_out[80];
    assign wire_14359 = lut_tile_2_10_chanxy_out[81];
    assign wire_14367 = lut_tile_2_10_chanxy_out[82];
    assign wire_14375 = lut_tile_2_10_chanxy_out[83];
    assign wire_14383 = lut_tile_2_10_chanxy_out[84];
    assign wire_14391 = lut_tile_2_10_chanxy_out[85];
    assign wire_14399 = lut_tile_2_10_chanxy_out[86];
    assign wire_14407 = lut_tile_2_10_chanxy_out[87];
    assign wire_14415 = lut_tile_2_10_chanxy_out[88];
    assign wire_14423 = lut_tile_2_10_chanxy_out[89];
    assign wire_14430 = lut_tile_2_10_chanxy_out[90];
    assign wire_14432 = lut_tile_2_10_chanxy_out[91];
    assign wire_14434 = lut_tile_2_10_chanxy_out[92];
    assign wire_14436 = lut_tile_2_10_chanxy_out[93];
    assign wire_14438 = lut_tile_2_10_chanxy_out[94];
    assign wire_14440 = lut_tile_2_10_chanxy_out[95];
    assign wire_14442 = lut_tile_2_10_chanxy_out[96];
    assign wire_14444 = lut_tile_2_10_chanxy_out[97];
    assign wire_14446 = lut_tile_2_10_chanxy_out[98];
    assign wire_14448 = lut_tile_2_10_chanxy_out[99];
    assign wire_14450 = lut_tile_2_10_chanxy_out[100];
    assign wire_14452 = lut_tile_2_10_chanxy_out[101];
    assign wire_14454 = lut_tile_2_10_chanxy_out[102];
    assign wire_14456 = lut_tile_2_10_chanxy_out[103];
    assign wire_14458 = lut_tile_2_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_3_1_chanxy_in = {wire_10918, wire_7021, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_6914, wire_1161, wire_10910, wire_7049, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_6922, wire_1161, wire_10902, wire_7047, wire_7013, wire_7012, wire_6973, wire_6972, wire_6933, wire_6932, wire_6930, wire_1161, wire_10894, wire_7045, wire_7009, wire_7008, wire_6969, wire_6968, wire_6938, wire_6929, wire_6928, wire_651, wire_10886, wire_7043, wire_7007, wire_7006, wire_6967, wire_6966, wire_6946, wire_6927, wire_6926, wire_651, wire_10878, wire_7041, wire_7005, wire_7004, wire_6965, wire_6964, wire_6954, wire_6925, wire_6924, wire_651, wire_10870, wire_7039, wire_7001, wire_7000, wire_6962, wire_6961, wire_6960, wire_6921, wire_6920, wire_1165, wire_651, wire_10862, wire_7037, wire_6999, wire_6998, wire_6970, wire_6959, wire_6958, wire_6919, wire_6918, wire_1165, wire_651, wire_10854, wire_7035, wire_6997, wire_6996, wire_6978, wire_6957, wire_6956, wire_6917, wire_6916, wire_1165, wire_651, wire_10846, wire_7033, wire_6993, wire_6992, wire_6986, wire_6953, wire_6952, wire_6913, wire_6912, wire_1165, wire_647, wire_10838, wire_7031, wire_6994, wire_6991, wire_6990, wire_6951, wire_6950, wire_6911, wire_6910, wire_1165, wire_647, wire_10830, wire_7029, wire_7002, wire_6989, wire_6988, wire_6949, wire_6948, wire_6909, wire_6908, wire_1165, wire_647, wire_10822, wire_7027, wire_7010, wire_6985, wire_6984, wire_6945, wire_6944, wire_6905, wire_6904, wire_1161, wire_647, wire_10814, wire_7025, wire_7018, wire_6983, wire_6982, wire_6943, wire_6942, wire_6903, wire_6902, wire_1161, wire_647, wire_10806, wire_7023, wire_6981, wire_6980, wire_6941, wire_6940, wire_6906, wire_6901, wire_6900, wire_1161, wire_647, wire_11009, wire_7439, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7290, wire_1161, wire_11007, wire_7411, wire_7407, wire_7406, wire_7402, wire_7367, wire_7366, wire_7327, wire_7326, wire_1161, wire_11005, wire_7413, wire_7405, wire_7404, wire_7394, wire_7365, wire_7364, wire_7325, wire_7324, wire_1161, wire_11003, wire_7415, wire_7401, wire_7400, wire_7386, wire_7361, wire_7360, wire_7321, wire_7320, wire_651, wire_11001, wire_7417, wire_7399, wire_7398, wire_7378, wire_7359, wire_7358, wire_7319, wire_7318, wire_651, wire_10999, wire_7419, wire_7397, wire_7396, wire_7370, wire_7357, wire_7356, wire_7317, wire_7316, wire_651, wire_10997, wire_7421, wire_7393, wire_7392, wire_7362, wire_7353, wire_7352, wire_7313, wire_7312, wire_1165, wire_651, wire_10995, wire_7423, wire_7391, wire_7390, wire_7354, wire_7351, wire_7350, wire_7311, wire_7310, wire_1165, wire_651, wire_10993, wire_7425, wire_7389, wire_7388, wire_7349, wire_7348, wire_7346, wire_7309, wire_7308, wire_1165, wire_651, wire_10991, wire_7427, wire_7385, wire_7384, wire_7345, wire_7344, wire_7338, wire_7305, wire_7304, wire_1165, wire_647, wire_10989, wire_7429, wire_7383, wire_7382, wire_7343, wire_7342, wire_7330, wire_7303, wire_7302, wire_1165, wire_647, wire_10987, wire_7431, wire_7381, wire_7380, wire_7341, wire_7340, wire_7322, wire_7301, wire_7300, wire_1165, wire_647, wire_10985, wire_7433, wire_7377, wire_7376, wire_7337, wire_7336, wire_7314, wire_7297, wire_7296, wire_1161, wire_647, wire_10983, wire_7435, wire_7375, wire_7374, wire_7335, wire_7334, wire_7306, wire_7295, wire_7294, wire_1161, wire_647, wire_10981, wire_7437, wire_7373, wire_7372, wire_7333, wire_7332, wire_7298, wire_7293, wire_7292, wire_1161, wire_647, wire_10603, wire_10464, wire_10619, wire_10528, wire_10589, wire_10588, wire_10983, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10904, wire_7439, wire_690, wire_10573, wire_10572, wire_10559, wire_10558, wire_10523, wire_10522, wire_10543, wire_10542, wire_10985, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10896, wire_7437, wire_690, wire_10617, wire_10520, wire_10587, wire_10586, wire_10459, wire_10458, wire_10557, wire_10556, wire_10987, wire_10915, wire_10914, wire_10888, wire_10875, wire_10874, wire_10835, wire_10834, wire_7435, wire_690, wire_10515, wire_10514, wire_10615, wire_10512, wire_10601, wire_10456, wire_10571, wire_10570, wire_10989, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10880, wire_7433, wire_650, wire_10585, wire_10584, wire_10541, wire_10540, wire_10451, wire_10450, wire_10555, wire_10554, wire_10991, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10872, wire_7431, wire_650, wire_10599, wire_10448, wire_10569, wire_10568, wire_10507, wire_10506, wire_10539, wire_10538, wire_10993, wire_10907, wire_10906, wire_10867, wire_10866, wire_10864, wire_10827, wire_10826, wire_7429, wire_650, wire_10443, wire_10442, wire_10597, wire_10440, wire_10613, wire_10504, wire_10583, wire_10582, wire_10995, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10856, wire_7427, wire_694, wire_650, wire_10567, wire_10566, wire_10553, wire_10552, wire_10499, wire_10498, wire_10537, wire_10536, wire_10997, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10848, wire_7425, wire_694, wire_650, wire_10611, wire_10496, wire_10581, wire_10580, wire_10435, wire_10434, wire_10551, wire_10550, wire_10999, wire_10899, wire_10898, wire_10859, wire_10858, wire_10840, wire_10819, wire_10818, wire_7423, wire_694, wire_650, wire_10491, wire_10490, wire_10609, wire_10488, wire_694, wire_10595, wire_10432, wire_694, wire_10565, wire_10564, wire_694, wire_11001, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10832, wire_7421, wire_694, wire_646, wire_10579, wire_10578, wire_694, wire_10535, wire_10534, wire_694, wire_10427, wire_10426, wire_694, wire_10549, wire_10548, wire_690, wire_11003, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10824, wire_7419, wire_694, wire_646, wire_10593, wire_10424, wire_690, wire_10563, wire_10562, wire_690, wire_10483, wire_10482, wire_690, wire_10533, wire_10532, wire_690, wire_11005, wire_10891, wire_10890, wire_10851, wire_10850, wire_10816, wire_10811, wire_10810, wire_7417, wire_694, wire_646, wire_10419, wire_10418, wire_690, wire_10591, wire_10416, wire_650, wire_10607, wire_10480, wire_650, wire_10577, wire_10576, wire_650, wire_11007, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10808, wire_7415, wire_690, wire_646, wire_10561, wire_10560, wire_650, wire_10547, wire_10546, wire_650, wire_10475, wire_10474, wire_650, wire_10531, wire_10530, wire_646, wire_11009, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10800, wire_7413, wire_690, wire_646, wire_10605, wire_10472, wire_646, wire_10575, wire_10574, wire_646, wire_10411, wire_10410, wire_646, wire_10545, wire_10544, wire_646, wire_10981, wire_10912, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_7411, wire_690, wire_646, wire_10467, wire_10466, wire_646};
    // CHNAXY TOTAL: 621
    assign wire_7290 = lut_tile_3_1_chanxy_out[0];
    assign wire_7291 = lut_tile_3_1_chanxy_out[1];
    assign wire_7292 = lut_tile_3_1_chanxy_out[2];
    assign wire_7294 = lut_tile_3_1_chanxy_out[3];
    assign wire_7296 = lut_tile_3_1_chanxy_out[4];
    assign wire_7298 = lut_tile_3_1_chanxy_out[5];
    assign wire_7299 = lut_tile_3_1_chanxy_out[6];
    assign wire_7300 = lut_tile_3_1_chanxy_out[7];
    assign wire_7302 = lut_tile_3_1_chanxy_out[8];
    assign wire_7304 = lut_tile_3_1_chanxy_out[9];
    assign wire_7306 = lut_tile_3_1_chanxy_out[10];
    assign wire_7307 = lut_tile_3_1_chanxy_out[11];
    assign wire_7308 = lut_tile_3_1_chanxy_out[12];
    assign wire_7310 = lut_tile_3_1_chanxy_out[13];
    assign wire_7312 = lut_tile_3_1_chanxy_out[14];
    assign wire_7314 = lut_tile_3_1_chanxy_out[15];
    assign wire_7315 = lut_tile_3_1_chanxy_out[16];
    assign wire_7316 = lut_tile_3_1_chanxy_out[17];
    assign wire_7318 = lut_tile_3_1_chanxy_out[18];
    assign wire_7320 = lut_tile_3_1_chanxy_out[19];
    assign wire_7322 = lut_tile_3_1_chanxy_out[20];
    assign wire_7323 = lut_tile_3_1_chanxy_out[21];
    assign wire_7324 = lut_tile_3_1_chanxy_out[22];
    assign wire_7326 = lut_tile_3_1_chanxy_out[23];
    assign wire_7328 = lut_tile_3_1_chanxy_out[24];
    assign wire_7330 = lut_tile_3_1_chanxy_out[25];
    assign wire_7331 = lut_tile_3_1_chanxy_out[26];
    assign wire_7332 = lut_tile_3_1_chanxy_out[27];
    assign wire_7334 = lut_tile_3_1_chanxy_out[28];
    assign wire_7336 = lut_tile_3_1_chanxy_out[29];
    assign wire_7338 = lut_tile_3_1_chanxy_out[30];
    assign wire_7339 = lut_tile_3_1_chanxy_out[31];
    assign wire_7340 = lut_tile_3_1_chanxy_out[32];
    assign wire_7342 = lut_tile_3_1_chanxy_out[33];
    assign wire_7344 = lut_tile_3_1_chanxy_out[34];
    assign wire_7346 = lut_tile_3_1_chanxy_out[35];
    assign wire_7347 = lut_tile_3_1_chanxy_out[36];
    assign wire_7348 = lut_tile_3_1_chanxy_out[37];
    assign wire_7350 = lut_tile_3_1_chanxy_out[38];
    assign wire_7352 = lut_tile_3_1_chanxy_out[39];
    assign wire_7354 = lut_tile_3_1_chanxy_out[40];
    assign wire_7355 = lut_tile_3_1_chanxy_out[41];
    assign wire_7356 = lut_tile_3_1_chanxy_out[42];
    assign wire_7358 = lut_tile_3_1_chanxy_out[43];
    assign wire_7360 = lut_tile_3_1_chanxy_out[44];
    assign wire_7362 = lut_tile_3_1_chanxy_out[45];
    assign wire_7363 = lut_tile_3_1_chanxy_out[46];
    assign wire_7364 = lut_tile_3_1_chanxy_out[47];
    assign wire_7366 = lut_tile_3_1_chanxy_out[48];
    assign wire_7368 = lut_tile_3_1_chanxy_out[49];
    assign wire_7370 = lut_tile_3_1_chanxy_out[50];
    assign wire_7371 = lut_tile_3_1_chanxy_out[51];
    assign wire_7372 = lut_tile_3_1_chanxy_out[52];
    assign wire_7374 = lut_tile_3_1_chanxy_out[53];
    assign wire_7376 = lut_tile_3_1_chanxy_out[54];
    assign wire_7378 = lut_tile_3_1_chanxy_out[55];
    assign wire_7379 = lut_tile_3_1_chanxy_out[56];
    assign wire_7380 = lut_tile_3_1_chanxy_out[57];
    assign wire_7382 = lut_tile_3_1_chanxy_out[58];
    assign wire_7384 = lut_tile_3_1_chanxy_out[59];
    assign wire_7386 = lut_tile_3_1_chanxy_out[60];
    assign wire_7387 = lut_tile_3_1_chanxy_out[61];
    assign wire_7388 = lut_tile_3_1_chanxy_out[62];
    assign wire_7390 = lut_tile_3_1_chanxy_out[63];
    assign wire_7392 = lut_tile_3_1_chanxy_out[64];
    assign wire_7394 = lut_tile_3_1_chanxy_out[65];
    assign wire_7395 = lut_tile_3_1_chanxy_out[66];
    assign wire_7396 = lut_tile_3_1_chanxy_out[67];
    assign wire_7398 = lut_tile_3_1_chanxy_out[68];
    assign wire_7400 = lut_tile_3_1_chanxy_out[69];
    assign wire_7402 = lut_tile_3_1_chanxy_out[70];
    assign wire_7403 = lut_tile_3_1_chanxy_out[71];
    assign wire_7404 = lut_tile_3_1_chanxy_out[72];
    assign wire_7406 = lut_tile_3_1_chanxy_out[73];
    assign wire_7408 = lut_tile_3_1_chanxy_out[74];
    assign wire_10801 = lut_tile_3_1_chanxy_out[75];
    assign wire_10809 = lut_tile_3_1_chanxy_out[76];
    assign wire_10817 = lut_tile_3_1_chanxy_out[77];
    assign wire_10825 = lut_tile_3_1_chanxy_out[78];
    assign wire_10833 = lut_tile_3_1_chanxy_out[79];
    assign wire_10841 = lut_tile_3_1_chanxy_out[80];
    assign wire_10849 = lut_tile_3_1_chanxy_out[81];
    assign wire_10857 = lut_tile_3_1_chanxy_out[82];
    assign wire_10865 = lut_tile_3_1_chanxy_out[83];
    assign wire_10873 = lut_tile_3_1_chanxy_out[84];
    assign wire_10881 = lut_tile_3_1_chanxy_out[85];
    assign wire_10889 = lut_tile_3_1_chanxy_out[86];
    assign wire_10897 = lut_tile_3_1_chanxy_out[87];
    assign wire_10905 = lut_tile_3_1_chanxy_out[88];
    assign wire_10913 = lut_tile_3_1_chanxy_out[89];
    assign wire_10950 = lut_tile_3_1_chanxy_out[90];
    assign wire_10952 = lut_tile_3_1_chanxy_out[91];
    assign wire_10954 = lut_tile_3_1_chanxy_out[92];
    assign wire_10956 = lut_tile_3_1_chanxy_out[93];
    assign wire_10958 = lut_tile_3_1_chanxy_out[94];
    assign wire_10960 = lut_tile_3_1_chanxy_out[95];
    assign wire_10962 = lut_tile_3_1_chanxy_out[96];
    assign wire_10964 = lut_tile_3_1_chanxy_out[97];
    assign wire_10966 = lut_tile_3_1_chanxy_out[98];
    assign wire_10968 = lut_tile_3_1_chanxy_out[99];
    assign wire_10970 = lut_tile_3_1_chanxy_out[100];
    assign wire_10972 = lut_tile_3_1_chanxy_out[101];
    assign wire_10974 = lut_tile_3_1_chanxy_out[102];
    assign wire_10976 = lut_tile_3_1_chanxy_out[103];
    assign wire_10978 = lut_tile_3_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_3_2_chanxy_in = {wire_11302, wire_7051, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6908, wire_1677, wire_11294, wire_7079, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_6916, wire_1677, wire_11286, wire_7077, wire_7015, wire_7014, wire_6975, wire_6974, wire_6935, wire_6934, wire_6924, wire_1677, wire_11278, wire_7075, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6932, wire_1167, wire_11270, wire_7073, wire_7009, wire_7008, wire_6969, wire_6968, wire_6940, wire_6929, wire_6928, wire_1167, wire_11262, wire_7071, wire_7007, wire_7006, wire_6967, wire_6966, wire_6948, wire_6927, wire_6926, wire_1167, wire_11254, wire_7069, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6956, wire_1681, wire_1167, wire_11246, wire_7067, wire_7001, wire_7000, wire_6964, wire_6961, wire_6960, wire_6921, wire_6920, wire_1681, wire_1167, wire_11238, wire_7065, wire_6999, wire_6998, wire_6972, wire_6959, wire_6958, wire_6919, wire_6918, wire_1681, wire_1167, wire_11230, wire_7063, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6980, wire_1681, wire_1163, wire_11222, wire_7061, wire_6993, wire_6992, wire_6988, wire_6953, wire_6952, wire_6913, wire_6912, wire_1681, wire_1163, wire_11214, wire_7059, wire_6996, wire_6991, wire_6990, wire_6951, wire_6950, wire_6911, wire_6910, wire_1681, wire_1163, wire_11206, wire_7057, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_7004, wire_1677, wire_1163, wire_11198, wire_7055, wire_7012, wire_6985, wire_6984, wire_6945, wire_6944, wire_6905, wire_6904, wire_1677, wire_1163, wire_11190, wire_7053, wire_6983, wire_6982, wire_6943, wire_6942, wire_6903, wire_6902, wire_6900, wire_1677, wire_1163, wire_11399, wire_7469, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7292, wire_1677, wire_11397, wire_7441, wire_7407, wire_7406, wire_7404, wire_7367, wire_7366, wire_7327, wire_7326, wire_1677, wire_11395, wire_7443, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7396, wire_1677, wire_11393, wire_7445, wire_7401, wire_7400, wire_7388, wire_7361, wire_7360, wire_7321, wire_7320, wire_1167, wire_11391, wire_7447, wire_7399, wire_7398, wire_7380, wire_7359, wire_7358, wire_7319, wire_7318, wire_1167, wire_11389, wire_7449, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7372, wire_1167, wire_11387, wire_7451, wire_7393, wire_7392, wire_7364, wire_7353, wire_7352, wire_7313, wire_7312, wire_1681, wire_1167, wire_11385, wire_7453, wire_7391, wire_7390, wire_7356, wire_7351, wire_7350, wire_7311, wire_7310, wire_1681, wire_1167, wire_11383, wire_7455, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7348, wire_1681, wire_1167, wire_11381, wire_7457, wire_7385, wire_7384, wire_7345, wire_7344, wire_7340, wire_7305, wire_7304, wire_1681, wire_1163, wire_11379, wire_7459, wire_7383, wire_7382, wire_7343, wire_7342, wire_7332, wire_7303, wire_7302, wire_1681, wire_1163, wire_11377, wire_7461, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7324, wire_1681, wire_1163, wire_11375, wire_7463, wire_7377, wire_7376, wire_7337, wire_7336, wire_7316, wire_7297, wire_7296, wire_1677, wire_1163, wire_11373, wire_7465, wire_7375, wire_7374, wire_7335, wire_7334, wire_7308, wire_7295, wire_7294, wire_1677, wire_1163, wire_11371, wire_7467, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7300, wire_1677, wire_1163, wire_11007, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10912, wire_7402, wire_1206, wire_11005, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10800, wire_7394, wire_1206, wire_11003, wire_10915, wire_10914, wire_10875, wire_10874, wire_10835, wire_10834, wire_10808, wire_7386, wire_1206, wire_11001, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10816, wire_7378, wire_1166, wire_10999, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10824, wire_7370, wire_1166, wire_10997, wire_10907, wire_10906, wire_10867, wire_10866, wire_10832, wire_10827, wire_10826, wire_7362, wire_1166, wire_10995, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10840, wire_7354, wire_1210, wire_1166, wire_10993, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10848, wire_7346, wire_1210, wire_1166, wire_10991, wire_10899, wire_10898, wire_10859, wire_10858, wire_10856, wire_10819, wire_10818, wire_7338, wire_1210, wire_1166, wire_10989, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10864, wire_7330, wire_1210, wire_1162, wire_10987, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10872, wire_7322, wire_1210, wire_1162, wire_10985, wire_10891, wire_10890, wire_10880, wire_10851, wire_10850, wire_10811, wire_10810, wire_7314, wire_1210, wire_1162, wire_10983, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10888, wire_7306, wire_1206, wire_1162, wire_10981, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10896, wire_7298, wire_1206, wire_1162, wire_11009, wire_10904, wire_10883, wire_10882, wire_10843, wire_10842, wire_10803, wire_10802, wire_7290, wire_1206, wire_1162, wire_11373, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11296, wire_7469, wire_1206, wire_11375, wire_11307, wire_11306, wire_11288, wire_11267, wire_11266, wire_11227, wire_11226, wire_7467, wire_1206, wire_11377, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11280, wire_7465, wire_1206, wire_11379, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11272, wire_7463, wire_1166, wire_11381, wire_11299, wire_11298, wire_11264, wire_11259, wire_11258, wire_11219, wire_11218, wire_7461, wire_1166, wire_11383, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11256, wire_7459, wire_1166, wire_11385, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11248, wire_7457, wire_1210, wire_1166, wire_11387, wire_11291, wire_11290, wire_11251, wire_11250, wire_11240, wire_11211, wire_11210, wire_7455, wire_1210, wire_1166, wire_11389, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11232, wire_7453, wire_1210, wire_1166, wire_11391, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11224, wire_7451, wire_1210, wire_1162, wire_11393, wire_11283, wire_11282, wire_11243, wire_11242, wire_11216, wire_11203, wire_11202, wire_7449, wire_1210, wire_1162, wire_11395, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11208, wire_7447, wire_1210, wire_1162, wire_11397, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11200, wire_7445, wire_1206, wire_1162, wire_11399, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_11192, wire_7443, wire_1206, wire_1162, wire_11371, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11304, wire_7441, wire_1206, wire_1162};
    // CHNAXY TOTAL: 636
    assign wire_7293 = lut_tile_3_2_chanxy_out[0];
    assign wire_7301 = lut_tile_3_2_chanxy_out[1];
    assign wire_7309 = lut_tile_3_2_chanxy_out[2];
    assign wire_7317 = lut_tile_3_2_chanxy_out[3];
    assign wire_7325 = lut_tile_3_2_chanxy_out[4];
    assign wire_7333 = lut_tile_3_2_chanxy_out[5];
    assign wire_7341 = lut_tile_3_2_chanxy_out[6];
    assign wire_7349 = lut_tile_3_2_chanxy_out[7];
    assign wire_7357 = lut_tile_3_2_chanxy_out[8];
    assign wire_7365 = lut_tile_3_2_chanxy_out[9];
    assign wire_7373 = lut_tile_3_2_chanxy_out[10];
    assign wire_7381 = lut_tile_3_2_chanxy_out[11];
    assign wire_7389 = lut_tile_3_2_chanxy_out[12];
    assign wire_7397 = lut_tile_3_2_chanxy_out[13];
    assign wire_7405 = lut_tile_3_2_chanxy_out[14];
    assign wire_7410 = lut_tile_3_2_chanxy_out[15];
    assign wire_7412 = lut_tile_3_2_chanxy_out[16];
    assign wire_7414 = lut_tile_3_2_chanxy_out[17];
    assign wire_7416 = lut_tile_3_2_chanxy_out[18];
    assign wire_7418 = lut_tile_3_2_chanxy_out[19];
    assign wire_7420 = lut_tile_3_2_chanxy_out[20];
    assign wire_7422 = lut_tile_3_2_chanxy_out[21];
    assign wire_7424 = lut_tile_3_2_chanxy_out[22];
    assign wire_7426 = lut_tile_3_2_chanxy_out[23];
    assign wire_7428 = lut_tile_3_2_chanxy_out[24];
    assign wire_7430 = lut_tile_3_2_chanxy_out[25];
    assign wire_7432 = lut_tile_3_2_chanxy_out[26];
    assign wire_7434 = lut_tile_3_2_chanxy_out[27];
    assign wire_7436 = lut_tile_3_2_chanxy_out[28];
    assign wire_7438 = lut_tile_3_2_chanxy_out[29];
    assign wire_11193 = lut_tile_3_2_chanxy_out[30];
    assign wire_11201 = lut_tile_3_2_chanxy_out[31];
    assign wire_11209 = lut_tile_3_2_chanxy_out[32];
    assign wire_11217 = lut_tile_3_2_chanxy_out[33];
    assign wire_11225 = lut_tile_3_2_chanxy_out[34];
    assign wire_11233 = lut_tile_3_2_chanxy_out[35];
    assign wire_11241 = lut_tile_3_2_chanxy_out[36];
    assign wire_11249 = lut_tile_3_2_chanxy_out[37];
    assign wire_11257 = lut_tile_3_2_chanxy_out[38];
    assign wire_11265 = lut_tile_3_2_chanxy_out[39];
    assign wire_11273 = lut_tile_3_2_chanxy_out[40];
    assign wire_11281 = lut_tile_3_2_chanxy_out[41];
    assign wire_11289 = lut_tile_3_2_chanxy_out[42];
    assign wire_11297 = lut_tile_3_2_chanxy_out[43];
    assign wire_11305 = lut_tile_3_2_chanxy_out[44];
    assign wire_11340 = lut_tile_3_2_chanxy_out[45];
    assign wire_11342 = lut_tile_3_2_chanxy_out[46];
    assign wire_11344 = lut_tile_3_2_chanxy_out[47];
    assign wire_11346 = lut_tile_3_2_chanxy_out[48];
    assign wire_11348 = lut_tile_3_2_chanxy_out[49];
    assign wire_11350 = lut_tile_3_2_chanxy_out[50];
    assign wire_11352 = lut_tile_3_2_chanxy_out[51];
    assign wire_11354 = lut_tile_3_2_chanxy_out[52];
    assign wire_11356 = lut_tile_3_2_chanxy_out[53];
    assign wire_11358 = lut_tile_3_2_chanxy_out[54];
    assign wire_11360 = lut_tile_3_2_chanxy_out[55];
    assign wire_11362 = lut_tile_3_2_chanxy_out[56];
    assign wire_11364 = lut_tile_3_2_chanxy_out[57];
    assign wire_11366 = lut_tile_3_2_chanxy_out[58];
    assign wire_11368 = lut_tile_3_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_3_chanxy_in = {wire_11694, wire_7081, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6910, wire_2193, wire_11686, wire_7109, wire_7017, wire_7016, wire_6977, wire_6976, wire_6937, wire_6936, wire_6918, wire_2193, wire_11678, wire_7107, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_6926, wire_2193, wire_11670, wire_7105, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6934, wire_1683, wire_11662, wire_7103, wire_7009, wire_7008, wire_6969, wire_6968, wire_6942, wire_6929, wire_6928, wire_1683, wire_11654, wire_7101, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6950, wire_1683, wire_11646, wire_7099, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6958, wire_2197, wire_1683, wire_11638, wire_7097, wire_7001, wire_7000, wire_6966, wire_6961, wire_6960, wire_6921, wire_6920, wire_2197, wire_1683, wire_11630, wire_7095, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_6974, wire_2197, wire_1683, wire_11622, wire_7093, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6982, wire_2197, wire_1679, wire_11614, wire_7091, wire_6993, wire_6992, wire_6990, wire_6953, wire_6952, wire_6913, wire_6912, wire_2197, wire_1679, wire_11606, wire_7089, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_6998, wire_2197, wire_1679, wire_11598, wire_7087, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_7006, wire_2193, wire_1679, wire_11590, wire_7085, wire_7014, wire_6985, wire_6984, wire_6945, wire_6944, wire_6905, wire_6904, wire_2193, wire_1679, wire_11582, wire_7083, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_6902, wire_2193, wire_1679, wire_11789, wire_7499, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7294, wire_2193, wire_11787, wire_7471, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7406, wire_2193, wire_11785, wire_7473, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7398, wire_2193, wire_11783, wire_7475, wire_7401, wire_7400, wire_7390, wire_7361, wire_7360, wire_7321, wire_7320, wire_1683, wire_11781, wire_7477, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7382, wire_1683, wire_11779, wire_7479, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7374, wire_1683, wire_11777, wire_7481, wire_7393, wire_7392, wire_7366, wire_7353, wire_7352, wire_7313, wire_7312, wire_2197, wire_1683, wire_11775, wire_7483, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7358, wire_2197, wire_1683, wire_11773, wire_7485, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7350, wire_2197, wire_1683, wire_11771, wire_7487, wire_7385, wire_7384, wire_7345, wire_7344, wire_7342, wire_7305, wire_7304, wire_2197, wire_1679, wire_11769, wire_7489, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7334, wire_2197, wire_1679, wire_11767, wire_7491, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7326, wire_2197, wire_1679, wire_11765, wire_7493, wire_7377, wire_7376, wire_7337, wire_7336, wire_7318, wire_7297, wire_7296, wire_2193, wire_1679, wire_11763, wire_7495, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7310, wire_2193, wire_1679, wire_11761, wire_7497, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7302, wire_2193, wire_1679, wire_11397, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11304, wire_7404, wire_1722, wire_11395, wire_11307, wire_11306, wire_11267, wire_11266, wire_11227, wire_11226, wire_11192, wire_7396, wire_1722, wire_11393, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11200, wire_7388, wire_1722, wire_11391, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11208, wire_7380, wire_1682, wire_11389, wire_11299, wire_11298, wire_11259, wire_11258, wire_11219, wire_11218, wire_11216, wire_7372, wire_1682, wire_11387, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11224, wire_7364, wire_1682, wire_11385, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11232, wire_7356, wire_1726, wire_1682, wire_11383, wire_11291, wire_11290, wire_11251, wire_11250, wire_11240, wire_11211, wire_11210, wire_7348, wire_1726, wire_1682, wire_11381, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11248, wire_7340, wire_1726, wire_1682, wire_11379, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11256, wire_7332, wire_1726, wire_1678, wire_11377, wire_11283, wire_11282, wire_11264, wire_11243, wire_11242, wire_11203, wire_11202, wire_7324, wire_1726, wire_1678, wire_11375, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11272, wire_7316, wire_1726, wire_1678, wire_11373, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11280, wire_7308, wire_1722, wire_1678, wire_11371, wire_11288, wire_11275, wire_11274, wire_11235, wire_11234, wire_11195, wire_11194, wire_7300, wire_1722, wire_1678, wire_11399, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11296, wire_7292, wire_1722, wire_1678, wire_11763, wire_11699, wire_11698, wire_11688, wire_11659, wire_11658, wire_11619, wire_11618, wire_7499, wire_1722, wire_11765, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11680, wire_7497, wire_1722, wire_11767, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11672, wire_7495, wire_1722, wire_11769, wire_11691, wire_11690, wire_11664, wire_11651, wire_11650, wire_11611, wire_11610, wire_7493, wire_1682, wire_11771, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11656, wire_7491, wire_1682, wire_11773, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11648, wire_7489, wire_1682, wire_11775, wire_11683, wire_11682, wire_11643, wire_11642, wire_11640, wire_11603, wire_11602, wire_7487, wire_1726, wire_1682, wire_11777, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11632, wire_7485, wire_1726, wire_1682, wire_11779, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11624, wire_7483, wire_1726, wire_1682, wire_11781, wire_11675, wire_11674, wire_11635, wire_11634, wire_11616, wire_11595, wire_11594, wire_7481, wire_1726, wire_1678, wire_11783, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11608, wire_7479, wire_1726, wire_1678, wire_11785, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11600, wire_7477, wire_1726, wire_1678, wire_11787, wire_11667, wire_11666, wire_11627, wire_11626, wire_11592, wire_11587, wire_11586, wire_7475, wire_1722, wire_1678, wire_11789, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11584, wire_7473, wire_1722, wire_1678, wire_11761, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11696, wire_7471, wire_1722, wire_1678};
    // CHNAXY TOTAL: 636
    assign wire_7295 = lut_tile_3_3_chanxy_out[0];
    assign wire_7303 = lut_tile_3_3_chanxy_out[1];
    assign wire_7311 = lut_tile_3_3_chanxy_out[2];
    assign wire_7319 = lut_tile_3_3_chanxy_out[3];
    assign wire_7327 = lut_tile_3_3_chanxy_out[4];
    assign wire_7335 = lut_tile_3_3_chanxy_out[5];
    assign wire_7343 = lut_tile_3_3_chanxy_out[6];
    assign wire_7351 = lut_tile_3_3_chanxy_out[7];
    assign wire_7359 = lut_tile_3_3_chanxy_out[8];
    assign wire_7367 = lut_tile_3_3_chanxy_out[9];
    assign wire_7375 = lut_tile_3_3_chanxy_out[10];
    assign wire_7383 = lut_tile_3_3_chanxy_out[11];
    assign wire_7391 = lut_tile_3_3_chanxy_out[12];
    assign wire_7399 = lut_tile_3_3_chanxy_out[13];
    assign wire_7407 = lut_tile_3_3_chanxy_out[14];
    assign wire_7440 = lut_tile_3_3_chanxy_out[15];
    assign wire_7442 = lut_tile_3_3_chanxy_out[16];
    assign wire_7444 = lut_tile_3_3_chanxy_out[17];
    assign wire_7446 = lut_tile_3_3_chanxy_out[18];
    assign wire_7448 = lut_tile_3_3_chanxy_out[19];
    assign wire_7450 = lut_tile_3_3_chanxy_out[20];
    assign wire_7452 = lut_tile_3_3_chanxy_out[21];
    assign wire_7454 = lut_tile_3_3_chanxy_out[22];
    assign wire_7456 = lut_tile_3_3_chanxy_out[23];
    assign wire_7458 = lut_tile_3_3_chanxy_out[24];
    assign wire_7460 = lut_tile_3_3_chanxy_out[25];
    assign wire_7462 = lut_tile_3_3_chanxy_out[26];
    assign wire_7464 = lut_tile_3_3_chanxy_out[27];
    assign wire_7466 = lut_tile_3_3_chanxy_out[28];
    assign wire_7468 = lut_tile_3_3_chanxy_out[29];
    assign wire_11585 = lut_tile_3_3_chanxy_out[30];
    assign wire_11593 = lut_tile_3_3_chanxy_out[31];
    assign wire_11601 = lut_tile_3_3_chanxy_out[32];
    assign wire_11609 = lut_tile_3_3_chanxy_out[33];
    assign wire_11617 = lut_tile_3_3_chanxy_out[34];
    assign wire_11625 = lut_tile_3_3_chanxy_out[35];
    assign wire_11633 = lut_tile_3_3_chanxy_out[36];
    assign wire_11641 = lut_tile_3_3_chanxy_out[37];
    assign wire_11649 = lut_tile_3_3_chanxy_out[38];
    assign wire_11657 = lut_tile_3_3_chanxy_out[39];
    assign wire_11665 = lut_tile_3_3_chanxy_out[40];
    assign wire_11673 = lut_tile_3_3_chanxy_out[41];
    assign wire_11681 = lut_tile_3_3_chanxy_out[42];
    assign wire_11689 = lut_tile_3_3_chanxy_out[43];
    assign wire_11697 = lut_tile_3_3_chanxy_out[44];
    assign wire_11730 = lut_tile_3_3_chanxy_out[45];
    assign wire_11732 = lut_tile_3_3_chanxy_out[46];
    assign wire_11734 = lut_tile_3_3_chanxy_out[47];
    assign wire_11736 = lut_tile_3_3_chanxy_out[48];
    assign wire_11738 = lut_tile_3_3_chanxy_out[49];
    assign wire_11740 = lut_tile_3_3_chanxy_out[50];
    assign wire_11742 = lut_tile_3_3_chanxy_out[51];
    assign wire_11744 = lut_tile_3_3_chanxy_out[52];
    assign wire_11746 = lut_tile_3_3_chanxy_out[53];
    assign wire_11748 = lut_tile_3_3_chanxy_out[54];
    assign wire_11750 = lut_tile_3_3_chanxy_out[55];
    assign wire_11752 = lut_tile_3_3_chanxy_out[56];
    assign wire_11754 = lut_tile_3_3_chanxy_out[57];
    assign wire_11756 = lut_tile_3_3_chanxy_out[58];
    assign wire_11758 = lut_tile_3_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_4_chanxy_in = {wire_12086, wire_7111, wire_7049, wire_7048, wire_7039, wire_7038, wire_7029, wire_7028, wire_6912, wire_2709, wire_12078, wire_7139, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_6920, wire_2709, wire_12070, wire_7137, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_6928, wire_2709, wire_12062, wire_7135, wire_7047, wire_7046, wire_7037, wire_7036, wire_7027, wire_7026, wire_6936, wire_2199, wire_12054, wire_7133, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_6944, wire_2199, wire_12046, wire_7131, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_6952, wire_2199, wire_12038, wire_7129, wire_7045, wire_7044, wire_7035, wire_7034, wire_7025, wire_7024, wire_6960, wire_2713, wire_2199, wire_12030, wire_7127, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_6968, wire_2713, wire_2199, wire_12022, wire_7125, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_6976, wire_2713, wire_2199, wire_12014, wire_7123, wire_7043, wire_7042, wire_7033, wire_7032, wire_7023, wire_7022, wire_6984, wire_2713, wire_2195, wire_12006, wire_7121, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_6992, wire_2713, wire_2195, wire_11998, wire_7119, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_7000, wire_2713, wire_2195, wire_11990, wire_7117, wire_7041, wire_7040, wire_7031, wire_7030, wire_7021, wire_7020, wire_7008, wire_2709, wire_2195, wire_11982, wire_7115, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7016, wire_2709, wire_2195, wire_11974, wire_7113, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_6904, wire_2709, wire_2195, wire_12179, wire_7529, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7296, wire_2709, wire_12177, wire_7501, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7408, wire_2709, wire_12175, wire_7503, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7400, wire_2709, wire_12173, wire_7505, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7392, wire_2199, wire_12171, wire_7507, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7384, wire_2199, wire_12169, wire_7509, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7376, wire_2199, wire_12167, wire_7511, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7368, wire_2713, wire_2199, wire_12165, wire_7513, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7360, wire_2713, wire_2199, wire_12163, wire_7515, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7352, wire_2713, wire_2199, wire_12161, wire_7517, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7344, wire_2713, wire_2195, wire_12159, wire_7519, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7336, wire_2713, wire_2195, wire_12157, wire_7521, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7328, wire_2713, wire_2195, wire_12155, wire_7523, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7320, wire_2709, wire_2195, wire_12153, wire_7525, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7312, wire_2709, wire_2195, wire_12151, wire_7527, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7304, wire_2709, wire_2195, wire_11787, wire_11699, wire_11698, wire_11696, wire_11659, wire_11658, wire_11619, wire_11618, wire_7406, wire_2238, wire_11785, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11584, wire_7398, wire_2238, wire_11783, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11592, wire_7390, wire_2238, wire_11781, wire_11691, wire_11690, wire_11651, wire_11650, wire_11611, wire_11610, wire_11600, wire_7382, wire_2198, wire_11779, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11608, wire_7374, wire_2198, wire_11777, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11616, wire_7366, wire_2198, wire_11775, wire_11683, wire_11682, wire_11643, wire_11642, wire_11624, wire_11603, wire_11602, wire_7358, wire_2242, wire_2198, wire_11773, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11632, wire_7350, wire_2242, wire_2198, wire_11771, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11640, wire_7342, wire_2242, wire_2198, wire_11769, wire_11675, wire_11674, wire_11648, wire_11635, wire_11634, wire_11595, wire_11594, wire_7334, wire_2242, wire_2194, wire_11767, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11656, wire_7326, wire_2242, wire_2194, wire_11765, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11664, wire_7318, wire_2242, wire_2194, wire_11763, wire_11672, wire_11667, wire_11666, wire_11627, wire_11626, wire_11587, wire_11586, wire_7310, wire_2238, wire_2194, wire_11761, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11680, wire_7302, wire_2238, wire_2194, wire_11789, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11688, wire_7294, wire_2238, wire_2194, wire_12153, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12080, wire_7529, wire_2238, wire_12155, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_12072, wire_7527, wire_2238, wire_12157, wire_12083, wire_12082, wire_12064, wire_12043, wire_12042, wire_12003, wire_12002, wire_7525, wire_2238, wire_12159, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12056, wire_7523, wire_2198, wire_12161, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12048, wire_7521, wire_2198, wire_12163, wire_12075, wire_12074, wire_12040, wire_12035, wire_12034, wire_11995, wire_11994, wire_7519, wire_2198, wire_12165, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12032, wire_7517, wire_2242, wire_2198, wire_12167, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12024, wire_7515, wire_2242, wire_2198, wire_12169, wire_12067, wire_12066, wire_12027, wire_12026, wire_12016, wire_11987, wire_11986, wire_7513, wire_2242, wire_2198, wire_12171, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12008, wire_7511, wire_2242, wire_2194, wire_12173, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12000, wire_7509, wire_2242, wire_2194, wire_12175, wire_12059, wire_12058, wire_12019, wire_12018, wire_11992, wire_11979, wire_11978, wire_7507, wire_2242, wire_2194, wire_12177, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_11984, wire_7505, wire_2238, wire_2194, wire_12179, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_11976, wire_7503, wire_2238, wire_2194, wire_12151, wire_12088, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7501, wire_2238, wire_2194};
    // CHNAXY TOTAL: 636
    assign wire_7297 = lut_tile_3_4_chanxy_out[0];
    assign wire_7305 = lut_tile_3_4_chanxy_out[1];
    assign wire_7313 = lut_tile_3_4_chanxy_out[2];
    assign wire_7321 = lut_tile_3_4_chanxy_out[3];
    assign wire_7329 = lut_tile_3_4_chanxy_out[4];
    assign wire_7337 = lut_tile_3_4_chanxy_out[5];
    assign wire_7345 = lut_tile_3_4_chanxy_out[6];
    assign wire_7353 = lut_tile_3_4_chanxy_out[7];
    assign wire_7361 = lut_tile_3_4_chanxy_out[8];
    assign wire_7369 = lut_tile_3_4_chanxy_out[9];
    assign wire_7377 = lut_tile_3_4_chanxy_out[10];
    assign wire_7385 = lut_tile_3_4_chanxy_out[11];
    assign wire_7393 = lut_tile_3_4_chanxy_out[12];
    assign wire_7401 = lut_tile_3_4_chanxy_out[13];
    assign wire_7409 = lut_tile_3_4_chanxy_out[14];
    assign wire_7470 = lut_tile_3_4_chanxy_out[15];
    assign wire_7472 = lut_tile_3_4_chanxy_out[16];
    assign wire_7474 = lut_tile_3_4_chanxy_out[17];
    assign wire_7476 = lut_tile_3_4_chanxy_out[18];
    assign wire_7478 = lut_tile_3_4_chanxy_out[19];
    assign wire_7480 = lut_tile_3_4_chanxy_out[20];
    assign wire_7482 = lut_tile_3_4_chanxy_out[21];
    assign wire_7484 = lut_tile_3_4_chanxy_out[22];
    assign wire_7486 = lut_tile_3_4_chanxy_out[23];
    assign wire_7488 = lut_tile_3_4_chanxy_out[24];
    assign wire_7490 = lut_tile_3_4_chanxy_out[25];
    assign wire_7492 = lut_tile_3_4_chanxy_out[26];
    assign wire_7494 = lut_tile_3_4_chanxy_out[27];
    assign wire_7496 = lut_tile_3_4_chanxy_out[28];
    assign wire_7498 = lut_tile_3_4_chanxy_out[29];
    assign wire_11977 = lut_tile_3_4_chanxy_out[30];
    assign wire_11985 = lut_tile_3_4_chanxy_out[31];
    assign wire_11993 = lut_tile_3_4_chanxy_out[32];
    assign wire_12001 = lut_tile_3_4_chanxy_out[33];
    assign wire_12009 = lut_tile_3_4_chanxy_out[34];
    assign wire_12017 = lut_tile_3_4_chanxy_out[35];
    assign wire_12025 = lut_tile_3_4_chanxy_out[36];
    assign wire_12033 = lut_tile_3_4_chanxy_out[37];
    assign wire_12041 = lut_tile_3_4_chanxy_out[38];
    assign wire_12049 = lut_tile_3_4_chanxy_out[39];
    assign wire_12057 = lut_tile_3_4_chanxy_out[40];
    assign wire_12065 = lut_tile_3_4_chanxy_out[41];
    assign wire_12073 = lut_tile_3_4_chanxy_out[42];
    assign wire_12081 = lut_tile_3_4_chanxy_out[43];
    assign wire_12089 = lut_tile_3_4_chanxy_out[44];
    assign wire_12120 = lut_tile_3_4_chanxy_out[45];
    assign wire_12122 = lut_tile_3_4_chanxy_out[46];
    assign wire_12124 = lut_tile_3_4_chanxy_out[47];
    assign wire_12126 = lut_tile_3_4_chanxy_out[48];
    assign wire_12128 = lut_tile_3_4_chanxy_out[49];
    assign wire_12130 = lut_tile_3_4_chanxy_out[50];
    assign wire_12132 = lut_tile_3_4_chanxy_out[51];
    assign wire_12134 = lut_tile_3_4_chanxy_out[52];
    assign wire_12136 = lut_tile_3_4_chanxy_out[53];
    assign wire_12138 = lut_tile_3_4_chanxy_out[54];
    assign wire_12140 = lut_tile_3_4_chanxy_out[55];
    assign wire_12142 = lut_tile_3_4_chanxy_out[56];
    assign wire_12144 = lut_tile_3_4_chanxy_out[57];
    assign wire_12146 = lut_tile_3_4_chanxy_out[58];
    assign wire_12148 = lut_tile_3_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_5_chanxy_in = {wire_12478, wire_7141, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7022, wire_3225, wire_12470, wire_7169, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7024, wire_3225, wire_12462, wire_7167, wire_7079, wire_7078, wire_7069, wire_7068, wire_7059, wire_7058, wire_7026, wire_3225, wire_12454, wire_7165, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7028, wire_2715, wire_12446, wire_7163, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7030, wire_2715, wire_12438, wire_7161, wire_7077, wire_7076, wire_7067, wire_7066, wire_7057, wire_7056, wire_7032, wire_2715, wire_12430, wire_7159, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7034, wire_3229, wire_2715, wire_12422, wire_7157, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7036, wire_3229, wire_2715, wire_12414, wire_7155, wire_7075, wire_7074, wire_7065, wire_7064, wire_7055, wire_7054, wire_7038, wire_3229, wire_2715, wire_12406, wire_7153, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7040, wire_3229, wire_2711, wire_12398, wire_7151, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7042, wire_3229, wire_2711, wire_12390, wire_7149, wire_7073, wire_7072, wire_7063, wire_7062, wire_7053, wire_7052, wire_7044, wire_3229, wire_2711, wire_12382, wire_7147, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7046, wire_3225, wire_2711, wire_12374, wire_7145, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7048, wire_3225, wire_2711, wire_12366, wire_7143, wire_7071, wire_7070, wire_7061, wire_7060, wire_7051, wire_7050, wire_7020, wire_3225, wire_2711, wire_12569, wire_7559, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7410, wire_3225, wire_12567, wire_7531, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7438, wire_3225, wire_12565, wire_7533, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7436, wire_3225, wire_12563, wire_7535, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7434, wire_2715, wire_12561, wire_7537, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7432, wire_2715, wire_12559, wire_7539, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7430, wire_2715, wire_12557, wire_7541, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7428, wire_3229, wire_2715, wire_12555, wire_7543, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7426, wire_3229, wire_2715, wire_12553, wire_7545, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7424, wire_3229, wire_2715, wire_12551, wire_7547, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7422, wire_3229, wire_2711, wire_12549, wire_7549, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7420, wire_3229, wire_2711, wire_12547, wire_7551, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7418, wire_3229, wire_2711, wire_12545, wire_7553, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7416, wire_3225, wire_2711, wire_12543, wire_7555, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7414, wire_3225, wire_2711, wire_12541, wire_7557, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7412, wire_3225, wire_2711, wire_12177, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12088, wire_7408, wire_2754, wire_12175, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_11976, wire_7400, wire_2754, wire_12173, wire_12083, wire_12082, wire_12043, wire_12042, wire_12003, wire_12002, wire_11984, wire_7392, wire_2754, wire_12171, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_11992, wire_7384, wire_2714, wire_12169, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12000, wire_7376, wire_2714, wire_12167, wire_12075, wire_12074, wire_12035, wire_12034, wire_12008, wire_11995, wire_11994, wire_7368, wire_2714, wire_12165, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12016, wire_7360, wire_2758, wire_2714, wire_12163, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12024, wire_7352, wire_2758, wire_2714, wire_12161, wire_12067, wire_12066, wire_12032, wire_12027, wire_12026, wire_11987, wire_11986, wire_7344, wire_2758, wire_2714, wire_12159, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12040, wire_7336, wire_2758, wire_2710, wire_12157, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12048, wire_7328, wire_2758, wire_2710, wire_12155, wire_12059, wire_12058, wire_12056, wire_12019, wire_12018, wire_11979, wire_11978, wire_7320, wire_2758, wire_2710, wire_12153, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12064, wire_7312, wire_2754, wire_2710, wire_12151, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12072, wire_7304, wire_2754, wire_2710, wire_12179, wire_12080, wire_12051, wire_12050, wire_12011, wire_12010, wire_11971, wire_11970, wire_7296, wire_2754, wire_2710, wire_12543, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12464, wire_7559, wire_2754, wire_12545, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12456, wire_7557, wire_2754, wire_12547, wire_12475, wire_12474, wire_12448, wire_12435, wire_12434, wire_12395, wire_12394, wire_7555, wire_2754, wire_12549, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12440, wire_7553, wire_2714, wire_12551, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12432, wire_7551, wire_2714, wire_12553, wire_12467, wire_12466, wire_12427, wire_12426, wire_12424, wire_12387, wire_12386, wire_7549, wire_2714, wire_12555, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12416, wire_7547, wire_2758, wire_2714, wire_12557, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12408, wire_7545, wire_2758, wire_2714, wire_12559, wire_12459, wire_12458, wire_12419, wire_12418, wire_12400, wire_12379, wire_12378, wire_7543, wire_2758, wire_2714, wire_12561, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12392, wire_7541, wire_2758, wire_2710, wire_12563, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12384, wire_7539, wire_2758, wire_2710, wire_12565, wire_12451, wire_12450, wire_12411, wire_12410, wire_12376, wire_12371, wire_12370, wire_7537, wire_2758, wire_2710, wire_12567, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12368, wire_7535, wire_2754, wire_2710, wire_12569, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12360, wire_7533, wire_2754, wire_2710, wire_12541, wire_12472, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_7531, wire_2754, wire_2710};
    // CHNAXY TOTAL: 636
    assign wire_7411 = lut_tile_3_5_chanxy_out[0];
    assign wire_7413 = lut_tile_3_5_chanxy_out[1];
    assign wire_7415 = lut_tile_3_5_chanxy_out[2];
    assign wire_7417 = lut_tile_3_5_chanxy_out[3];
    assign wire_7419 = lut_tile_3_5_chanxy_out[4];
    assign wire_7421 = lut_tile_3_5_chanxy_out[5];
    assign wire_7423 = lut_tile_3_5_chanxy_out[6];
    assign wire_7425 = lut_tile_3_5_chanxy_out[7];
    assign wire_7427 = lut_tile_3_5_chanxy_out[8];
    assign wire_7429 = lut_tile_3_5_chanxy_out[9];
    assign wire_7431 = lut_tile_3_5_chanxy_out[10];
    assign wire_7433 = lut_tile_3_5_chanxy_out[11];
    assign wire_7435 = lut_tile_3_5_chanxy_out[12];
    assign wire_7437 = lut_tile_3_5_chanxy_out[13];
    assign wire_7439 = lut_tile_3_5_chanxy_out[14];
    assign wire_7500 = lut_tile_3_5_chanxy_out[15];
    assign wire_7502 = lut_tile_3_5_chanxy_out[16];
    assign wire_7504 = lut_tile_3_5_chanxy_out[17];
    assign wire_7506 = lut_tile_3_5_chanxy_out[18];
    assign wire_7508 = lut_tile_3_5_chanxy_out[19];
    assign wire_7510 = lut_tile_3_5_chanxy_out[20];
    assign wire_7512 = lut_tile_3_5_chanxy_out[21];
    assign wire_7514 = lut_tile_3_5_chanxy_out[22];
    assign wire_7516 = lut_tile_3_5_chanxy_out[23];
    assign wire_7518 = lut_tile_3_5_chanxy_out[24];
    assign wire_7520 = lut_tile_3_5_chanxy_out[25];
    assign wire_7522 = lut_tile_3_5_chanxy_out[26];
    assign wire_7524 = lut_tile_3_5_chanxy_out[27];
    assign wire_7526 = lut_tile_3_5_chanxy_out[28];
    assign wire_7528 = lut_tile_3_5_chanxy_out[29];
    assign wire_12361 = lut_tile_3_5_chanxy_out[30];
    assign wire_12369 = lut_tile_3_5_chanxy_out[31];
    assign wire_12377 = lut_tile_3_5_chanxy_out[32];
    assign wire_12385 = lut_tile_3_5_chanxy_out[33];
    assign wire_12393 = lut_tile_3_5_chanxy_out[34];
    assign wire_12401 = lut_tile_3_5_chanxy_out[35];
    assign wire_12409 = lut_tile_3_5_chanxy_out[36];
    assign wire_12417 = lut_tile_3_5_chanxy_out[37];
    assign wire_12425 = lut_tile_3_5_chanxy_out[38];
    assign wire_12433 = lut_tile_3_5_chanxy_out[39];
    assign wire_12441 = lut_tile_3_5_chanxy_out[40];
    assign wire_12449 = lut_tile_3_5_chanxy_out[41];
    assign wire_12457 = lut_tile_3_5_chanxy_out[42];
    assign wire_12465 = lut_tile_3_5_chanxy_out[43];
    assign wire_12473 = lut_tile_3_5_chanxy_out[44];
    assign wire_12510 = lut_tile_3_5_chanxy_out[45];
    assign wire_12512 = lut_tile_3_5_chanxy_out[46];
    assign wire_12514 = lut_tile_3_5_chanxy_out[47];
    assign wire_12516 = lut_tile_3_5_chanxy_out[48];
    assign wire_12518 = lut_tile_3_5_chanxy_out[49];
    assign wire_12520 = lut_tile_3_5_chanxy_out[50];
    assign wire_12522 = lut_tile_3_5_chanxy_out[51];
    assign wire_12524 = lut_tile_3_5_chanxy_out[52];
    assign wire_12526 = lut_tile_3_5_chanxy_out[53];
    assign wire_12528 = lut_tile_3_5_chanxy_out[54];
    assign wire_12530 = lut_tile_3_5_chanxy_out[55];
    assign wire_12532 = lut_tile_3_5_chanxy_out[56];
    assign wire_12534 = lut_tile_3_5_chanxy_out[57];
    assign wire_12536 = lut_tile_3_5_chanxy_out[58];
    assign wire_12538 = lut_tile_3_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_6_chanxy_in = {wire_12862, wire_7171, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7052, wire_3741, wire_12854, wire_7199, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7054, wire_3741, wire_12846, wire_7197, wire_7109, wire_7108, wire_7099, wire_7098, wire_7089, wire_7088, wire_7056, wire_3741, wire_12838, wire_7195, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7058, wire_3231, wire_12830, wire_7193, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7060, wire_3231, wire_12822, wire_7191, wire_7107, wire_7106, wire_7097, wire_7096, wire_7087, wire_7086, wire_7062, wire_3231, wire_12814, wire_7189, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7064, wire_3745, wire_3231, wire_12806, wire_7187, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7066, wire_3745, wire_3231, wire_12798, wire_7185, wire_7105, wire_7104, wire_7095, wire_7094, wire_7085, wire_7084, wire_7068, wire_3745, wire_3231, wire_12790, wire_7183, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7070, wire_3745, wire_3227, wire_12782, wire_7181, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7072, wire_3745, wire_3227, wire_12774, wire_7179, wire_7103, wire_7102, wire_7093, wire_7092, wire_7083, wire_7082, wire_7074, wire_3745, wire_3227, wire_12766, wire_7177, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7076, wire_3741, wire_3227, wire_12758, wire_7175, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7078, wire_3741, wire_3227, wire_12750, wire_7173, wire_7101, wire_7100, wire_7091, wire_7090, wire_7081, wire_7080, wire_7050, wire_3741, wire_3227, wire_12959, wire_7589, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7440, wire_3741, wire_12957, wire_7561, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7468, wire_3741, wire_12955, wire_7563, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7466, wire_3741, wire_12953, wire_7565, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7464, wire_3231, wire_12951, wire_7567, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7462, wire_3231, wire_12949, wire_7569, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7460, wire_3231, wire_12947, wire_7571, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7458, wire_3745, wire_3231, wire_12945, wire_7573, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7456, wire_3745, wire_3231, wire_12943, wire_7575, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7454, wire_3745, wire_3231, wire_12941, wire_7577, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7452, wire_3745, wire_3227, wire_12939, wire_7579, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7450, wire_3745, wire_3227, wire_12937, wire_7581, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7448, wire_3745, wire_3227, wire_12935, wire_7583, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7446, wire_3741, wire_3227, wire_12933, wire_7585, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7444, wire_3741, wire_3227, wire_12931, wire_7587, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7442, wire_3741, wire_3227, wire_12567, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12472, wire_7438, wire_3270, wire_12565, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12360, wire_7436, wire_3270, wire_12563, wire_12475, wire_12474, wire_12435, wire_12434, wire_12395, wire_12394, wire_12368, wire_7434, wire_3270, wire_12561, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12376, wire_7432, wire_3230, wire_12559, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12384, wire_7430, wire_3230, wire_12557, wire_12467, wire_12466, wire_12427, wire_12426, wire_12392, wire_12387, wire_12386, wire_7428, wire_3230, wire_12555, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12400, wire_7426, wire_3274, wire_3230, wire_12553, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12408, wire_7424, wire_3274, wire_3230, wire_12551, wire_12459, wire_12458, wire_12419, wire_12418, wire_12416, wire_12379, wire_12378, wire_7422, wire_3274, wire_3230, wire_12549, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12424, wire_7420, wire_3274, wire_3226, wire_12547, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12432, wire_7418, wire_3274, wire_3226, wire_12545, wire_12451, wire_12450, wire_12440, wire_12411, wire_12410, wire_12371, wire_12370, wire_7416, wire_3274, wire_3226, wire_12543, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12448, wire_7414, wire_3270, wire_3226, wire_12541, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12456, wire_7412, wire_3270, wire_3226, wire_12569, wire_12464, wire_12443, wire_12442, wire_12403, wire_12402, wire_12363, wire_12362, wire_7410, wire_3270, wire_3226, wire_12933, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12856, wire_7589, wire_3270, wire_12935, wire_12867, wire_12866, wire_12848, wire_12827, wire_12826, wire_12787, wire_12786, wire_7587, wire_3270, wire_12937, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12840, wire_7585, wire_3270, wire_12939, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12832, wire_7583, wire_3230, wire_12941, wire_12859, wire_12858, wire_12824, wire_12819, wire_12818, wire_12779, wire_12778, wire_7581, wire_3230, wire_12943, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12816, wire_7579, wire_3230, wire_12945, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12808, wire_7577, wire_3274, wire_3230, wire_12947, wire_12851, wire_12850, wire_12811, wire_12810, wire_12800, wire_12771, wire_12770, wire_7575, wire_3274, wire_3230, wire_12949, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12792, wire_7573, wire_3274, wire_3230, wire_12951, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12784, wire_7571, wire_3274, wire_3226, wire_12953, wire_12843, wire_12842, wire_12803, wire_12802, wire_12776, wire_12763, wire_12762, wire_7569, wire_3274, wire_3226, wire_12955, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12768, wire_7567, wire_3274, wire_3226, wire_12957, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12760, wire_7565, wire_3270, wire_3226, wire_12959, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_12752, wire_7563, wire_3270, wire_3226, wire_12931, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12864, wire_7561, wire_3270, wire_3226};
    // CHNAXY TOTAL: 636
    assign wire_7441 = lut_tile_3_6_chanxy_out[0];
    assign wire_7443 = lut_tile_3_6_chanxy_out[1];
    assign wire_7445 = lut_tile_3_6_chanxy_out[2];
    assign wire_7447 = lut_tile_3_6_chanxy_out[3];
    assign wire_7449 = lut_tile_3_6_chanxy_out[4];
    assign wire_7451 = lut_tile_3_6_chanxy_out[5];
    assign wire_7453 = lut_tile_3_6_chanxy_out[6];
    assign wire_7455 = lut_tile_3_6_chanxy_out[7];
    assign wire_7457 = lut_tile_3_6_chanxy_out[8];
    assign wire_7459 = lut_tile_3_6_chanxy_out[9];
    assign wire_7461 = lut_tile_3_6_chanxy_out[10];
    assign wire_7463 = lut_tile_3_6_chanxy_out[11];
    assign wire_7465 = lut_tile_3_6_chanxy_out[12];
    assign wire_7467 = lut_tile_3_6_chanxy_out[13];
    assign wire_7469 = lut_tile_3_6_chanxy_out[14];
    assign wire_7530 = lut_tile_3_6_chanxy_out[15];
    assign wire_7532 = lut_tile_3_6_chanxy_out[16];
    assign wire_7534 = lut_tile_3_6_chanxy_out[17];
    assign wire_7536 = lut_tile_3_6_chanxy_out[18];
    assign wire_7538 = lut_tile_3_6_chanxy_out[19];
    assign wire_7540 = lut_tile_3_6_chanxy_out[20];
    assign wire_7542 = lut_tile_3_6_chanxy_out[21];
    assign wire_7544 = lut_tile_3_6_chanxy_out[22];
    assign wire_7546 = lut_tile_3_6_chanxy_out[23];
    assign wire_7548 = lut_tile_3_6_chanxy_out[24];
    assign wire_7550 = lut_tile_3_6_chanxy_out[25];
    assign wire_7552 = lut_tile_3_6_chanxy_out[26];
    assign wire_7554 = lut_tile_3_6_chanxy_out[27];
    assign wire_7556 = lut_tile_3_6_chanxy_out[28];
    assign wire_7558 = lut_tile_3_6_chanxy_out[29];
    assign wire_12753 = lut_tile_3_6_chanxy_out[30];
    assign wire_12761 = lut_tile_3_6_chanxy_out[31];
    assign wire_12769 = lut_tile_3_6_chanxy_out[32];
    assign wire_12777 = lut_tile_3_6_chanxy_out[33];
    assign wire_12785 = lut_tile_3_6_chanxy_out[34];
    assign wire_12793 = lut_tile_3_6_chanxy_out[35];
    assign wire_12801 = lut_tile_3_6_chanxy_out[36];
    assign wire_12809 = lut_tile_3_6_chanxy_out[37];
    assign wire_12817 = lut_tile_3_6_chanxy_out[38];
    assign wire_12825 = lut_tile_3_6_chanxy_out[39];
    assign wire_12833 = lut_tile_3_6_chanxy_out[40];
    assign wire_12841 = lut_tile_3_6_chanxy_out[41];
    assign wire_12849 = lut_tile_3_6_chanxy_out[42];
    assign wire_12857 = lut_tile_3_6_chanxy_out[43];
    assign wire_12865 = lut_tile_3_6_chanxy_out[44];
    assign wire_12900 = lut_tile_3_6_chanxy_out[45];
    assign wire_12902 = lut_tile_3_6_chanxy_out[46];
    assign wire_12904 = lut_tile_3_6_chanxy_out[47];
    assign wire_12906 = lut_tile_3_6_chanxy_out[48];
    assign wire_12908 = lut_tile_3_6_chanxy_out[49];
    assign wire_12910 = lut_tile_3_6_chanxy_out[50];
    assign wire_12912 = lut_tile_3_6_chanxy_out[51];
    assign wire_12914 = lut_tile_3_6_chanxy_out[52];
    assign wire_12916 = lut_tile_3_6_chanxy_out[53];
    assign wire_12918 = lut_tile_3_6_chanxy_out[54];
    assign wire_12920 = lut_tile_3_6_chanxy_out[55];
    assign wire_12922 = lut_tile_3_6_chanxy_out[56];
    assign wire_12924 = lut_tile_3_6_chanxy_out[57];
    assign wire_12926 = lut_tile_3_6_chanxy_out[58];
    assign wire_12928 = lut_tile_3_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_7_chanxy_in = {wire_13254, wire_7201, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7082, wire_4257, wire_13246, wire_7229, wire_7139, wire_7138, wire_7129, wire_7128, wire_7119, wire_7118, wire_7084, wire_4257, wire_13238, wire_7227, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7086, wire_4257, wire_13230, wire_7225, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7088, wire_3747, wire_13222, wire_7223, wire_7137, wire_7136, wire_7127, wire_7126, wire_7117, wire_7116, wire_7090, wire_3747, wire_13214, wire_7221, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7092, wire_3747, wire_13206, wire_7219, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7094, wire_4261, wire_3747, wire_13198, wire_7217, wire_7135, wire_7134, wire_7125, wire_7124, wire_7115, wire_7114, wire_7096, wire_4261, wire_3747, wire_13190, wire_7215, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7098, wire_4261, wire_3747, wire_13182, wire_7213, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7100, wire_4261, wire_3743, wire_13174, wire_7211, wire_7133, wire_7132, wire_7123, wire_7122, wire_7113, wire_7112, wire_7102, wire_4261, wire_3743, wire_13166, wire_7209, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7104, wire_4261, wire_3743, wire_13158, wire_7207, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7106, wire_4257, wire_3743, wire_13150, wire_7205, wire_7131, wire_7130, wire_7121, wire_7120, wire_7111, wire_7110, wire_7108, wire_4257, wire_3743, wire_13142, wire_7203, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7080, wire_4257, wire_3743, wire_13349, wire_7619, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7470, wire_4257, wire_13347, wire_7591, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7498, wire_4257, wire_13345, wire_7593, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7496, wire_4257, wire_13343, wire_7595, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7494, wire_3747, wire_13341, wire_7597, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7492, wire_3747, wire_13339, wire_7599, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7490, wire_3747, wire_13337, wire_7601, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7488, wire_4261, wire_3747, wire_13335, wire_7603, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7486, wire_4261, wire_3747, wire_13333, wire_7605, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7484, wire_4261, wire_3747, wire_13331, wire_7607, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7482, wire_4261, wire_3743, wire_13329, wire_7609, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7480, wire_4261, wire_3743, wire_13327, wire_7611, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7478, wire_4261, wire_3743, wire_13325, wire_7613, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7476, wire_4257, wire_3743, wire_13323, wire_7615, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7474, wire_4257, wire_3743, wire_13321, wire_7617, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7472, wire_4257, wire_3743, wire_12957, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12864, wire_7468, wire_3786, wire_12955, wire_12867, wire_12866, wire_12827, wire_12826, wire_12787, wire_12786, wire_12752, wire_7466, wire_3786, wire_12953, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12760, wire_7464, wire_3786, wire_12951, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12768, wire_7462, wire_3746, wire_12949, wire_12859, wire_12858, wire_12819, wire_12818, wire_12779, wire_12778, wire_12776, wire_7460, wire_3746, wire_12947, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12784, wire_7458, wire_3746, wire_12945, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12792, wire_7456, wire_3790, wire_3746, wire_12943, wire_12851, wire_12850, wire_12811, wire_12810, wire_12800, wire_12771, wire_12770, wire_7454, wire_3790, wire_3746, wire_12941, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12808, wire_7452, wire_3790, wire_3746, wire_12939, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12816, wire_7450, wire_3790, wire_3742, wire_12937, wire_12843, wire_12842, wire_12824, wire_12803, wire_12802, wire_12763, wire_12762, wire_7448, wire_3790, wire_3742, wire_12935, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12832, wire_7446, wire_3790, wire_3742, wire_12933, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12840, wire_7444, wire_3786, wire_3742, wire_12931, wire_12848, wire_12835, wire_12834, wire_12795, wire_12794, wire_12755, wire_12754, wire_7442, wire_3786, wire_3742, wire_12959, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12856, wire_7440, wire_3786, wire_3742, wire_13323, wire_13259, wire_13258, wire_13248, wire_13219, wire_13218, wire_13179, wire_13178, wire_7619, wire_3786, wire_13325, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13240, wire_7617, wire_3786, wire_13327, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13232, wire_7615, wire_3786, wire_13329, wire_13251, wire_13250, wire_13224, wire_13211, wire_13210, wire_13171, wire_13170, wire_7613, wire_3746, wire_13331, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13216, wire_7611, wire_3746, wire_13333, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13208, wire_7609, wire_3746, wire_13335, wire_13243, wire_13242, wire_13203, wire_13202, wire_13200, wire_13163, wire_13162, wire_7607, wire_3790, wire_3746, wire_13337, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13192, wire_7605, wire_3790, wire_3746, wire_13339, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13184, wire_7603, wire_3790, wire_3746, wire_13341, wire_13235, wire_13234, wire_13195, wire_13194, wire_13176, wire_13155, wire_13154, wire_7601, wire_3790, wire_3742, wire_13343, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13168, wire_7599, wire_3790, wire_3742, wire_13345, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13160, wire_7597, wire_3790, wire_3742, wire_13347, wire_13227, wire_13226, wire_13187, wire_13186, wire_13152, wire_13147, wire_13146, wire_7595, wire_3786, wire_3742, wire_13349, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13144, wire_7593, wire_3786, wire_3742, wire_13321, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13256, wire_7591, wire_3786, wire_3742};
    // CHNAXY TOTAL: 636
    assign wire_7471 = lut_tile_3_7_chanxy_out[0];
    assign wire_7473 = lut_tile_3_7_chanxy_out[1];
    assign wire_7475 = lut_tile_3_7_chanxy_out[2];
    assign wire_7477 = lut_tile_3_7_chanxy_out[3];
    assign wire_7479 = lut_tile_3_7_chanxy_out[4];
    assign wire_7481 = lut_tile_3_7_chanxy_out[5];
    assign wire_7483 = lut_tile_3_7_chanxy_out[6];
    assign wire_7485 = lut_tile_3_7_chanxy_out[7];
    assign wire_7487 = lut_tile_3_7_chanxy_out[8];
    assign wire_7489 = lut_tile_3_7_chanxy_out[9];
    assign wire_7491 = lut_tile_3_7_chanxy_out[10];
    assign wire_7493 = lut_tile_3_7_chanxy_out[11];
    assign wire_7495 = lut_tile_3_7_chanxy_out[12];
    assign wire_7497 = lut_tile_3_7_chanxy_out[13];
    assign wire_7499 = lut_tile_3_7_chanxy_out[14];
    assign wire_7560 = lut_tile_3_7_chanxy_out[15];
    assign wire_7562 = lut_tile_3_7_chanxy_out[16];
    assign wire_7564 = lut_tile_3_7_chanxy_out[17];
    assign wire_7566 = lut_tile_3_7_chanxy_out[18];
    assign wire_7568 = lut_tile_3_7_chanxy_out[19];
    assign wire_7570 = lut_tile_3_7_chanxy_out[20];
    assign wire_7572 = lut_tile_3_7_chanxy_out[21];
    assign wire_7574 = lut_tile_3_7_chanxy_out[22];
    assign wire_7576 = lut_tile_3_7_chanxy_out[23];
    assign wire_7578 = lut_tile_3_7_chanxy_out[24];
    assign wire_7580 = lut_tile_3_7_chanxy_out[25];
    assign wire_7582 = lut_tile_3_7_chanxy_out[26];
    assign wire_7584 = lut_tile_3_7_chanxy_out[27];
    assign wire_7586 = lut_tile_3_7_chanxy_out[28];
    assign wire_7588 = lut_tile_3_7_chanxy_out[29];
    assign wire_13145 = lut_tile_3_7_chanxy_out[30];
    assign wire_13153 = lut_tile_3_7_chanxy_out[31];
    assign wire_13161 = lut_tile_3_7_chanxy_out[32];
    assign wire_13169 = lut_tile_3_7_chanxy_out[33];
    assign wire_13177 = lut_tile_3_7_chanxy_out[34];
    assign wire_13185 = lut_tile_3_7_chanxy_out[35];
    assign wire_13193 = lut_tile_3_7_chanxy_out[36];
    assign wire_13201 = lut_tile_3_7_chanxy_out[37];
    assign wire_13209 = lut_tile_3_7_chanxy_out[38];
    assign wire_13217 = lut_tile_3_7_chanxy_out[39];
    assign wire_13225 = lut_tile_3_7_chanxy_out[40];
    assign wire_13233 = lut_tile_3_7_chanxy_out[41];
    assign wire_13241 = lut_tile_3_7_chanxy_out[42];
    assign wire_13249 = lut_tile_3_7_chanxy_out[43];
    assign wire_13257 = lut_tile_3_7_chanxy_out[44];
    assign wire_13290 = lut_tile_3_7_chanxy_out[45];
    assign wire_13292 = lut_tile_3_7_chanxy_out[46];
    assign wire_13294 = lut_tile_3_7_chanxy_out[47];
    assign wire_13296 = lut_tile_3_7_chanxy_out[48];
    assign wire_13298 = lut_tile_3_7_chanxy_out[49];
    assign wire_13300 = lut_tile_3_7_chanxy_out[50];
    assign wire_13302 = lut_tile_3_7_chanxy_out[51];
    assign wire_13304 = lut_tile_3_7_chanxy_out[52];
    assign wire_13306 = lut_tile_3_7_chanxy_out[53];
    assign wire_13308 = lut_tile_3_7_chanxy_out[54];
    assign wire_13310 = lut_tile_3_7_chanxy_out[55];
    assign wire_13312 = lut_tile_3_7_chanxy_out[56];
    assign wire_13314 = lut_tile_3_7_chanxy_out[57];
    assign wire_13316 = lut_tile_3_7_chanxy_out[58];
    assign wire_13318 = lut_tile_3_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_8_chanxy_in = {wire_13646, wire_7231, wire_7169, wire_7168, wire_7159, wire_7158, wire_7149, wire_7148, wire_7112, wire_4773, wire_13638, wire_7259, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7114, wire_4773, wire_13630, wire_7257, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7116, wire_4773, wire_13622, wire_7255, wire_7167, wire_7166, wire_7157, wire_7156, wire_7147, wire_7146, wire_7118, wire_4263, wire_13614, wire_7253, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7120, wire_4263, wire_13606, wire_7251, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7122, wire_4263, wire_13598, wire_7249, wire_7165, wire_7164, wire_7155, wire_7154, wire_7145, wire_7144, wire_7124, wire_4777, wire_4263, wire_13590, wire_7247, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7126, wire_4777, wire_4263, wire_13582, wire_7245, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7128, wire_4777, wire_4263, wire_13574, wire_7243, wire_7163, wire_7162, wire_7153, wire_7152, wire_7143, wire_7142, wire_7130, wire_4777, wire_4259, wire_13566, wire_7241, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7132, wire_4777, wire_4259, wire_13558, wire_7239, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7134, wire_4777, wire_4259, wire_13550, wire_7237, wire_7161, wire_7160, wire_7151, wire_7150, wire_7141, wire_7140, wire_7136, wire_4773, wire_4259, wire_13542, wire_7235, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7138, wire_4773, wire_4259, wire_13534, wire_7233, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7110, wire_4773, wire_4259, wire_13739, wire_7649, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7500, wire_4773, wire_13737, wire_7621, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7528, wire_4773, wire_13735, wire_7623, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7526, wire_4773, wire_13733, wire_7625, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7524, wire_4263, wire_13731, wire_7627, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7522, wire_4263, wire_13729, wire_7629, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7520, wire_4263, wire_13727, wire_7631, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7518, wire_4777, wire_4263, wire_13725, wire_7633, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7516, wire_4777, wire_4263, wire_13723, wire_7635, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7514, wire_4777, wire_4263, wire_13721, wire_7637, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7512, wire_4777, wire_4259, wire_13719, wire_7639, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7510, wire_4777, wire_4259, wire_13717, wire_7641, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7508, wire_4777, wire_4259, wire_13715, wire_7643, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7506, wire_4773, wire_4259, wire_13713, wire_7645, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7504, wire_4773, wire_4259, wire_13711, wire_7647, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7502, wire_4773, wire_4259, wire_13347, wire_13259, wire_13258, wire_13256, wire_13219, wire_13218, wire_13179, wire_13178, wire_7498, wire_4302, wire_13345, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13144, wire_7496, wire_4302, wire_13343, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13152, wire_7494, wire_4302, wire_13341, wire_13251, wire_13250, wire_13211, wire_13210, wire_13171, wire_13170, wire_13160, wire_7492, wire_4262, wire_13339, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13168, wire_7490, wire_4262, wire_13337, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13176, wire_7488, wire_4262, wire_13335, wire_13243, wire_13242, wire_13203, wire_13202, wire_13184, wire_13163, wire_13162, wire_7486, wire_4306, wire_4262, wire_13333, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13192, wire_7484, wire_4306, wire_4262, wire_13331, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13200, wire_7482, wire_4306, wire_4262, wire_13329, wire_13235, wire_13234, wire_13208, wire_13195, wire_13194, wire_13155, wire_13154, wire_7480, wire_4306, wire_4258, wire_13327, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13216, wire_7478, wire_4306, wire_4258, wire_13325, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13224, wire_7476, wire_4306, wire_4258, wire_13323, wire_13232, wire_13227, wire_13226, wire_13187, wire_13186, wire_13147, wire_13146, wire_7474, wire_4302, wire_4258, wire_13321, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13240, wire_7472, wire_4302, wire_4258, wire_13349, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13248, wire_7470, wire_4302, wire_4258, wire_13713, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13640, wire_7649, wire_4302, wire_13715, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13632, wire_7647, wire_4302, wire_13717, wire_13643, wire_13642, wire_13624, wire_13603, wire_13602, wire_13563, wire_13562, wire_7645, wire_4302, wire_13719, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13616, wire_7643, wire_4262, wire_13721, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13608, wire_7641, wire_4262, wire_13723, wire_13635, wire_13634, wire_13600, wire_13595, wire_13594, wire_13555, wire_13554, wire_7639, wire_4262, wire_13725, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13592, wire_7637, wire_4306, wire_4262, wire_13727, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13584, wire_7635, wire_4306, wire_4262, wire_13729, wire_13627, wire_13626, wire_13587, wire_13586, wire_13576, wire_13547, wire_13546, wire_7633, wire_4306, wire_4262, wire_13731, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13568, wire_7631, wire_4306, wire_4258, wire_13733, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13560, wire_7629, wire_4306, wire_4258, wire_13735, wire_13619, wire_13618, wire_13579, wire_13578, wire_13552, wire_13539, wire_13538, wire_7627, wire_4306, wire_4258, wire_13737, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13544, wire_7625, wire_4302, wire_4258, wire_13739, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13536, wire_7623, wire_4302, wire_4258, wire_13711, wire_13648, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7621, wire_4302, wire_4258};
    // CHNAXY TOTAL: 636
    assign wire_7501 = lut_tile_3_8_chanxy_out[0];
    assign wire_7503 = lut_tile_3_8_chanxy_out[1];
    assign wire_7505 = lut_tile_3_8_chanxy_out[2];
    assign wire_7507 = lut_tile_3_8_chanxy_out[3];
    assign wire_7509 = lut_tile_3_8_chanxy_out[4];
    assign wire_7511 = lut_tile_3_8_chanxy_out[5];
    assign wire_7513 = lut_tile_3_8_chanxy_out[6];
    assign wire_7515 = lut_tile_3_8_chanxy_out[7];
    assign wire_7517 = lut_tile_3_8_chanxy_out[8];
    assign wire_7519 = lut_tile_3_8_chanxy_out[9];
    assign wire_7521 = lut_tile_3_8_chanxy_out[10];
    assign wire_7523 = lut_tile_3_8_chanxy_out[11];
    assign wire_7525 = lut_tile_3_8_chanxy_out[12];
    assign wire_7527 = lut_tile_3_8_chanxy_out[13];
    assign wire_7529 = lut_tile_3_8_chanxy_out[14];
    assign wire_7590 = lut_tile_3_8_chanxy_out[15];
    assign wire_7592 = lut_tile_3_8_chanxy_out[16];
    assign wire_7594 = lut_tile_3_8_chanxy_out[17];
    assign wire_7596 = lut_tile_3_8_chanxy_out[18];
    assign wire_7598 = lut_tile_3_8_chanxy_out[19];
    assign wire_7600 = lut_tile_3_8_chanxy_out[20];
    assign wire_7602 = lut_tile_3_8_chanxy_out[21];
    assign wire_7604 = lut_tile_3_8_chanxy_out[22];
    assign wire_7606 = lut_tile_3_8_chanxy_out[23];
    assign wire_7608 = lut_tile_3_8_chanxy_out[24];
    assign wire_7610 = lut_tile_3_8_chanxy_out[25];
    assign wire_7612 = lut_tile_3_8_chanxy_out[26];
    assign wire_7614 = lut_tile_3_8_chanxy_out[27];
    assign wire_7616 = lut_tile_3_8_chanxy_out[28];
    assign wire_7618 = lut_tile_3_8_chanxy_out[29];
    assign wire_13537 = lut_tile_3_8_chanxy_out[30];
    assign wire_13545 = lut_tile_3_8_chanxy_out[31];
    assign wire_13553 = lut_tile_3_8_chanxy_out[32];
    assign wire_13561 = lut_tile_3_8_chanxy_out[33];
    assign wire_13569 = lut_tile_3_8_chanxy_out[34];
    assign wire_13577 = lut_tile_3_8_chanxy_out[35];
    assign wire_13585 = lut_tile_3_8_chanxy_out[36];
    assign wire_13593 = lut_tile_3_8_chanxy_out[37];
    assign wire_13601 = lut_tile_3_8_chanxy_out[38];
    assign wire_13609 = lut_tile_3_8_chanxy_out[39];
    assign wire_13617 = lut_tile_3_8_chanxy_out[40];
    assign wire_13625 = lut_tile_3_8_chanxy_out[41];
    assign wire_13633 = lut_tile_3_8_chanxy_out[42];
    assign wire_13641 = lut_tile_3_8_chanxy_out[43];
    assign wire_13649 = lut_tile_3_8_chanxy_out[44];
    assign wire_13680 = lut_tile_3_8_chanxy_out[45];
    assign wire_13682 = lut_tile_3_8_chanxy_out[46];
    assign wire_13684 = lut_tile_3_8_chanxy_out[47];
    assign wire_13686 = lut_tile_3_8_chanxy_out[48];
    assign wire_13688 = lut_tile_3_8_chanxy_out[49];
    assign wire_13690 = lut_tile_3_8_chanxy_out[50];
    assign wire_13692 = lut_tile_3_8_chanxy_out[51];
    assign wire_13694 = lut_tile_3_8_chanxy_out[52];
    assign wire_13696 = lut_tile_3_8_chanxy_out[53];
    assign wire_13698 = lut_tile_3_8_chanxy_out[54];
    assign wire_13700 = lut_tile_3_8_chanxy_out[55];
    assign wire_13702 = lut_tile_3_8_chanxy_out[56];
    assign wire_13704 = lut_tile_3_8_chanxy_out[57];
    assign wire_13706 = lut_tile_3_8_chanxy_out[58];
    assign wire_13708 = lut_tile_3_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_9_chanxy_in = {wire_14038, wire_7261, wire_7259, wire_7258, wire_7249, wire_7248, wire_7239, wire_7238, wire_7142, wire_5289, wire_14030, wire_7289, wire_7229, wire_7228, wire_7219, wire_7218, wire_7209, wire_7208, wire_7144, wire_5289, wire_14022, wire_7287, wire_7199, wire_7198, wire_7189, wire_7188, wire_7179, wire_7178, wire_7146, wire_5289, wire_14014, wire_7285, wire_7257, wire_7256, wire_7247, wire_7246, wire_7237, wire_7236, wire_7148, wire_4779, wire_14006, wire_7283, wire_7227, wire_7226, wire_7217, wire_7216, wire_7207, wire_7206, wire_7150, wire_4779, wire_13998, wire_7281, wire_7197, wire_7196, wire_7187, wire_7186, wire_7177, wire_7176, wire_7152, wire_4779, wire_13990, wire_7279, wire_7255, wire_7254, wire_7245, wire_7244, wire_7235, wire_7234, wire_7154, wire_5293, wire_4779, wire_13982, wire_7277, wire_7225, wire_7224, wire_7215, wire_7214, wire_7205, wire_7204, wire_7156, wire_5293, wire_4779, wire_13974, wire_7275, wire_7195, wire_7194, wire_7185, wire_7184, wire_7175, wire_7174, wire_7158, wire_5293, wire_4779, wire_13966, wire_7273, wire_7253, wire_7252, wire_7243, wire_7242, wire_7233, wire_7232, wire_7160, wire_5293, wire_4775, wire_13958, wire_7271, wire_7223, wire_7222, wire_7213, wire_7212, wire_7203, wire_7202, wire_7162, wire_5293, wire_4775, wire_13950, wire_7269, wire_7193, wire_7192, wire_7183, wire_7182, wire_7173, wire_7172, wire_7164, wire_5293, wire_4775, wire_13942, wire_7267, wire_7251, wire_7250, wire_7241, wire_7240, wire_7231, wire_7230, wire_7166, wire_5289, wire_4775, wire_13934, wire_7265, wire_7221, wire_7220, wire_7211, wire_7210, wire_7201, wire_7200, wire_7168, wire_5289, wire_4775, wire_13926, wire_7263, wire_7191, wire_7190, wire_7181, wire_7180, wire_7171, wire_7170, wire_7140, wire_5289, wire_4775, wire_14129, wire_7679, wire_7649, wire_7648, wire_7639, wire_7638, wire_7629, wire_7628, wire_7530, wire_5289, wire_14127, wire_7651, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7558, wire_5289, wire_14125, wire_7653, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7556, wire_5289, wire_14123, wire_7655, wire_7647, wire_7646, wire_7637, wire_7636, wire_7627, wire_7626, wire_7554, wire_4779, wire_14121, wire_7657, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7552, wire_4779, wire_14119, wire_7659, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7550, wire_4779, wire_14117, wire_7661, wire_7645, wire_7644, wire_7635, wire_7634, wire_7625, wire_7624, wire_7548, wire_5293, wire_4779, wire_14115, wire_7663, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7546, wire_5293, wire_4779, wire_14113, wire_7665, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7544, wire_5293, wire_4779, wire_14111, wire_7667, wire_7643, wire_7642, wire_7633, wire_7632, wire_7623, wire_7622, wire_7542, wire_5293, wire_4775, wire_14109, wire_7669, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7540, wire_5293, wire_4775, wire_14107, wire_7671, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7538, wire_5293, wire_4775, wire_14105, wire_7673, wire_7641, wire_7640, wire_7631, wire_7630, wire_7621, wire_7620, wire_7536, wire_5289, wire_4775, wire_14103, wire_7675, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7534, wire_5289, wire_4775, wire_14101, wire_7677, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7532, wire_5289, wire_4775, wire_13737, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13648, wire_7528, wire_4818, wire_13735, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13536, wire_7526, wire_4818, wire_13733, wire_13643, wire_13642, wire_13603, wire_13602, wire_13563, wire_13562, wire_13544, wire_7524, wire_4818, wire_13731, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13552, wire_7522, wire_4778, wire_13729, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13560, wire_7520, wire_4778, wire_13727, wire_13635, wire_13634, wire_13595, wire_13594, wire_13568, wire_13555, wire_13554, wire_7518, wire_4778, wire_13725, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13576, wire_7516, wire_4822, wire_4778, wire_13723, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13584, wire_7514, wire_4822, wire_4778, wire_13721, wire_13627, wire_13626, wire_13592, wire_13587, wire_13586, wire_13547, wire_13546, wire_7512, wire_4822, wire_4778, wire_13719, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13600, wire_7510, wire_4822, wire_4774, wire_13717, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13608, wire_7508, wire_4822, wire_4774, wire_13715, wire_13619, wire_13618, wire_13616, wire_13579, wire_13578, wire_13539, wire_13538, wire_7506, wire_4822, wire_4774, wire_13713, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13624, wire_7504, wire_4818, wire_4774, wire_13711, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13632, wire_7502, wire_4818, wire_4774, wire_13739, wire_13640, wire_13611, wire_13610, wire_13571, wire_13570, wire_13531, wire_13530, wire_7500, wire_4818, wire_4774, wire_14103, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14024, wire_7679, wire_4818, wire_14105, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14016, wire_7677, wire_4818, wire_14107, wire_14035, wire_14034, wire_14008, wire_13995, wire_13994, wire_13955, wire_13954, wire_7675, wire_4818, wire_14109, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14000, wire_7673, wire_4778, wire_14111, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_13992, wire_7671, wire_4778, wire_14113, wire_14027, wire_14026, wire_13987, wire_13986, wire_13984, wire_13947, wire_13946, wire_7669, wire_4778, wire_14115, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_13976, wire_7667, wire_4822, wire_4778, wire_14117, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13968, wire_7665, wire_4822, wire_4778, wire_14119, wire_14019, wire_14018, wire_13979, wire_13978, wire_13960, wire_13939, wire_13938, wire_7663, wire_4822, wire_4778, wire_14121, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_13952, wire_7661, wire_4822, wire_4774, wire_14123, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13944, wire_7659, wire_4822, wire_4774, wire_14125, wire_14011, wire_14010, wire_13971, wire_13970, wire_13936, wire_13931, wire_13930, wire_7657, wire_4822, wire_4774, wire_14127, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_13928, wire_7655, wire_4818, wire_4774, wire_14129, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_13920, wire_7653, wire_4818, wire_4774, wire_14101, wire_14032, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_7651, wire_4818, wire_4774};
    // CHNAXY TOTAL: 636
    assign wire_7531 = lut_tile_3_9_chanxy_out[0];
    assign wire_7533 = lut_tile_3_9_chanxy_out[1];
    assign wire_7535 = lut_tile_3_9_chanxy_out[2];
    assign wire_7537 = lut_tile_3_9_chanxy_out[3];
    assign wire_7539 = lut_tile_3_9_chanxy_out[4];
    assign wire_7541 = lut_tile_3_9_chanxy_out[5];
    assign wire_7543 = lut_tile_3_9_chanxy_out[6];
    assign wire_7545 = lut_tile_3_9_chanxy_out[7];
    assign wire_7547 = lut_tile_3_9_chanxy_out[8];
    assign wire_7549 = lut_tile_3_9_chanxy_out[9];
    assign wire_7551 = lut_tile_3_9_chanxy_out[10];
    assign wire_7553 = lut_tile_3_9_chanxy_out[11];
    assign wire_7555 = lut_tile_3_9_chanxy_out[12];
    assign wire_7557 = lut_tile_3_9_chanxy_out[13];
    assign wire_7559 = lut_tile_3_9_chanxy_out[14];
    assign wire_7620 = lut_tile_3_9_chanxy_out[15];
    assign wire_7622 = lut_tile_3_9_chanxy_out[16];
    assign wire_7624 = lut_tile_3_9_chanxy_out[17];
    assign wire_7626 = lut_tile_3_9_chanxy_out[18];
    assign wire_7628 = lut_tile_3_9_chanxy_out[19];
    assign wire_7630 = lut_tile_3_9_chanxy_out[20];
    assign wire_7632 = lut_tile_3_9_chanxy_out[21];
    assign wire_7634 = lut_tile_3_9_chanxy_out[22];
    assign wire_7636 = lut_tile_3_9_chanxy_out[23];
    assign wire_7638 = lut_tile_3_9_chanxy_out[24];
    assign wire_7640 = lut_tile_3_9_chanxy_out[25];
    assign wire_7642 = lut_tile_3_9_chanxy_out[26];
    assign wire_7644 = lut_tile_3_9_chanxy_out[27];
    assign wire_7646 = lut_tile_3_9_chanxy_out[28];
    assign wire_7648 = lut_tile_3_9_chanxy_out[29];
    assign wire_13921 = lut_tile_3_9_chanxy_out[30];
    assign wire_13929 = lut_tile_3_9_chanxy_out[31];
    assign wire_13937 = lut_tile_3_9_chanxy_out[32];
    assign wire_13945 = lut_tile_3_9_chanxy_out[33];
    assign wire_13953 = lut_tile_3_9_chanxy_out[34];
    assign wire_13961 = lut_tile_3_9_chanxy_out[35];
    assign wire_13969 = lut_tile_3_9_chanxy_out[36];
    assign wire_13977 = lut_tile_3_9_chanxy_out[37];
    assign wire_13985 = lut_tile_3_9_chanxy_out[38];
    assign wire_13993 = lut_tile_3_9_chanxy_out[39];
    assign wire_14001 = lut_tile_3_9_chanxy_out[40];
    assign wire_14009 = lut_tile_3_9_chanxy_out[41];
    assign wire_14017 = lut_tile_3_9_chanxy_out[42];
    assign wire_14025 = lut_tile_3_9_chanxy_out[43];
    assign wire_14033 = lut_tile_3_9_chanxy_out[44];
    assign wire_14070 = lut_tile_3_9_chanxy_out[45];
    assign wire_14072 = lut_tile_3_9_chanxy_out[46];
    assign wire_14074 = lut_tile_3_9_chanxy_out[47];
    assign wire_14076 = lut_tile_3_9_chanxy_out[48];
    assign wire_14078 = lut_tile_3_9_chanxy_out[49];
    assign wire_14080 = lut_tile_3_9_chanxy_out[50];
    assign wire_14082 = lut_tile_3_9_chanxy_out[51];
    assign wire_14084 = lut_tile_3_9_chanxy_out[52];
    assign wire_14086 = lut_tile_3_9_chanxy_out[53];
    assign wire_14088 = lut_tile_3_9_chanxy_out[54];
    assign wire_14090 = lut_tile_3_9_chanxy_out[55];
    assign wire_14092 = lut_tile_3_9_chanxy_out[56];
    assign wire_14094 = lut_tile_3_9_chanxy_out[57];
    assign wire_14096 = lut_tile_3_9_chanxy_out[58];
    assign wire_14098 = lut_tile_3_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_3_10_chanxy_in = {wire_14422, wire_7288, wire_7236, wire_7214, wire_7192, wire_5782, wire_5776, wire_5767, wire_5761, wire_14414, wire_7280, wire_7258, wire_7206, wire_7184, wire_5782, wire_5776, wire_5767, wire_5761, wire_14406, wire_7272, wire_7250, wire_7228, wire_7176, wire_5782, wire_5776, wire_5767, wire_5761, wire_14398, wire_7264, wire_7242, wire_7220, wire_7198, wire_5782, wire_5773, wire_5767, wire_5295, wire_14390, wire_7286, wire_7234, wire_7212, wire_7190, wire_5782, wire_5773, wire_5767, wire_5295, wire_14382, wire_7278, wire_7256, wire_7204, wire_7182, wire_5782, wire_5773, wire_5767, wire_5295, wire_14374, wire_7270, wire_7248, wire_7226, wire_7174, wire_5779, wire_5773, wire_5764, wire_5295, wire_14366, wire_7262, wire_7240, wire_7218, wire_7196, wire_5779, wire_5773, wire_5764, wire_5295, wire_14358, wire_7284, wire_7232, wire_7210, wire_7188, wire_5779, wire_5773, wire_5764, wire_5295, wire_14350, wire_7276, wire_7254, wire_7202, wire_7180, wire_5779, wire_5770, wire_5764, wire_5291, wire_14342, wire_7268, wire_7246, wire_7224, wire_7172, wire_5779, wire_5770, wire_5764, wire_5291, wire_14334, wire_7260, wire_7238, wire_7216, wire_7194, wire_5779, wire_5770, wire_5764, wire_5291, wire_14326, wire_7282, wire_7230, wire_7208, wire_7186, wire_5776, wire_5770, wire_5761, wire_5291, wire_14318, wire_7274, wire_7252, wire_7200, wire_7178, wire_5776, wire_5770, wire_5761, wire_5291, wire_14310, wire_7266, wire_7244, wire_7222, wire_7170, wire_5776, wire_5770, wire_5761, wire_5291, wire_14519, wire_7672, wire_7648, wire_7596, wire_7574, wire_5782, wire_5776, wire_5767, wire_5761, wire_14517, wire_7664, wire_7640, wire_7618, wire_7566, wire_5782, wire_5776, wire_5767, wire_5761, wire_14515, wire_7656, wire_7632, wire_7610, wire_7588, wire_5782, wire_5776, wire_5767, wire_5761, wire_14513, wire_7678, wire_7624, wire_7602, wire_7580, wire_5782, wire_5773, wire_5767, wire_5295, wire_14511, wire_7670, wire_7646, wire_7594, wire_7572, wire_5782, wire_5773, wire_5767, wire_5295, wire_14509, wire_7662, wire_7638, wire_7616, wire_7564, wire_5782, wire_5773, wire_5767, wire_5295, wire_14507, wire_7654, wire_7630, wire_7608, wire_7586, wire_5779, wire_5773, wire_5764, wire_5295, wire_14505, wire_7676, wire_7622, wire_7600, wire_7578, wire_5779, wire_5773, wire_5764, wire_5295, wire_14503, wire_7668, wire_7644, wire_7592, wire_7570, wire_5779, wire_5773, wire_5764, wire_5295, wire_14501, wire_7660, wire_7636, wire_7614, wire_7562, wire_5779, wire_5770, wire_5764, wire_5291, wire_14499, wire_7652, wire_7628, wire_7606, wire_7584, wire_5779, wire_5770, wire_5764, wire_5291, wire_14497, wire_7674, wire_7620, wire_7598, wire_7576, wire_5779, wire_5770, wire_5764, wire_5291, wire_14495, wire_7666, wire_7642, wire_7590, wire_7568, wire_5776, wire_5770, wire_5761, wire_5291, wire_14493, wire_7658, wire_7634, wire_7612, wire_7560, wire_5776, wire_5770, wire_5761, wire_5291, wire_14491, wire_7650, wire_7626, wire_7604, wire_7582, wire_5776, wire_5770, wire_5761, wire_5291, wire_14519, wire_14424, wire_14127, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14032, wire_7558, wire_5334, wire_14419, wire_14418, wire_14125, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_13920, wire_7556, wire_5334, wire_14473, wire_14472, wire_14123, wire_14035, wire_14034, wire_13995, wire_13994, wire_13955, wire_13954, wire_13928, wire_7554, wire_5334, wire_14501, wire_14352, wire_14121, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_13936, wire_7552, wire_5294, wire_14347, wire_14346, wire_14119, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_13944, wire_7550, wire_5294, wire_14485, wire_14484, wire_14117, wire_14027, wire_14026, wire_13987, wire_13986, wire_13952, wire_13947, wire_13946, wire_7548, wire_5294, wire_14513, wire_14400, wire_14115, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_13960, wire_7546, wire_5338, wire_5294, wire_14395, wire_14394, wire_14113, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13968, wire_7544, wire_5338, wire_5294, wire_14467, wire_14466, wire_14111, wire_14019, wire_14018, wire_13979, wire_13978, wire_13976, wire_13939, wire_13938, wire_7542, wire_5338, wire_5294, wire_14495, wire_14328, wire_5338, wire_14109, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_13984, wire_7540, wire_5338, wire_5290, wire_14323, wire_14322, wire_5334, wire_14107, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13992, wire_7538, wire_5338, wire_5290, wire_14479, wire_14478, wire_5334, wire_14105, wire_14011, wire_14010, wire_14000, wire_13971, wire_13970, wire_13931, wire_13930, wire_7536, wire_5338, wire_5290, wire_14507, wire_14376, wire_5294, wire_14103, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14008, wire_7534, wire_5334, wire_5290, wire_14371, wire_14370, wire_5290, wire_14101, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_14016, wire_7532, wire_5334, wire_5290, wire_14461, wire_14460, wire_5290, wire_14129, wire_14024, wire_14003, wire_14002, wire_13963, wire_13962, wire_13923, wire_13922, wire_7530, wire_5334, wire_5290, wire_14459, wire_14458, wire_14489, wire_14488, wire_14503, wire_14360, wire_14441, wire_14440, wire_14471, wire_14470, wire_14515, wire_14408, wire_14453, wire_14452, wire_14483, wire_14482, wire_14497, wire_14336, wire_14435, wire_14434, wire_5338, wire_14465, wire_14464, wire_5338, wire_14509, wire_14384, wire_5334, wire_14447, wire_14446, wire_5294, wire_14477, wire_14476, wire_5294, wire_14491, wire_14312, wire_5290, wire_14427, wire_14426, wire_14363, wire_14362, wire_14517, wire_14416, wire_14355, wire_14354, wire_14411, wire_14410, wire_14499, wire_14344, wire_14403, wire_14402, wire_14339, wire_14338, wire_14511, wire_14392, wire_14331, wire_14330, wire_5338, wire_14387, wire_14386, wire_5338, wire_14493, wire_14320, wire_5334, wire_14379, wire_14378, wire_5294, wire_14315, wire_14314, wire_5294, wire_14505, wire_14368, wire_5290, wire_14443, wire_14442, wire_14457, wire_14456, wire_14487, wire_14486, wire_14455, wire_14454, wire_14439, wire_14438, wire_14469, wire_14468, wire_14437, wire_14436, wire_14451, wire_14450, wire_14481, wire_14480, wire_14449, wire_14448, wire_5338, wire_14433, wire_14432, wire_5334, wire_14463, wire_14462, wire_5334, wire_14431, wire_14430, wire_5294, wire_14445, wire_14444, wire_5290, wire_14475, wire_14474, wire_5290};
    // CHNAXY TOTAL: 573
    assign wire_7561 = lut_tile_3_10_chanxy_out[0];
    assign wire_7563 = lut_tile_3_10_chanxy_out[1];
    assign wire_7565 = lut_tile_3_10_chanxy_out[2];
    assign wire_7567 = lut_tile_3_10_chanxy_out[3];
    assign wire_7569 = lut_tile_3_10_chanxy_out[4];
    assign wire_7571 = lut_tile_3_10_chanxy_out[5];
    assign wire_7573 = lut_tile_3_10_chanxy_out[6];
    assign wire_7575 = lut_tile_3_10_chanxy_out[7];
    assign wire_7577 = lut_tile_3_10_chanxy_out[8];
    assign wire_7579 = lut_tile_3_10_chanxy_out[9];
    assign wire_7581 = lut_tile_3_10_chanxy_out[10];
    assign wire_7583 = lut_tile_3_10_chanxy_out[11];
    assign wire_7585 = lut_tile_3_10_chanxy_out[12];
    assign wire_7587 = lut_tile_3_10_chanxy_out[13];
    assign wire_7589 = lut_tile_3_10_chanxy_out[14];
    assign wire_7591 = lut_tile_3_10_chanxy_out[15];
    assign wire_7593 = lut_tile_3_10_chanxy_out[16];
    assign wire_7595 = lut_tile_3_10_chanxy_out[17];
    assign wire_7597 = lut_tile_3_10_chanxy_out[18];
    assign wire_7599 = lut_tile_3_10_chanxy_out[19];
    assign wire_7601 = lut_tile_3_10_chanxy_out[20];
    assign wire_7603 = lut_tile_3_10_chanxy_out[21];
    assign wire_7605 = lut_tile_3_10_chanxy_out[22];
    assign wire_7607 = lut_tile_3_10_chanxy_out[23];
    assign wire_7609 = lut_tile_3_10_chanxy_out[24];
    assign wire_7611 = lut_tile_3_10_chanxy_out[25];
    assign wire_7613 = lut_tile_3_10_chanxy_out[26];
    assign wire_7615 = lut_tile_3_10_chanxy_out[27];
    assign wire_7617 = lut_tile_3_10_chanxy_out[28];
    assign wire_7619 = lut_tile_3_10_chanxy_out[29];
    assign wire_7621 = lut_tile_3_10_chanxy_out[30];
    assign wire_7623 = lut_tile_3_10_chanxy_out[31];
    assign wire_7625 = lut_tile_3_10_chanxy_out[32];
    assign wire_7627 = lut_tile_3_10_chanxy_out[33];
    assign wire_7629 = lut_tile_3_10_chanxy_out[34];
    assign wire_7631 = lut_tile_3_10_chanxy_out[35];
    assign wire_7633 = lut_tile_3_10_chanxy_out[36];
    assign wire_7635 = lut_tile_3_10_chanxy_out[37];
    assign wire_7637 = lut_tile_3_10_chanxy_out[38];
    assign wire_7639 = lut_tile_3_10_chanxy_out[39];
    assign wire_7641 = lut_tile_3_10_chanxy_out[40];
    assign wire_7643 = lut_tile_3_10_chanxy_out[41];
    assign wire_7645 = lut_tile_3_10_chanxy_out[42];
    assign wire_7647 = lut_tile_3_10_chanxy_out[43];
    assign wire_7649 = lut_tile_3_10_chanxy_out[44];
    assign wire_7650 = lut_tile_3_10_chanxy_out[45];
    assign wire_7651 = lut_tile_3_10_chanxy_out[46];
    assign wire_7652 = lut_tile_3_10_chanxy_out[47];
    assign wire_7653 = lut_tile_3_10_chanxy_out[48];
    assign wire_7654 = lut_tile_3_10_chanxy_out[49];
    assign wire_7655 = lut_tile_3_10_chanxy_out[50];
    assign wire_7656 = lut_tile_3_10_chanxy_out[51];
    assign wire_7657 = lut_tile_3_10_chanxy_out[52];
    assign wire_7658 = lut_tile_3_10_chanxy_out[53];
    assign wire_7659 = lut_tile_3_10_chanxy_out[54];
    assign wire_7660 = lut_tile_3_10_chanxy_out[55];
    assign wire_7661 = lut_tile_3_10_chanxy_out[56];
    assign wire_7662 = lut_tile_3_10_chanxy_out[57];
    assign wire_7663 = lut_tile_3_10_chanxy_out[58];
    assign wire_7664 = lut_tile_3_10_chanxy_out[59];
    assign wire_7665 = lut_tile_3_10_chanxy_out[60];
    assign wire_7666 = lut_tile_3_10_chanxy_out[61];
    assign wire_7667 = lut_tile_3_10_chanxy_out[62];
    assign wire_7668 = lut_tile_3_10_chanxy_out[63];
    assign wire_7669 = lut_tile_3_10_chanxy_out[64];
    assign wire_7670 = lut_tile_3_10_chanxy_out[65];
    assign wire_7671 = lut_tile_3_10_chanxy_out[66];
    assign wire_7672 = lut_tile_3_10_chanxy_out[67];
    assign wire_7673 = lut_tile_3_10_chanxy_out[68];
    assign wire_7674 = lut_tile_3_10_chanxy_out[69];
    assign wire_7675 = lut_tile_3_10_chanxy_out[70];
    assign wire_7676 = lut_tile_3_10_chanxy_out[71];
    assign wire_7677 = lut_tile_3_10_chanxy_out[72];
    assign wire_7678 = lut_tile_3_10_chanxy_out[73];
    assign wire_7679 = lut_tile_3_10_chanxy_out[74];
    assign wire_14313 = lut_tile_3_10_chanxy_out[75];
    assign wire_14321 = lut_tile_3_10_chanxy_out[76];
    assign wire_14329 = lut_tile_3_10_chanxy_out[77];
    assign wire_14337 = lut_tile_3_10_chanxy_out[78];
    assign wire_14345 = lut_tile_3_10_chanxy_out[79];
    assign wire_14353 = lut_tile_3_10_chanxy_out[80];
    assign wire_14361 = lut_tile_3_10_chanxy_out[81];
    assign wire_14369 = lut_tile_3_10_chanxy_out[82];
    assign wire_14377 = lut_tile_3_10_chanxy_out[83];
    assign wire_14385 = lut_tile_3_10_chanxy_out[84];
    assign wire_14393 = lut_tile_3_10_chanxy_out[85];
    assign wire_14401 = lut_tile_3_10_chanxy_out[86];
    assign wire_14409 = lut_tile_3_10_chanxy_out[87];
    assign wire_14417 = lut_tile_3_10_chanxy_out[88];
    assign wire_14425 = lut_tile_3_10_chanxy_out[89];
    assign wire_14460 = lut_tile_3_10_chanxy_out[90];
    assign wire_14462 = lut_tile_3_10_chanxy_out[91];
    assign wire_14464 = lut_tile_3_10_chanxy_out[92];
    assign wire_14466 = lut_tile_3_10_chanxy_out[93];
    assign wire_14468 = lut_tile_3_10_chanxy_out[94];
    assign wire_14470 = lut_tile_3_10_chanxy_out[95];
    assign wire_14472 = lut_tile_3_10_chanxy_out[96];
    assign wire_14474 = lut_tile_3_10_chanxy_out[97];
    assign wire_14476 = lut_tile_3_10_chanxy_out[98];
    assign wire_14478 = lut_tile_3_10_chanxy_out[99];
    assign wire_14480 = lut_tile_3_10_chanxy_out[100];
    assign wire_14482 = lut_tile_3_10_chanxy_out[101];
    assign wire_14484 = lut_tile_3_10_chanxy_out[102];
    assign wire_14486 = lut_tile_3_10_chanxy_out[103];
    assign wire_14488 = lut_tile_3_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_4_1_chanxy_in = {wire_10912, wire_7411, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7298, wire_1203, wire_10904, wire_7439, wire_7407, wire_7406, wire_7367, wire_7366, wire_7327, wire_7326, wire_7306, wire_1203, wire_10896, wire_7437, wire_7405, wire_7404, wire_7365, wire_7364, wire_7325, wire_7324, wire_7314, wire_1203, wire_10888, wire_7435, wire_7401, wire_7400, wire_7361, wire_7360, wire_7322, wire_7321, wire_7320, wire_693, wire_10880, wire_7433, wire_7399, wire_7398, wire_7359, wire_7358, wire_7330, wire_7319, wire_7318, wire_693, wire_10872, wire_7431, wire_7397, wire_7396, wire_7357, wire_7356, wire_7338, wire_7317, wire_7316, wire_693, wire_10864, wire_7429, wire_7393, wire_7392, wire_7353, wire_7352, wire_7346, wire_7313, wire_7312, wire_1207, wire_693, wire_10856, wire_7427, wire_7391, wire_7390, wire_7354, wire_7351, wire_7350, wire_7311, wire_7310, wire_1207, wire_693, wire_10848, wire_7425, wire_7389, wire_7388, wire_7362, wire_7349, wire_7348, wire_7309, wire_7308, wire_1207, wire_693, wire_10840, wire_7423, wire_7385, wire_7384, wire_7370, wire_7345, wire_7344, wire_7305, wire_7304, wire_1207, wire_689, wire_10832, wire_7421, wire_7383, wire_7382, wire_7378, wire_7343, wire_7342, wire_7303, wire_7302, wire_1207, wire_689, wire_10824, wire_7419, wire_7386, wire_7381, wire_7380, wire_7341, wire_7340, wire_7301, wire_7300, wire_1207, wire_689, wire_10816, wire_7417, wire_7394, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296, wire_1203, wire_689, wire_10808, wire_7415, wire_7402, wire_7375, wire_7374, wire_7335, wire_7334, wire_7295, wire_7294, wire_1203, wire_689, wire_10800, wire_7413, wire_7373, wire_7372, wire_7333, wire_7332, wire_7293, wire_7292, wire_7290, wire_1203, wire_689, wire_11039, wire_7829, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_7682, wire_1203, wire_11037, wire_7801, wire_7797, wire_7796, wire_7794, wire_7757, wire_7756, wire_7717, wire_7716, wire_1203, wire_11035, wire_7803, wire_7793, wire_7792, wire_7786, wire_7753, wire_7752, wire_7713, wire_7712, wire_1203, wire_11033, wire_7805, wire_7791, wire_7790, wire_7778, wire_7751, wire_7750, wire_7711, wire_7710, wire_693, wire_11031, wire_7807, wire_7789, wire_7788, wire_7770, wire_7749, wire_7748, wire_7709, wire_7708, wire_693, wire_11029, wire_7809, wire_7785, wire_7784, wire_7762, wire_7745, wire_7744, wire_7705, wire_7704, wire_693, wire_11027, wire_7811, wire_7783, wire_7782, wire_7754, wire_7743, wire_7742, wire_7703, wire_7702, wire_1207, wire_693, wire_11025, wire_7813, wire_7781, wire_7780, wire_7746, wire_7741, wire_7740, wire_7701, wire_7700, wire_1207, wire_693, wire_11023, wire_7815, wire_7777, wire_7776, wire_7738, wire_7737, wire_7736, wire_7697, wire_7696, wire_1207, wire_693, wire_11021, wire_7817, wire_7775, wire_7774, wire_7735, wire_7734, wire_7730, wire_7695, wire_7694, wire_1207, wire_689, wire_11019, wire_7819, wire_7773, wire_7772, wire_7733, wire_7732, wire_7722, wire_7693, wire_7692, wire_1207, wire_689, wire_11017, wire_7821, wire_7769, wire_7768, wire_7729, wire_7728, wire_7714, wire_7689, wire_7688, wire_1207, wire_689, wire_11015, wire_7823, wire_7767, wire_7766, wire_7727, wire_7726, wire_7706, wire_7687, wire_7686, wire_1203, wire_689, wire_11013, wire_7825, wire_7765, wire_7764, wire_7725, wire_7724, wire_7698, wire_7685, wire_7684, wire_1203, wire_689, wire_11011, wire_7827, wire_7761, wire_7760, wire_7721, wire_7720, wire_7690, wire_7681, wire_7680, wire_1203, wire_689, wire_10603, wire_10602, wire_10619, wire_10618, wire_11013, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10906, wire_7829, wire_732, wire_10589, wire_10588, wire_10573, wire_10572, wire_10559, wire_10558, wire_10649, wire_10522, wire_11015, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10898, wire_7827, wire_732, wire_10543, wire_10542, wire_10617, wire_10616, wire_10587, wire_10586, wire_10633, wire_10458, wire_11017, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10890, wire_7825, wire_732, wire_10557, wire_10556, wire_10647, wire_10514, wire_10615, wire_10614, wire_10601, wire_10600, wire_11019, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10882, wire_7823, wire_692, wire_10571, wire_10570, wire_10585, wire_10584, wire_10541, wire_10540, wire_10631, wire_10450, wire_11021, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10874, wire_7821, wire_692, wire_10555, wire_10554, wire_10599, wire_10598, wire_10569, wire_10568, wire_10645, wire_10506, wire_11023, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10866, wire_7819, wire_692, wire_10539, wire_10538, wire_10629, wire_10442, wire_10597, wire_10596, wire_10613, wire_10612, wire_11025, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10858, wire_7817, wire_736, wire_692, wire_10583, wire_10582, wire_10567, wire_10566, wire_10553, wire_10552, wire_10643, wire_10498, wire_11027, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10850, wire_7815, wire_736, wire_692, wire_10537, wire_10536, wire_10611, wire_10610, wire_10581, wire_10580, wire_10627, wire_10434, wire_11029, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10842, wire_7813, wire_736, wire_692, wire_10551, wire_10550, wire_10641, wire_10490, wire_10609, wire_10608, wire_736, wire_10595, wire_10594, wire_736, wire_11031, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10834, wire_7811, wire_736, wire_688, wire_10565, wire_10564, wire_736, wire_10579, wire_10578, wire_736, wire_10535, wire_10534, wire_736, wire_10625, wire_10426, wire_736, wire_11033, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10826, wire_7809, wire_736, wire_688, wire_10549, wire_10548, wire_732, wire_10593, wire_10592, wire_732, wire_10563, wire_10562, wire_732, wire_10639, wire_10482, wire_732, wire_11035, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10818, wire_7807, wire_736, wire_688, wire_10533, wire_10532, wire_732, wire_10623, wire_10418, wire_732, wire_10591, wire_10590, wire_692, wire_10607, wire_10606, wire_692, wire_11037, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10810, wire_7805, wire_732, wire_688, wire_10577, wire_10576, wire_692, wire_10561, wire_10560, wire_692, wire_10547, wire_10546, wire_692, wire_10637, wire_10474, wire_692, wire_11039, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10802, wire_7803, wire_732, wire_688, wire_10531, wire_10530, wire_688, wire_10605, wire_10604, wire_688, wire_10575, wire_10574, wire_688, wire_10621, wire_10410, wire_688, wire_11011, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10914, wire_7801, wire_732, wire_688, wire_10545, wire_10544, wire_688, wire_10635, wire_10466, wire_688};
    // CHNAXY TOTAL: 621
    assign wire_7680 = lut_tile_4_1_chanxy_out[0];
    assign wire_7682 = lut_tile_4_1_chanxy_out[1];
    assign wire_7683 = lut_tile_4_1_chanxy_out[2];
    assign wire_7684 = lut_tile_4_1_chanxy_out[3];
    assign wire_7686 = lut_tile_4_1_chanxy_out[4];
    assign wire_7688 = lut_tile_4_1_chanxy_out[5];
    assign wire_7690 = lut_tile_4_1_chanxy_out[6];
    assign wire_7691 = lut_tile_4_1_chanxy_out[7];
    assign wire_7692 = lut_tile_4_1_chanxy_out[8];
    assign wire_7694 = lut_tile_4_1_chanxy_out[9];
    assign wire_7696 = lut_tile_4_1_chanxy_out[10];
    assign wire_7698 = lut_tile_4_1_chanxy_out[11];
    assign wire_7699 = lut_tile_4_1_chanxy_out[12];
    assign wire_7700 = lut_tile_4_1_chanxy_out[13];
    assign wire_7702 = lut_tile_4_1_chanxy_out[14];
    assign wire_7704 = lut_tile_4_1_chanxy_out[15];
    assign wire_7706 = lut_tile_4_1_chanxy_out[16];
    assign wire_7707 = lut_tile_4_1_chanxy_out[17];
    assign wire_7708 = lut_tile_4_1_chanxy_out[18];
    assign wire_7710 = lut_tile_4_1_chanxy_out[19];
    assign wire_7712 = lut_tile_4_1_chanxy_out[20];
    assign wire_7714 = lut_tile_4_1_chanxy_out[21];
    assign wire_7715 = lut_tile_4_1_chanxy_out[22];
    assign wire_7716 = lut_tile_4_1_chanxy_out[23];
    assign wire_7718 = lut_tile_4_1_chanxy_out[24];
    assign wire_7720 = lut_tile_4_1_chanxy_out[25];
    assign wire_7722 = lut_tile_4_1_chanxy_out[26];
    assign wire_7723 = lut_tile_4_1_chanxy_out[27];
    assign wire_7724 = lut_tile_4_1_chanxy_out[28];
    assign wire_7726 = lut_tile_4_1_chanxy_out[29];
    assign wire_7728 = lut_tile_4_1_chanxy_out[30];
    assign wire_7730 = lut_tile_4_1_chanxy_out[31];
    assign wire_7731 = lut_tile_4_1_chanxy_out[32];
    assign wire_7732 = lut_tile_4_1_chanxy_out[33];
    assign wire_7734 = lut_tile_4_1_chanxy_out[34];
    assign wire_7736 = lut_tile_4_1_chanxy_out[35];
    assign wire_7738 = lut_tile_4_1_chanxy_out[36];
    assign wire_7739 = lut_tile_4_1_chanxy_out[37];
    assign wire_7740 = lut_tile_4_1_chanxy_out[38];
    assign wire_7742 = lut_tile_4_1_chanxy_out[39];
    assign wire_7744 = lut_tile_4_1_chanxy_out[40];
    assign wire_7746 = lut_tile_4_1_chanxy_out[41];
    assign wire_7747 = lut_tile_4_1_chanxy_out[42];
    assign wire_7748 = lut_tile_4_1_chanxy_out[43];
    assign wire_7750 = lut_tile_4_1_chanxy_out[44];
    assign wire_7752 = lut_tile_4_1_chanxy_out[45];
    assign wire_7754 = lut_tile_4_1_chanxy_out[46];
    assign wire_7755 = lut_tile_4_1_chanxy_out[47];
    assign wire_7756 = lut_tile_4_1_chanxy_out[48];
    assign wire_7758 = lut_tile_4_1_chanxy_out[49];
    assign wire_7760 = lut_tile_4_1_chanxy_out[50];
    assign wire_7762 = lut_tile_4_1_chanxy_out[51];
    assign wire_7763 = lut_tile_4_1_chanxy_out[52];
    assign wire_7764 = lut_tile_4_1_chanxy_out[53];
    assign wire_7766 = lut_tile_4_1_chanxy_out[54];
    assign wire_7768 = lut_tile_4_1_chanxy_out[55];
    assign wire_7770 = lut_tile_4_1_chanxy_out[56];
    assign wire_7771 = lut_tile_4_1_chanxy_out[57];
    assign wire_7772 = lut_tile_4_1_chanxy_out[58];
    assign wire_7774 = lut_tile_4_1_chanxy_out[59];
    assign wire_7776 = lut_tile_4_1_chanxy_out[60];
    assign wire_7778 = lut_tile_4_1_chanxy_out[61];
    assign wire_7779 = lut_tile_4_1_chanxy_out[62];
    assign wire_7780 = lut_tile_4_1_chanxy_out[63];
    assign wire_7782 = lut_tile_4_1_chanxy_out[64];
    assign wire_7784 = lut_tile_4_1_chanxy_out[65];
    assign wire_7786 = lut_tile_4_1_chanxy_out[66];
    assign wire_7787 = lut_tile_4_1_chanxy_out[67];
    assign wire_7788 = lut_tile_4_1_chanxy_out[68];
    assign wire_7790 = lut_tile_4_1_chanxy_out[69];
    assign wire_7792 = lut_tile_4_1_chanxy_out[70];
    assign wire_7794 = lut_tile_4_1_chanxy_out[71];
    assign wire_7795 = lut_tile_4_1_chanxy_out[72];
    assign wire_7796 = lut_tile_4_1_chanxy_out[73];
    assign wire_7798 = lut_tile_4_1_chanxy_out[74];
    assign wire_10803 = lut_tile_4_1_chanxy_out[75];
    assign wire_10811 = lut_tile_4_1_chanxy_out[76];
    assign wire_10819 = lut_tile_4_1_chanxy_out[77];
    assign wire_10827 = lut_tile_4_1_chanxy_out[78];
    assign wire_10835 = lut_tile_4_1_chanxy_out[79];
    assign wire_10843 = lut_tile_4_1_chanxy_out[80];
    assign wire_10851 = lut_tile_4_1_chanxy_out[81];
    assign wire_10859 = lut_tile_4_1_chanxy_out[82];
    assign wire_10867 = lut_tile_4_1_chanxy_out[83];
    assign wire_10875 = lut_tile_4_1_chanxy_out[84];
    assign wire_10883 = lut_tile_4_1_chanxy_out[85];
    assign wire_10891 = lut_tile_4_1_chanxy_out[86];
    assign wire_10899 = lut_tile_4_1_chanxy_out[87];
    assign wire_10907 = lut_tile_4_1_chanxy_out[88];
    assign wire_10915 = lut_tile_4_1_chanxy_out[89];
    assign wire_10980 = lut_tile_4_1_chanxy_out[90];
    assign wire_10982 = lut_tile_4_1_chanxy_out[91];
    assign wire_10984 = lut_tile_4_1_chanxy_out[92];
    assign wire_10986 = lut_tile_4_1_chanxy_out[93];
    assign wire_10988 = lut_tile_4_1_chanxy_out[94];
    assign wire_10990 = lut_tile_4_1_chanxy_out[95];
    assign wire_10992 = lut_tile_4_1_chanxy_out[96];
    assign wire_10994 = lut_tile_4_1_chanxy_out[97];
    assign wire_10996 = lut_tile_4_1_chanxy_out[98];
    assign wire_10998 = lut_tile_4_1_chanxy_out[99];
    assign wire_11000 = lut_tile_4_1_chanxy_out[100];
    assign wire_11002 = lut_tile_4_1_chanxy_out[101];
    assign wire_11004 = lut_tile_4_1_chanxy_out[102];
    assign wire_11006 = lut_tile_4_1_chanxy_out[103];
    assign wire_11008 = lut_tile_4_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_4_2_chanxy_in = {wire_11304, wire_7441, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7300, wire_1719, wire_11296, wire_7469, wire_7407, wire_7406, wire_7367, wire_7366, wire_7327, wire_7326, wire_7308, wire_1719, wire_11288, wire_7467, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7316, wire_1719, wire_11280, wire_7465, wire_7401, wire_7400, wire_7361, wire_7360, wire_7324, wire_7321, wire_7320, wire_1209, wire_11272, wire_7463, wire_7399, wire_7398, wire_7359, wire_7358, wire_7332, wire_7319, wire_7318, wire_1209, wire_11264, wire_7461, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7340, wire_1209, wire_11256, wire_7459, wire_7393, wire_7392, wire_7353, wire_7352, wire_7348, wire_7313, wire_7312, wire_1723, wire_1209, wire_11248, wire_7457, wire_7391, wire_7390, wire_7356, wire_7351, wire_7350, wire_7311, wire_7310, wire_1723, wire_1209, wire_11240, wire_7455, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7364, wire_1723, wire_1209, wire_11232, wire_7453, wire_7385, wire_7384, wire_7372, wire_7345, wire_7344, wire_7305, wire_7304, wire_1723, wire_1205, wire_11224, wire_7451, wire_7383, wire_7382, wire_7380, wire_7343, wire_7342, wire_7303, wire_7302, wire_1723, wire_1205, wire_11216, wire_7449, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7388, wire_1723, wire_1205, wire_11208, wire_7447, wire_7396, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296, wire_1719, wire_1205, wire_11200, wire_7445, wire_7404, wire_7375, wire_7374, wire_7335, wire_7334, wire_7295, wire_7294, wire_1719, wire_1205, wire_11192, wire_7443, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7292, wire_1719, wire_1205, wire_11429, wire_7859, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_7684, wire_1719, wire_11427, wire_7831, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7796, wire_1719, wire_11425, wire_7833, wire_7793, wire_7792, wire_7788, wire_7753, wire_7752, wire_7713, wire_7712, wire_1719, wire_11423, wire_7835, wire_7791, wire_7790, wire_7780, wire_7751, wire_7750, wire_7711, wire_7710, wire_1209, wire_11421, wire_7837, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7772, wire_1209, wire_11419, wire_7839, wire_7785, wire_7784, wire_7764, wire_7745, wire_7744, wire_7705, wire_7704, wire_1209, wire_11417, wire_7841, wire_7783, wire_7782, wire_7756, wire_7743, wire_7742, wire_7703, wire_7702, wire_1723, wire_1209, wire_11415, wire_7843, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7748, wire_1723, wire_1209, wire_11413, wire_7845, wire_7777, wire_7776, wire_7740, wire_7737, wire_7736, wire_7697, wire_7696, wire_1723, wire_1209, wire_11411, wire_7847, wire_7775, wire_7774, wire_7735, wire_7734, wire_7732, wire_7695, wire_7694, wire_1723, wire_1205, wire_11409, wire_7849, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7724, wire_1723, wire_1205, wire_11407, wire_7851, wire_7769, wire_7768, wire_7729, wire_7728, wire_7716, wire_7689, wire_7688, wire_1723, wire_1205, wire_11405, wire_7853, wire_7767, wire_7766, wire_7727, wire_7726, wire_7708, wire_7687, wire_7686, wire_1719, wire_1205, wire_11403, wire_7855, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7700, wire_1719, wire_1205, wire_11401, wire_7857, wire_7761, wire_7760, wire_7721, wire_7720, wire_7692, wire_7681, wire_7680, wire_1719, wire_1205, wire_11037, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10914, wire_7794, wire_1248, wire_11035, wire_10949, wire_10948, wire_10939, wire_10938, wire_10929, wire_10928, wire_10802, wire_7786, wire_1248, wire_11033, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10810, wire_7778, wire_1248, wire_11031, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10818, wire_7770, wire_1208, wire_11029, wire_10947, wire_10946, wire_10937, wire_10936, wire_10927, wire_10926, wire_10826, wire_7762, wire_1208, wire_11027, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10834, wire_7754, wire_1208, wire_11025, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10842, wire_7746, wire_1252, wire_1208, wire_11023, wire_10945, wire_10944, wire_10935, wire_10934, wire_10925, wire_10924, wire_10850, wire_7738, wire_1252, wire_1208, wire_11021, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10858, wire_7730, wire_1252, wire_1208, wire_11019, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10866, wire_7722, wire_1252, wire_1204, wire_11017, wire_10943, wire_10942, wire_10933, wire_10932, wire_10923, wire_10922, wire_10874, wire_7714, wire_1252, wire_1204, wire_11015, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10882, wire_7706, wire_1252, wire_1204, wire_11013, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10890, wire_7698, wire_1248, wire_1204, wire_11011, wire_10941, wire_10940, wire_10931, wire_10930, wire_10921, wire_10920, wire_10898, wire_7690, wire_1248, wire_1204, wire_11039, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10906, wire_7682, wire_1248, wire_1204, wire_11403, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11298, wire_7859, wire_1248, wire_11405, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11290, wire_7857, wire_1248, wire_11407, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11282, wire_7855, wire_1248, wire_11409, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11274, wire_7853, wire_1208, wire_11411, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11266, wire_7851, wire_1208, wire_11413, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11258, wire_7849, wire_1208, wire_11415, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11250, wire_7847, wire_1252, wire_1208, wire_11417, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11242, wire_7845, wire_1252, wire_1208, wire_11419, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11234, wire_7843, wire_1252, wire_1208, wire_11421, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11226, wire_7841, wire_1252, wire_1204, wire_11423, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11218, wire_7839, wire_1252, wire_1204, wire_11425, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11210, wire_7837, wire_1252, wire_1204, wire_11427, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11202, wire_7835, wire_1248, wire_1204, wire_11429, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11194, wire_7833, wire_1248, wire_1204, wire_11401, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11306, wire_7831, wire_1248, wire_1204};
    // CHNAXY TOTAL: 636
    assign wire_7685 = lut_tile_4_2_chanxy_out[0];
    assign wire_7693 = lut_tile_4_2_chanxy_out[1];
    assign wire_7701 = lut_tile_4_2_chanxy_out[2];
    assign wire_7709 = lut_tile_4_2_chanxy_out[3];
    assign wire_7717 = lut_tile_4_2_chanxy_out[4];
    assign wire_7725 = lut_tile_4_2_chanxy_out[5];
    assign wire_7733 = lut_tile_4_2_chanxy_out[6];
    assign wire_7741 = lut_tile_4_2_chanxy_out[7];
    assign wire_7749 = lut_tile_4_2_chanxy_out[8];
    assign wire_7757 = lut_tile_4_2_chanxy_out[9];
    assign wire_7765 = lut_tile_4_2_chanxy_out[10];
    assign wire_7773 = lut_tile_4_2_chanxy_out[11];
    assign wire_7781 = lut_tile_4_2_chanxy_out[12];
    assign wire_7789 = lut_tile_4_2_chanxy_out[13];
    assign wire_7797 = lut_tile_4_2_chanxy_out[14];
    assign wire_7800 = lut_tile_4_2_chanxy_out[15];
    assign wire_7802 = lut_tile_4_2_chanxy_out[16];
    assign wire_7804 = lut_tile_4_2_chanxy_out[17];
    assign wire_7806 = lut_tile_4_2_chanxy_out[18];
    assign wire_7808 = lut_tile_4_2_chanxy_out[19];
    assign wire_7810 = lut_tile_4_2_chanxy_out[20];
    assign wire_7812 = lut_tile_4_2_chanxy_out[21];
    assign wire_7814 = lut_tile_4_2_chanxy_out[22];
    assign wire_7816 = lut_tile_4_2_chanxy_out[23];
    assign wire_7818 = lut_tile_4_2_chanxy_out[24];
    assign wire_7820 = lut_tile_4_2_chanxy_out[25];
    assign wire_7822 = lut_tile_4_2_chanxy_out[26];
    assign wire_7824 = lut_tile_4_2_chanxy_out[27];
    assign wire_7826 = lut_tile_4_2_chanxy_out[28];
    assign wire_7828 = lut_tile_4_2_chanxy_out[29];
    assign wire_11195 = lut_tile_4_2_chanxy_out[30];
    assign wire_11203 = lut_tile_4_2_chanxy_out[31];
    assign wire_11211 = lut_tile_4_2_chanxy_out[32];
    assign wire_11219 = lut_tile_4_2_chanxy_out[33];
    assign wire_11227 = lut_tile_4_2_chanxy_out[34];
    assign wire_11235 = lut_tile_4_2_chanxy_out[35];
    assign wire_11243 = lut_tile_4_2_chanxy_out[36];
    assign wire_11251 = lut_tile_4_2_chanxy_out[37];
    assign wire_11259 = lut_tile_4_2_chanxy_out[38];
    assign wire_11267 = lut_tile_4_2_chanxy_out[39];
    assign wire_11275 = lut_tile_4_2_chanxy_out[40];
    assign wire_11283 = lut_tile_4_2_chanxy_out[41];
    assign wire_11291 = lut_tile_4_2_chanxy_out[42];
    assign wire_11299 = lut_tile_4_2_chanxy_out[43];
    assign wire_11307 = lut_tile_4_2_chanxy_out[44];
    assign wire_11370 = lut_tile_4_2_chanxy_out[45];
    assign wire_11372 = lut_tile_4_2_chanxy_out[46];
    assign wire_11374 = lut_tile_4_2_chanxy_out[47];
    assign wire_11376 = lut_tile_4_2_chanxy_out[48];
    assign wire_11378 = lut_tile_4_2_chanxy_out[49];
    assign wire_11380 = lut_tile_4_2_chanxy_out[50];
    assign wire_11382 = lut_tile_4_2_chanxy_out[51];
    assign wire_11384 = lut_tile_4_2_chanxy_out[52];
    assign wire_11386 = lut_tile_4_2_chanxy_out[53];
    assign wire_11388 = lut_tile_4_2_chanxy_out[54];
    assign wire_11390 = lut_tile_4_2_chanxy_out[55];
    assign wire_11392 = lut_tile_4_2_chanxy_out[56];
    assign wire_11394 = lut_tile_4_2_chanxy_out[57];
    assign wire_11396 = lut_tile_4_2_chanxy_out[58];
    assign wire_11398 = lut_tile_4_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_3_chanxy_in = {wire_11696, wire_7471, wire_7409, wire_7408, wire_7369, wire_7368, wire_7329, wire_7328, wire_7302, wire_2235, wire_11688, wire_7499, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7310, wire_2235, wire_11680, wire_7497, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7318, wire_2235, wire_11672, wire_7495, wire_7401, wire_7400, wire_7361, wire_7360, wire_7326, wire_7321, wire_7320, wire_1725, wire_11664, wire_7493, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7334, wire_1725, wire_11656, wire_7491, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7342, wire_1725, wire_11648, wire_7489, wire_7393, wire_7392, wire_7353, wire_7352, wire_7350, wire_7313, wire_7312, wire_2239, wire_1725, wire_11640, wire_7487, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7358, wire_2239, wire_1725, wire_11632, wire_7485, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7366, wire_2239, wire_1725, wire_11624, wire_7483, wire_7385, wire_7384, wire_7374, wire_7345, wire_7344, wire_7305, wire_7304, wire_2239, wire_1721, wire_11616, wire_7481, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7382, wire_2239, wire_1721, wire_11608, wire_7479, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7390, wire_2239, wire_1721, wire_11600, wire_7477, wire_7398, wire_7377, wire_7376, wire_7337, wire_7336, wire_7297, wire_7296, wire_2235, wire_1721, wire_11592, wire_7475, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7406, wire_2235, wire_1721, wire_11584, wire_7473, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7294, wire_2235, wire_1721, wire_11819, wire_7889, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7686, wire_2235, wire_11817, wire_7861, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7798, wire_2235, wire_11815, wire_7863, wire_7793, wire_7792, wire_7790, wire_7753, wire_7752, wire_7713, wire_7712, wire_2235, wire_11813, wire_7865, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7782, wire_1725, wire_11811, wire_7867, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7774, wire_1725, wire_11809, wire_7869, wire_7785, wire_7784, wire_7766, wire_7745, wire_7744, wire_7705, wire_7704, wire_1725, wire_11807, wire_7871, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7758, wire_2239, wire_1725, wire_11805, wire_7873, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7750, wire_2239, wire_1725, wire_11803, wire_7875, wire_7777, wire_7776, wire_7742, wire_7737, wire_7736, wire_7697, wire_7696, wire_2239, wire_1725, wire_11801, wire_7877, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7734, wire_2239, wire_1721, wire_11799, wire_7879, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7726, wire_2239, wire_1721, wire_11797, wire_7881, wire_7769, wire_7768, wire_7729, wire_7728, wire_7718, wire_7689, wire_7688, wire_2239, wire_1721, wire_11795, wire_7883, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7710, wire_2235, wire_1721, wire_11793, wire_7885, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7702, wire_2235, wire_1721, wire_11791, wire_7887, wire_7761, wire_7760, wire_7721, wire_7720, wire_7694, wire_7681, wire_7680, wire_2235, wire_1721, wire_11427, wire_11339, wire_11338, wire_11329, wire_11328, wire_11319, wire_11318, wire_11306, wire_7796, wire_1764, wire_11425, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11194, wire_7788, wire_1764, wire_11423, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11202, wire_7780, wire_1764, wire_11421, wire_11337, wire_11336, wire_11327, wire_11326, wire_11317, wire_11316, wire_11210, wire_7772, wire_1724, wire_11419, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11218, wire_7764, wire_1724, wire_11417, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11226, wire_7756, wire_1724, wire_11415, wire_11335, wire_11334, wire_11325, wire_11324, wire_11315, wire_11314, wire_11234, wire_7748, wire_1768, wire_1724, wire_11413, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11242, wire_7740, wire_1768, wire_1724, wire_11411, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11250, wire_7732, wire_1768, wire_1724, wire_11409, wire_11333, wire_11332, wire_11323, wire_11322, wire_11313, wire_11312, wire_11258, wire_7724, wire_1768, wire_1720, wire_11407, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11266, wire_7716, wire_1768, wire_1720, wire_11405, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11274, wire_7708, wire_1768, wire_1720, wire_11403, wire_11331, wire_11330, wire_11321, wire_11320, wire_11311, wire_11310, wire_11282, wire_7700, wire_1764, wire_1720, wire_11401, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11290, wire_7692, wire_1764, wire_1720, wire_11429, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11298, wire_7684, wire_1764, wire_1720, wire_11793, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11690, wire_7889, wire_1764, wire_11795, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11682, wire_7887, wire_1764, wire_11797, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11674, wire_7885, wire_1764, wire_11799, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11666, wire_7883, wire_1724, wire_11801, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11658, wire_7881, wire_1724, wire_11803, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11650, wire_7879, wire_1724, wire_11805, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11642, wire_7877, wire_1768, wire_1724, wire_11807, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11634, wire_7875, wire_1768, wire_1724, wire_11809, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11626, wire_7873, wire_1768, wire_1724, wire_11811, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11618, wire_7871, wire_1768, wire_1720, wire_11813, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11610, wire_7869, wire_1768, wire_1720, wire_11815, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11602, wire_7867, wire_1768, wire_1720, wire_11817, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11594, wire_7865, wire_1764, wire_1720, wire_11819, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11586, wire_7863, wire_1764, wire_1720, wire_11791, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11698, wire_7861, wire_1764, wire_1720};
    // CHNAXY TOTAL: 636
    assign wire_7687 = lut_tile_4_3_chanxy_out[0];
    assign wire_7695 = lut_tile_4_3_chanxy_out[1];
    assign wire_7703 = lut_tile_4_3_chanxy_out[2];
    assign wire_7711 = lut_tile_4_3_chanxy_out[3];
    assign wire_7719 = lut_tile_4_3_chanxy_out[4];
    assign wire_7727 = lut_tile_4_3_chanxy_out[5];
    assign wire_7735 = lut_tile_4_3_chanxy_out[6];
    assign wire_7743 = lut_tile_4_3_chanxy_out[7];
    assign wire_7751 = lut_tile_4_3_chanxy_out[8];
    assign wire_7759 = lut_tile_4_3_chanxy_out[9];
    assign wire_7767 = lut_tile_4_3_chanxy_out[10];
    assign wire_7775 = lut_tile_4_3_chanxy_out[11];
    assign wire_7783 = lut_tile_4_3_chanxy_out[12];
    assign wire_7791 = lut_tile_4_3_chanxy_out[13];
    assign wire_7799 = lut_tile_4_3_chanxy_out[14];
    assign wire_7830 = lut_tile_4_3_chanxy_out[15];
    assign wire_7832 = lut_tile_4_3_chanxy_out[16];
    assign wire_7834 = lut_tile_4_3_chanxy_out[17];
    assign wire_7836 = lut_tile_4_3_chanxy_out[18];
    assign wire_7838 = lut_tile_4_3_chanxy_out[19];
    assign wire_7840 = lut_tile_4_3_chanxy_out[20];
    assign wire_7842 = lut_tile_4_3_chanxy_out[21];
    assign wire_7844 = lut_tile_4_3_chanxy_out[22];
    assign wire_7846 = lut_tile_4_3_chanxy_out[23];
    assign wire_7848 = lut_tile_4_3_chanxy_out[24];
    assign wire_7850 = lut_tile_4_3_chanxy_out[25];
    assign wire_7852 = lut_tile_4_3_chanxy_out[26];
    assign wire_7854 = lut_tile_4_3_chanxy_out[27];
    assign wire_7856 = lut_tile_4_3_chanxy_out[28];
    assign wire_7858 = lut_tile_4_3_chanxy_out[29];
    assign wire_11587 = lut_tile_4_3_chanxy_out[30];
    assign wire_11595 = lut_tile_4_3_chanxy_out[31];
    assign wire_11603 = lut_tile_4_3_chanxy_out[32];
    assign wire_11611 = lut_tile_4_3_chanxy_out[33];
    assign wire_11619 = lut_tile_4_3_chanxy_out[34];
    assign wire_11627 = lut_tile_4_3_chanxy_out[35];
    assign wire_11635 = lut_tile_4_3_chanxy_out[36];
    assign wire_11643 = lut_tile_4_3_chanxy_out[37];
    assign wire_11651 = lut_tile_4_3_chanxy_out[38];
    assign wire_11659 = lut_tile_4_3_chanxy_out[39];
    assign wire_11667 = lut_tile_4_3_chanxy_out[40];
    assign wire_11675 = lut_tile_4_3_chanxy_out[41];
    assign wire_11683 = lut_tile_4_3_chanxy_out[42];
    assign wire_11691 = lut_tile_4_3_chanxy_out[43];
    assign wire_11699 = lut_tile_4_3_chanxy_out[44];
    assign wire_11760 = lut_tile_4_3_chanxy_out[45];
    assign wire_11762 = lut_tile_4_3_chanxy_out[46];
    assign wire_11764 = lut_tile_4_3_chanxy_out[47];
    assign wire_11766 = lut_tile_4_3_chanxy_out[48];
    assign wire_11768 = lut_tile_4_3_chanxy_out[49];
    assign wire_11770 = lut_tile_4_3_chanxy_out[50];
    assign wire_11772 = lut_tile_4_3_chanxy_out[51];
    assign wire_11774 = lut_tile_4_3_chanxy_out[52];
    assign wire_11776 = lut_tile_4_3_chanxy_out[53];
    assign wire_11778 = lut_tile_4_3_chanxy_out[54];
    assign wire_11780 = lut_tile_4_3_chanxy_out[55];
    assign wire_11782 = lut_tile_4_3_chanxy_out[56];
    assign wire_11784 = lut_tile_4_3_chanxy_out[57];
    assign wire_11786 = lut_tile_4_3_chanxy_out[58];
    assign wire_11788 = lut_tile_4_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_4_chanxy_in = {wire_12088, wire_7501, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7304, wire_2751, wire_12080, wire_7529, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7312, wire_2751, wire_12072, wire_7527, wire_7439, wire_7438, wire_7429, wire_7428, wire_7419, wire_7418, wire_7320, wire_2751, wire_12064, wire_7525, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7328, wire_2241, wire_12056, wire_7523, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7336, wire_2241, wire_12048, wire_7521, wire_7437, wire_7436, wire_7427, wire_7426, wire_7417, wire_7416, wire_7344, wire_2241, wire_12040, wire_7519, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7352, wire_2755, wire_2241, wire_12032, wire_7517, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7360, wire_2755, wire_2241, wire_12024, wire_7515, wire_7435, wire_7434, wire_7425, wire_7424, wire_7415, wire_7414, wire_7368, wire_2755, wire_2241, wire_12016, wire_7513, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7376, wire_2755, wire_2237, wire_12008, wire_7511, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7384, wire_2755, wire_2237, wire_12000, wire_7509, wire_7433, wire_7432, wire_7423, wire_7422, wire_7413, wire_7412, wire_7392, wire_2755, wire_2237, wire_11992, wire_7507, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7400, wire_2751, wire_2237, wire_11984, wire_7505, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7408, wire_2751, wire_2237, wire_11976, wire_7503, wire_7431, wire_7430, wire_7421, wire_7420, wire_7411, wire_7410, wire_7296, wire_2751, wire_2237, wire_12209, wire_7919, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7680, wire_2751, wire_12207, wire_7891, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7792, wire_2751, wire_12205, wire_7893, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7784, wire_2751, wire_12203, wire_7895, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7776, wire_2241, wire_12201, wire_7897, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7768, wire_2241, wire_12199, wire_7899, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7760, wire_2241, wire_12197, wire_7901, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7752, wire_2755, wire_2241, wire_12195, wire_7903, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7744, wire_2755, wire_2241, wire_12193, wire_7905, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7736, wire_2755, wire_2241, wire_12191, wire_7907, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7728, wire_2755, wire_2237, wire_12189, wire_7909, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7720, wire_2755, wire_2237, wire_12187, wire_7911, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7712, wire_2755, wire_2237, wire_12185, wire_7913, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7704, wire_2751, wire_2237, wire_12183, wire_7915, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7696, wire_2751, wire_2237, wire_12181, wire_7917, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7688, wire_2751, wire_2237, wire_11817, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11698, wire_7798, wire_2280, wire_11815, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11586, wire_7790, wire_2280, wire_11813, wire_11729, wire_11728, wire_11719, wire_11718, wire_11709, wire_11708, wire_11594, wire_7782, wire_2280, wire_11811, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11602, wire_7774, wire_2240, wire_11809, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11610, wire_7766, wire_2240, wire_11807, wire_11727, wire_11726, wire_11717, wire_11716, wire_11707, wire_11706, wire_11618, wire_7758, wire_2240, wire_11805, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11626, wire_7750, wire_2284, wire_2240, wire_11803, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11634, wire_7742, wire_2284, wire_2240, wire_11801, wire_11725, wire_11724, wire_11715, wire_11714, wire_11705, wire_11704, wire_11642, wire_7734, wire_2284, wire_2240, wire_11799, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11650, wire_7726, wire_2284, wire_2236, wire_11797, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11658, wire_7718, wire_2284, wire_2236, wire_11795, wire_11723, wire_11722, wire_11713, wire_11712, wire_11703, wire_11702, wire_11666, wire_7710, wire_2284, wire_2236, wire_11793, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11674, wire_7702, wire_2280, wire_2236, wire_11791, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11682, wire_7694, wire_2280, wire_2236, wire_11819, wire_11721, wire_11720, wire_11711, wire_11710, wire_11701, wire_11700, wire_11690, wire_7686, wire_2280, wire_2236, wire_12183, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12074, wire_7919, wire_2280, wire_12185, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12066, wire_7917, wire_2280, wire_12187, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_12058, wire_7915, wire_2280, wire_12189, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12050, wire_7913, wire_2240, wire_12191, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12042, wire_7911, wire_2240, wire_12193, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12034, wire_7909, wire_2240, wire_12195, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12026, wire_7907, wire_2284, wire_2240, wire_12197, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12018, wire_7905, wire_2284, wire_2240, wire_12199, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12010, wire_7903, wire_2284, wire_2240, wire_12201, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12002, wire_7901, wire_2284, wire_2236, wire_12203, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_11994, wire_7899, wire_2284, wire_2236, wire_12205, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_11986, wire_7897, wire_2284, wire_2236, wire_12207, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_11978, wire_7895, wire_2280, wire_2236, wire_12209, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_11970, wire_7893, wire_2280, wire_2236, wire_12181, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12082, wire_7891, wire_2280, wire_2236};
    // CHNAXY TOTAL: 636
    assign wire_7681 = lut_tile_4_4_chanxy_out[0];
    assign wire_7689 = lut_tile_4_4_chanxy_out[1];
    assign wire_7697 = lut_tile_4_4_chanxy_out[2];
    assign wire_7705 = lut_tile_4_4_chanxy_out[3];
    assign wire_7713 = lut_tile_4_4_chanxy_out[4];
    assign wire_7721 = lut_tile_4_4_chanxy_out[5];
    assign wire_7729 = lut_tile_4_4_chanxy_out[6];
    assign wire_7737 = lut_tile_4_4_chanxy_out[7];
    assign wire_7745 = lut_tile_4_4_chanxy_out[8];
    assign wire_7753 = lut_tile_4_4_chanxy_out[9];
    assign wire_7761 = lut_tile_4_4_chanxy_out[10];
    assign wire_7769 = lut_tile_4_4_chanxy_out[11];
    assign wire_7777 = lut_tile_4_4_chanxy_out[12];
    assign wire_7785 = lut_tile_4_4_chanxy_out[13];
    assign wire_7793 = lut_tile_4_4_chanxy_out[14];
    assign wire_7860 = lut_tile_4_4_chanxy_out[15];
    assign wire_7862 = lut_tile_4_4_chanxy_out[16];
    assign wire_7864 = lut_tile_4_4_chanxy_out[17];
    assign wire_7866 = lut_tile_4_4_chanxy_out[18];
    assign wire_7868 = lut_tile_4_4_chanxy_out[19];
    assign wire_7870 = lut_tile_4_4_chanxy_out[20];
    assign wire_7872 = lut_tile_4_4_chanxy_out[21];
    assign wire_7874 = lut_tile_4_4_chanxy_out[22];
    assign wire_7876 = lut_tile_4_4_chanxy_out[23];
    assign wire_7878 = lut_tile_4_4_chanxy_out[24];
    assign wire_7880 = lut_tile_4_4_chanxy_out[25];
    assign wire_7882 = lut_tile_4_4_chanxy_out[26];
    assign wire_7884 = lut_tile_4_4_chanxy_out[27];
    assign wire_7886 = lut_tile_4_4_chanxy_out[28];
    assign wire_7888 = lut_tile_4_4_chanxy_out[29];
    assign wire_11971 = lut_tile_4_4_chanxy_out[30];
    assign wire_11979 = lut_tile_4_4_chanxy_out[31];
    assign wire_11987 = lut_tile_4_4_chanxy_out[32];
    assign wire_11995 = lut_tile_4_4_chanxy_out[33];
    assign wire_12003 = lut_tile_4_4_chanxy_out[34];
    assign wire_12011 = lut_tile_4_4_chanxy_out[35];
    assign wire_12019 = lut_tile_4_4_chanxy_out[36];
    assign wire_12027 = lut_tile_4_4_chanxy_out[37];
    assign wire_12035 = lut_tile_4_4_chanxy_out[38];
    assign wire_12043 = lut_tile_4_4_chanxy_out[39];
    assign wire_12051 = lut_tile_4_4_chanxy_out[40];
    assign wire_12059 = lut_tile_4_4_chanxy_out[41];
    assign wire_12067 = lut_tile_4_4_chanxy_out[42];
    assign wire_12075 = lut_tile_4_4_chanxy_out[43];
    assign wire_12083 = lut_tile_4_4_chanxy_out[44];
    assign wire_12150 = lut_tile_4_4_chanxy_out[45];
    assign wire_12152 = lut_tile_4_4_chanxy_out[46];
    assign wire_12154 = lut_tile_4_4_chanxy_out[47];
    assign wire_12156 = lut_tile_4_4_chanxy_out[48];
    assign wire_12158 = lut_tile_4_4_chanxy_out[49];
    assign wire_12160 = lut_tile_4_4_chanxy_out[50];
    assign wire_12162 = lut_tile_4_4_chanxy_out[51];
    assign wire_12164 = lut_tile_4_4_chanxy_out[52];
    assign wire_12166 = lut_tile_4_4_chanxy_out[53];
    assign wire_12168 = lut_tile_4_4_chanxy_out[54];
    assign wire_12170 = lut_tile_4_4_chanxy_out[55];
    assign wire_12172 = lut_tile_4_4_chanxy_out[56];
    assign wire_12174 = lut_tile_4_4_chanxy_out[57];
    assign wire_12176 = lut_tile_4_4_chanxy_out[58];
    assign wire_12178 = lut_tile_4_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_5_chanxy_in = {wire_12472, wire_7531, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7412, wire_3267, wire_12464, wire_7559, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7414, wire_3267, wire_12456, wire_7557, wire_7469, wire_7468, wire_7459, wire_7458, wire_7449, wire_7448, wire_7416, wire_3267, wire_12448, wire_7555, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7418, wire_2757, wire_12440, wire_7553, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7420, wire_2757, wire_12432, wire_7551, wire_7467, wire_7466, wire_7457, wire_7456, wire_7447, wire_7446, wire_7422, wire_2757, wire_12424, wire_7549, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7424, wire_3271, wire_2757, wire_12416, wire_7547, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7426, wire_3271, wire_2757, wire_12408, wire_7545, wire_7465, wire_7464, wire_7455, wire_7454, wire_7445, wire_7444, wire_7428, wire_3271, wire_2757, wire_12400, wire_7543, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7430, wire_3271, wire_2753, wire_12392, wire_7541, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7432, wire_3271, wire_2753, wire_12384, wire_7539, wire_7463, wire_7462, wire_7453, wire_7452, wire_7443, wire_7442, wire_7434, wire_3271, wire_2753, wire_12376, wire_7537, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7436, wire_3267, wire_2753, wire_12368, wire_7535, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7438, wire_3267, wire_2753, wire_12360, wire_7533, wire_7461, wire_7460, wire_7451, wire_7450, wire_7441, wire_7440, wire_7410, wire_3267, wire_2753, wire_12599, wire_7949, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7800, wire_3267, wire_12597, wire_7921, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7828, wire_3267, wire_12595, wire_7923, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7826, wire_3267, wire_12593, wire_7925, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7824, wire_2757, wire_12591, wire_7927, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7822, wire_2757, wire_12589, wire_7929, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7820, wire_2757, wire_12587, wire_7931, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7818, wire_3271, wire_2757, wire_12585, wire_7933, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7816, wire_3271, wire_2757, wire_12583, wire_7935, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7814, wire_3271, wire_2757, wire_12581, wire_7937, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7812, wire_3271, wire_2753, wire_12579, wire_7939, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7810, wire_3271, wire_2753, wire_12577, wire_7941, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7808, wire_3271, wire_2753, wire_12575, wire_7943, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7806, wire_3267, wire_2753, wire_12573, wire_7945, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7804, wire_3267, wire_2753, wire_12571, wire_7947, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7802, wire_3267, wire_2753, wire_12207, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12082, wire_7792, wire_2796, wire_12205, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_11970, wire_7784, wire_2796, wire_12203, wire_12119, wire_12118, wire_12109, wire_12108, wire_12099, wire_12098, wire_11978, wire_7776, wire_2796, wire_12201, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_11986, wire_7768, wire_2756, wire_12199, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_11994, wire_7760, wire_2756, wire_12197, wire_12117, wire_12116, wire_12107, wire_12106, wire_12097, wire_12096, wire_12002, wire_7752, wire_2756, wire_12195, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12010, wire_7744, wire_2800, wire_2756, wire_12193, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12018, wire_7736, wire_2800, wire_2756, wire_12191, wire_12115, wire_12114, wire_12105, wire_12104, wire_12095, wire_12094, wire_12026, wire_7728, wire_2800, wire_2756, wire_12189, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12034, wire_7720, wire_2800, wire_2752, wire_12187, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12042, wire_7712, wire_2800, wire_2752, wire_12185, wire_12113, wire_12112, wire_12103, wire_12102, wire_12093, wire_12092, wire_12050, wire_7704, wire_2800, wire_2752, wire_12183, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12058, wire_7696, wire_2796, wire_2752, wire_12181, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12066, wire_7688, wire_2796, wire_2752, wire_12209, wire_12111, wire_12110, wire_12101, wire_12100, wire_12091, wire_12090, wire_12074, wire_7680, wire_2796, wire_2752, wire_12573, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12466, wire_7949, wire_2796, wire_12575, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12458, wire_7947, wire_2796, wire_12577, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12450, wire_7945, wire_2796, wire_12579, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12442, wire_7943, wire_2756, wire_12581, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12434, wire_7941, wire_2756, wire_12583, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12426, wire_7939, wire_2756, wire_12585, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12418, wire_7937, wire_2800, wire_2756, wire_12587, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12410, wire_7935, wire_2800, wire_2756, wire_12589, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12402, wire_7933, wire_2800, wire_2756, wire_12591, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12394, wire_7931, wire_2800, wire_2752, wire_12593, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12386, wire_7929, wire_2800, wire_2752, wire_12595, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12378, wire_7927, wire_2800, wire_2752, wire_12597, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12370, wire_7925, wire_2796, wire_2752, wire_12599, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12362, wire_7923, wire_2796, wire_2752, wire_12571, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12474, wire_7921, wire_2796, wire_2752};
    // CHNAXY TOTAL: 636
    assign wire_7801 = lut_tile_4_5_chanxy_out[0];
    assign wire_7803 = lut_tile_4_5_chanxy_out[1];
    assign wire_7805 = lut_tile_4_5_chanxy_out[2];
    assign wire_7807 = lut_tile_4_5_chanxy_out[3];
    assign wire_7809 = lut_tile_4_5_chanxy_out[4];
    assign wire_7811 = lut_tile_4_5_chanxy_out[5];
    assign wire_7813 = lut_tile_4_5_chanxy_out[6];
    assign wire_7815 = lut_tile_4_5_chanxy_out[7];
    assign wire_7817 = lut_tile_4_5_chanxy_out[8];
    assign wire_7819 = lut_tile_4_5_chanxy_out[9];
    assign wire_7821 = lut_tile_4_5_chanxy_out[10];
    assign wire_7823 = lut_tile_4_5_chanxy_out[11];
    assign wire_7825 = lut_tile_4_5_chanxy_out[12];
    assign wire_7827 = lut_tile_4_5_chanxy_out[13];
    assign wire_7829 = lut_tile_4_5_chanxy_out[14];
    assign wire_7890 = lut_tile_4_5_chanxy_out[15];
    assign wire_7892 = lut_tile_4_5_chanxy_out[16];
    assign wire_7894 = lut_tile_4_5_chanxy_out[17];
    assign wire_7896 = lut_tile_4_5_chanxy_out[18];
    assign wire_7898 = lut_tile_4_5_chanxy_out[19];
    assign wire_7900 = lut_tile_4_5_chanxy_out[20];
    assign wire_7902 = lut_tile_4_5_chanxy_out[21];
    assign wire_7904 = lut_tile_4_5_chanxy_out[22];
    assign wire_7906 = lut_tile_4_5_chanxy_out[23];
    assign wire_7908 = lut_tile_4_5_chanxy_out[24];
    assign wire_7910 = lut_tile_4_5_chanxy_out[25];
    assign wire_7912 = lut_tile_4_5_chanxy_out[26];
    assign wire_7914 = lut_tile_4_5_chanxy_out[27];
    assign wire_7916 = lut_tile_4_5_chanxy_out[28];
    assign wire_7918 = lut_tile_4_5_chanxy_out[29];
    assign wire_12363 = lut_tile_4_5_chanxy_out[30];
    assign wire_12371 = lut_tile_4_5_chanxy_out[31];
    assign wire_12379 = lut_tile_4_5_chanxy_out[32];
    assign wire_12387 = lut_tile_4_5_chanxy_out[33];
    assign wire_12395 = lut_tile_4_5_chanxy_out[34];
    assign wire_12403 = lut_tile_4_5_chanxy_out[35];
    assign wire_12411 = lut_tile_4_5_chanxy_out[36];
    assign wire_12419 = lut_tile_4_5_chanxy_out[37];
    assign wire_12427 = lut_tile_4_5_chanxy_out[38];
    assign wire_12435 = lut_tile_4_5_chanxy_out[39];
    assign wire_12443 = lut_tile_4_5_chanxy_out[40];
    assign wire_12451 = lut_tile_4_5_chanxy_out[41];
    assign wire_12459 = lut_tile_4_5_chanxy_out[42];
    assign wire_12467 = lut_tile_4_5_chanxy_out[43];
    assign wire_12475 = lut_tile_4_5_chanxy_out[44];
    assign wire_12540 = lut_tile_4_5_chanxy_out[45];
    assign wire_12542 = lut_tile_4_5_chanxy_out[46];
    assign wire_12544 = lut_tile_4_5_chanxy_out[47];
    assign wire_12546 = lut_tile_4_5_chanxy_out[48];
    assign wire_12548 = lut_tile_4_5_chanxy_out[49];
    assign wire_12550 = lut_tile_4_5_chanxy_out[50];
    assign wire_12552 = lut_tile_4_5_chanxy_out[51];
    assign wire_12554 = lut_tile_4_5_chanxy_out[52];
    assign wire_12556 = lut_tile_4_5_chanxy_out[53];
    assign wire_12558 = lut_tile_4_5_chanxy_out[54];
    assign wire_12560 = lut_tile_4_5_chanxy_out[55];
    assign wire_12562 = lut_tile_4_5_chanxy_out[56];
    assign wire_12564 = lut_tile_4_5_chanxy_out[57];
    assign wire_12566 = lut_tile_4_5_chanxy_out[58];
    assign wire_12568 = lut_tile_4_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_6_chanxy_in = {wire_12864, wire_7561, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7442, wire_3783, wire_12856, wire_7589, wire_7499, wire_7498, wire_7489, wire_7488, wire_7479, wire_7478, wire_7444, wire_3783, wire_12848, wire_7587, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7446, wire_3783, wire_12840, wire_7585, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7448, wire_3273, wire_12832, wire_7583, wire_7497, wire_7496, wire_7487, wire_7486, wire_7477, wire_7476, wire_7450, wire_3273, wire_12824, wire_7581, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7452, wire_3273, wire_12816, wire_7579, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7454, wire_3787, wire_3273, wire_12808, wire_7577, wire_7495, wire_7494, wire_7485, wire_7484, wire_7475, wire_7474, wire_7456, wire_3787, wire_3273, wire_12800, wire_7575, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7458, wire_3787, wire_3273, wire_12792, wire_7573, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7460, wire_3787, wire_3269, wire_12784, wire_7571, wire_7493, wire_7492, wire_7483, wire_7482, wire_7473, wire_7472, wire_7462, wire_3787, wire_3269, wire_12776, wire_7569, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7464, wire_3787, wire_3269, wire_12768, wire_7567, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7466, wire_3783, wire_3269, wire_12760, wire_7565, wire_7491, wire_7490, wire_7481, wire_7480, wire_7471, wire_7470, wire_7468, wire_3783, wire_3269, wire_12752, wire_7563, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7440, wire_3783, wire_3269, wire_12989, wire_7979, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7830, wire_3783, wire_12987, wire_7951, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7858, wire_3783, wire_12985, wire_7953, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7856, wire_3783, wire_12983, wire_7955, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7854, wire_3273, wire_12981, wire_7957, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7852, wire_3273, wire_12979, wire_7959, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7850, wire_3273, wire_12977, wire_7961, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7848, wire_3787, wire_3273, wire_12975, wire_7963, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7846, wire_3787, wire_3273, wire_12973, wire_7965, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7844, wire_3787, wire_3273, wire_12971, wire_7967, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7842, wire_3787, wire_3269, wire_12969, wire_7969, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7840, wire_3787, wire_3269, wire_12967, wire_7971, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7838, wire_3787, wire_3269, wire_12965, wire_7973, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7836, wire_3783, wire_3269, wire_12963, wire_7975, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7834, wire_3783, wire_3269, wire_12961, wire_7977, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7832, wire_3783, wire_3269, wire_12597, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12474, wire_7828, wire_3312, wire_12595, wire_12509, wire_12508, wire_12499, wire_12498, wire_12489, wire_12488, wire_12362, wire_7826, wire_3312, wire_12593, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12370, wire_7824, wire_3312, wire_12591, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12378, wire_7822, wire_3272, wire_12589, wire_12507, wire_12506, wire_12497, wire_12496, wire_12487, wire_12486, wire_12386, wire_7820, wire_3272, wire_12587, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12394, wire_7818, wire_3272, wire_12585, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12402, wire_7816, wire_3316, wire_3272, wire_12583, wire_12505, wire_12504, wire_12495, wire_12494, wire_12485, wire_12484, wire_12410, wire_7814, wire_3316, wire_3272, wire_12581, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12418, wire_7812, wire_3316, wire_3272, wire_12579, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12426, wire_7810, wire_3316, wire_3268, wire_12577, wire_12503, wire_12502, wire_12493, wire_12492, wire_12483, wire_12482, wire_12434, wire_7808, wire_3316, wire_3268, wire_12575, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12442, wire_7806, wire_3316, wire_3268, wire_12573, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12450, wire_7804, wire_3312, wire_3268, wire_12571, wire_12501, wire_12500, wire_12491, wire_12490, wire_12481, wire_12480, wire_12458, wire_7802, wire_3312, wire_3268, wire_12599, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12466, wire_7800, wire_3312, wire_3268, wire_12963, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12858, wire_7979, wire_3312, wire_12965, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12850, wire_7977, wire_3312, wire_12967, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12842, wire_7975, wire_3312, wire_12969, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12834, wire_7973, wire_3272, wire_12971, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12826, wire_7971, wire_3272, wire_12973, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12818, wire_7969, wire_3272, wire_12975, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12810, wire_7967, wire_3316, wire_3272, wire_12977, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12802, wire_7965, wire_3316, wire_3272, wire_12979, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12794, wire_7963, wire_3316, wire_3272, wire_12981, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12786, wire_7961, wire_3316, wire_3268, wire_12983, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12778, wire_7959, wire_3316, wire_3268, wire_12985, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12770, wire_7957, wire_3316, wire_3268, wire_12987, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12762, wire_7955, wire_3312, wire_3268, wire_12989, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12754, wire_7953, wire_3312, wire_3268, wire_12961, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12866, wire_7951, wire_3312, wire_3268};
    // CHNAXY TOTAL: 636
    assign wire_7831 = lut_tile_4_6_chanxy_out[0];
    assign wire_7833 = lut_tile_4_6_chanxy_out[1];
    assign wire_7835 = lut_tile_4_6_chanxy_out[2];
    assign wire_7837 = lut_tile_4_6_chanxy_out[3];
    assign wire_7839 = lut_tile_4_6_chanxy_out[4];
    assign wire_7841 = lut_tile_4_6_chanxy_out[5];
    assign wire_7843 = lut_tile_4_6_chanxy_out[6];
    assign wire_7845 = lut_tile_4_6_chanxy_out[7];
    assign wire_7847 = lut_tile_4_6_chanxy_out[8];
    assign wire_7849 = lut_tile_4_6_chanxy_out[9];
    assign wire_7851 = lut_tile_4_6_chanxy_out[10];
    assign wire_7853 = lut_tile_4_6_chanxy_out[11];
    assign wire_7855 = lut_tile_4_6_chanxy_out[12];
    assign wire_7857 = lut_tile_4_6_chanxy_out[13];
    assign wire_7859 = lut_tile_4_6_chanxy_out[14];
    assign wire_7920 = lut_tile_4_6_chanxy_out[15];
    assign wire_7922 = lut_tile_4_6_chanxy_out[16];
    assign wire_7924 = lut_tile_4_6_chanxy_out[17];
    assign wire_7926 = lut_tile_4_6_chanxy_out[18];
    assign wire_7928 = lut_tile_4_6_chanxy_out[19];
    assign wire_7930 = lut_tile_4_6_chanxy_out[20];
    assign wire_7932 = lut_tile_4_6_chanxy_out[21];
    assign wire_7934 = lut_tile_4_6_chanxy_out[22];
    assign wire_7936 = lut_tile_4_6_chanxy_out[23];
    assign wire_7938 = lut_tile_4_6_chanxy_out[24];
    assign wire_7940 = lut_tile_4_6_chanxy_out[25];
    assign wire_7942 = lut_tile_4_6_chanxy_out[26];
    assign wire_7944 = lut_tile_4_6_chanxy_out[27];
    assign wire_7946 = lut_tile_4_6_chanxy_out[28];
    assign wire_7948 = lut_tile_4_6_chanxy_out[29];
    assign wire_12755 = lut_tile_4_6_chanxy_out[30];
    assign wire_12763 = lut_tile_4_6_chanxy_out[31];
    assign wire_12771 = lut_tile_4_6_chanxy_out[32];
    assign wire_12779 = lut_tile_4_6_chanxy_out[33];
    assign wire_12787 = lut_tile_4_6_chanxy_out[34];
    assign wire_12795 = lut_tile_4_6_chanxy_out[35];
    assign wire_12803 = lut_tile_4_6_chanxy_out[36];
    assign wire_12811 = lut_tile_4_6_chanxy_out[37];
    assign wire_12819 = lut_tile_4_6_chanxy_out[38];
    assign wire_12827 = lut_tile_4_6_chanxy_out[39];
    assign wire_12835 = lut_tile_4_6_chanxy_out[40];
    assign wire_12843 = lut_tile_4_6_chanxy_out[41];
    assign wire_12851 = lut_tile_4_6_chanxy_out[42];
    assign wire_12859 = lut_tile_4_6_chanxy_out[43];
    assign wire_12867 = lut_tile_4_6_chanxy_out[44];
    assign wire_12930 = lut_tile_4_6_chanxy_out[45];
    assign wire_12932 = lut_tile_4_6_chanxy_out[46];
    assign wire_12934 = lut_tile_4_6_chanxy_out[47];
    assign wire_12936 = lut_tile_4_6_chanxy_out[48];
    assign wire_12938 = lut_tile_4_6_chanxy_out[49];
    assign wire_12940 = lut_tile_4_6_chanxy_out[50];
    assign wire_12942 = lut_tile_4_6_chanxy_out[51];
    assign wire_12944 = lut_tile_4_6_chanxy_out[52];
    assign wire_12946 = lut_tile_4_6_chanxy_out[53];
    assign wire_12948 = lut_tile_4_6_chanxy_out[54];
    assign wire_12950 = lut_tile_4_6_chanxy_out[55];
    assign wire_12952 = lut_tile_4_6_chanxy_out[56];
    assign wire_12954 = lut_tile_4_6_chanxy_out[57];
    assign wire_12956 = lut_tile_4_6_chanxy_out[58];
    assign wire_12958 = lut_tile_4_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_7_chanxy_in = {wire_13256, wire_7591, wire_7529, wire_7528, wire_7519, wire_7518, wire_7509, wire_7508, wire_7472, wire_4299, wire_13248, wire_7619, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7474, wire_4299, wire_13240, wire_7617, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7476, wire_4299, wire_13232, wire_7615, wire_7527, wire_7526, wire_7517, wire_7516, wire_7507, wire_7506, wire_7478, wire_3789, wire_13224, wire_7613, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7480, wire_3789, wire_13216, wire_7611, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7482, wire_3789, wire_13208, wire_7609, wire_7525, wire_7524, wire_7515, wire_7514, wire_7505, wire_7504, wire_7484, wire_4303, wire_3789, wire_13200, wire_7607, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7486, wire_4303, wire_3789, wire_13192, wire_7605, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7488, wire_4303, wire_3789, wire_13184, wire_7603, wire_7523, wire_7522, wire_7513, wire_7512, wire_7503, wire_7502, wire_7490, wire_4303, wire_3785, wire_13176, wire_7601, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7492, wire_4303, wire_3785, wire_13168, wire_7599, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7494, wire_4303, wire_3785, wire_13160, wire_7597, wire_7521, wire_7520, wire_7511, wire_7510, wire_7501, wire_7500, wire_7496, wire_4299, wire_3785, wire_13152, wire_7595, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7498, wire_4299, wire_3785, wire_13144, wire_7593, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7470, wire_4299, wire_3785, wire_13379, wire_8009, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7860, wire_4299, wire_13377, wire_7981, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7888, wire_4299, wire_13375, wire_7983, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7886, wire_4299, wire_13373, wire_7985, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7884, wire_3789, wire_13371, wire_7987, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7882, wire_3789, wire_13369, wire_7989, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7880, wire_3789, wire_13367, wire_7991, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7878, wire_4303, wire_3789, wire_13365, wire_7993, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7876, wire_4303, wire_3789, wire_13363, wire_7995, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7874, wire_4303, wire_3789, wire_13361, wire_7997, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7872, wire_4303, wire_3785, wire_13359, wire_7999, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7870, wire_4303, wire_3785, wire_13357, wire_8001, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7868, wire_4303, wire_3785, wire_13355, wire_8003, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7866, wire_4299, wire_3785, wire_13353, wire_8005, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7864, wire_4299, wire_3785, wire_13351, wire_8007, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7862, wire_4299, wire_3785, wire_12987, wire_12899, wire_12898, wire_12889, wire_12888, wire_12879, wire_12878, wire_12866, wire_7858, wire_3828, wire_12985, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12754, wire_7856, wire_3828, wire_12983, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12762, wire_7854, wire_3828, wire_12981, wire_12897, wire_12896, wire_12887, wire_12886, wire_12877, wire_12876, wire_12770, wire_7852, wire_3788, wire_12979, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12778, wire_7850, wire_3788, wire_12977, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12786, wire_7848, wire_3788, wire_12975, wire_12895, wire_12894, wire_12885, wire_12884, wire_12875, wire_12874, wire_12794, wire_7846, wire_3832, wire_3788, wire_12973, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12802, wire_7844, wire_3832, wire_3788, wire_12971, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12810, wire_7842, wire_3832, wire_3788, wire_12969, wire_12893, wire_12892, wire_12883, wire_12882, wire_12873, wire_12872, wire_12818, wire_7840, wire_3832, wire_3784, wire_12967, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12826, wire_7838, wire_3832, wire_3784, wire_12965, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12834, wire_7836, wire_3832, wire_3784, wire_12963, wire_12891, wire_12890, wire_12881, wire_12880, wire_12871, wire_12870, wire_12842, wire_7834, wire_3828, wire_3784, wire_12961, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12850, wire_7832, wire_3828, wire_3784, wire_12989, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12858, wire_7830, wire_3828, wire_3784, wire_13353, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13250, wire_8009, wire_3828, wire_13355, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13242, wire_8007, wire_3828, wire_13357, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13234, wire_8005, wire_3828, wire_13359, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13226, wire_8003, wire_3788, wire_13361, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13218, wire_8001, wire_3788, wire_13363, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13210, wire_7999, wire_3788, wire_13365, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13202, wire_7997, wire_3832, wire_3788, wire_13367, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13194, wire_7995, wire_3832, wire_3788, wire_13369, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13186, wire_7993, wire_3832, wire_3788, wire_13371, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13178, wire_7991, wire_3832, wire_3784, wire_13373, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13170, wire_7989, wire_3832, wire_3784, wire_13375, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13162, wire_7987, wire_3832, wire_3784, wire_13377, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13154, wire_7985, wire_3828, wire_3784, wire_13379, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13146, wire_7983, wire_3828, wire_3784, wire_13351, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13258, wire_7981, wire_3828, wire_3784};
    // CHNAXY TOTAL: 636
    assign wire_7861 = lut_tile_4_7_chanxy_out[0];
    assign wire_7863 = lut_tile_4_7_chanxy_out[1];
    assign wire_7865 = lut_tile_4_7_chanxy_out[2];
    assign wire_7867 = lut_tile_4_7_chanxy_out[3];
    assign wire_7869 = lut_tile_4_7_chanxy_out[4];
    assign wire_7871 = lut_tile_4_7_chanxy_out[5];
    assign wire_7873 = lut_tile_4_7_chanxy_out[6];
    assign wire_7875 = lut_tile_4_7_chanxy_out[7];
    assign wire_7877 = lut_tile_4_7_chanxy_out[8];
    assign wire_7879 = lut_tile_4_7_chanxy_out[9];
    assign wire_7881 = lut_tile_4_7_chanxy_out[10];
    assign wire_7883 = lut_tile_4_7_chanxy_out[11];
    assign wire_7885 = lut_tile_4_7_chanxy_out[12];
    assign wire_7887 = lut_tile_4_7_chanxy_out[13];
    assign wire_7889 = lut_tile_4_7_chanxy_out[14];
    assign wire_7950 = lut_tile_4_7_chanxy_out[15];
    assign wire_7952 = lut_tile_4_7_chanxy_out[16];
    assign wire_7954 = lut_tile_4_7_chanxy_out[17];
    assign wire_7956 = lut_tile_4_7_chanxy_out[18];
    assign wire_7958 = lut_tile_4_7_chanxy_out[19];
    assign wire_7960 = lut_tile_4_7_chanxy_out[20];
    assign wire_7962 = lut_tile_4_7_chanxy_out[21];
    assign wire_7964 = lut_tile_4_7_chanxy_out[22];
    assign wire_7966 = lut_tile_4_7_chanxy_out[23];
    assign wire_7968 = lut_tile_4_7_chanxy_out[24];
    assign wire_7970 = lut_tile_4_7_chanxy_out[25];
    assign wire_7972 = lut_tile_4_7_chanxy_out[26];
    assign wire_7974 = lut_tile_4_7_chanxy_out[27];
    assign wire_7976 = lut_tile_4_7_chanxy_out[28];
    assign wire_7978 = lut_tile_4_7_chanxy_out[29];
    assign wire_13147 = lut_tile_4_7_chanxy_out[30];
    assign wire_13155 = lut_tile_4_7_chanxy_out[31];
    assign wire_13163 = lut_tile_4_7_chanxy_out[32];
    assign wire_13171 = lut_tile_4_7_chanxy_out[33];
    assign wire_13179 = lut_tile_4_7_chanxy_out[34];
    assign wire_13187 = lut_tile_4_7_chanxy_out[35];
    assign wire_13195 = lut_tile_4_7_chanxy_out[36];
    assign wire_13203 = lut_tile_4_7_chanxy_out[37];
    assign wire_13211 = lut_tile_4_7_chanxy_out[38];
    assign wire_13219 = lut_tile_4_7_chanxy_out[39];
    assign wire_13227 = lut_tile_4_7_chanxy_out[40];
    assign wire_13235 = lut_tile_4_7_chanxy_out[41];
    assign wire_13243 = lut_tile_4_7_chanxy_out[42];
    assign wire_13251 = lut_tile_4_7_chanxy_out[43];
    assign wire_13259 = lut_tile_4_7_chanxy_out[44];
    assign wire_13320 = lut_tile_4_7_chanxy_out[45];
    assign wire_13322 = lut_tile_4_7_chanxy_out[46];
    assign wire_13324 = lut_tile_4_7_chanxy_out[47];
    assign wire_13326 = lut_tile_4_7_chanxy_out[48];
    assign wire_13328 = lut_tile_4_7_chanxy_out[49];
    assign wire_13330 = lut_tile_4_7_chanxy_out[50];
    assign wire_13332 = lut_tile_4_7_chanxy_out[51];
    assign wire_13334 = lut_tile_4_7_chanxy_out[52];
    assign wire_13336 = lut_tile_4_7_chanxy_out[53];
    assign wire_13338 = lut_tile_4_7_chanxy_out[54];
    assign wire_13340 = lut_tile_4_7_chanxy_out[55];
    assign wire_13342 = lut_tile_4_7_chanxy_out[56];
    assign wire_13344 = lut_tile_4_7_chanxy_out[57];
    assign wire_13346 = lut_tile_4_7_chanxy_out[58];
    assign wire_13348 = lut_tile_4_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_8_chanxy_in = {wire_13648, wire_7621, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7502, wire_4815, wire_13640, wire_7649, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7504, wire_4815, wire_13632, wire_7647, wire_7559, wire_7558, wire_7549, wire_7548, wire_7539, wire_7538, wire_7506, wire_4815, wire_13624, wire_7645, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7508, wire_4305, wire_13616, wire_7643, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7510, wire_4305, wire_13608, wire_7641, wire_7557, wire_7556, wire_7547, wire_7546, wire_7537, wire_7536, wire_7512, wire_4305, wire_13600, wire_7639, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7514, wire_4819, wire_4305, wire_13592, wire_7637, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7516, wire_4819, wire_4305, wire_13584, wire_7635, wire_7555, wire_7554, wire_7545, wire_7544, wire_7535, wire_7534, wire_7518, wire_4819, wire_4305, wire_13576, wire_7633, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7520, wire_4819, wire_4301, wire_13568, wire_7631, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7522, wire_4819, wire_4301, wire_13560, wire_7629, wire_7553, wire_7552, wire_7543, wire_7542, wire_7533, wire_7532, wire_7524, wire_4819, wire_4301, wire_13552, wire_7627, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7526, wire_4815, wire_4301, wire_13544, wire_7625, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7528, wire_4815, wire_4301, wire_13536, wire_7623, wire_7551, wire_7550, wire_7541, wire_7540, wire_7531, wire_7530, wire_7500, wire_4815, wire_4301, wire_13769, wire_8039, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7890, wire_4815, wire_13767, wire_8011, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7918, wire_4815, wire_13765, wire_8013, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7916, wire_4815, wire_13763, wire_8015, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7914, wire_4305, wire_13761, wire_8017, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7912, wire_4305, wire_13759, wire_8019, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7910, wire_4305, wire_13757, wire_8021, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7908, wire_4819, wire_4305, wire_13755, wire_8023, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7906, wire_4819, wire_4305, wire_13753, wire_8025, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7904, wire_4819, wire_4305, wire_13751, wire_8027, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7902, wire_4819, wire_4301, wire_13749, wire_8029, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7900, wire_4819, wire_4301, wire_13747, wire_8031, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7898, wire_4819, wire_4301, wire_13745, wire_8033, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7896, wire_4815, wire_4301, wire_13743, wire_8035, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7894, wire_4815, wire_4301, wire_13741, wire_8037, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7892, wire_4815, wire_4301, wire_13377, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13258, wire_7888, wire_4344, wire_13375, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13146, wire_7886, wire_4344, wire_13373, wire_13289, wire_13288, wire_13279, wire_13278, wire_13269, wire_13268, wire_13154, wire_7884, wire_4344, wire_13371, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13162, wire_7882, wire_4304, wire_13369, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13170, wire_7880, wire_4304, wire_13367, wire_13287, wire_13286, wire_13277, wire_13276, wire_13267, wire_13266, wire_13178, wire_7878, wire_4304, wire_13365, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13186, wire_7876, wire_4348, wire_4304, wire_13363, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13194, wire_7874, wire_4348, wire_4304, wire_13361, wire_13285, wire_13284, wire_13275, wire_13274, wire_13265, wire_13264, wire_13202, wire_7872, wire_4348, wire_4304, wire_13359, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13210, wire_7870, wire_4348, wire_4300, wire_13357, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13218, wire_7868, wire_4348, wire_4300, wire_13355, wire_13283, wire_13282, wire_13273, wire_13272, wire_13263, wire_13262, wire_13226, wire_7866, wire_4348, wire_4300, wire_13353, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13234, wire_7864, wire_4344, wire_4300, wire_13351, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13242, wire_7862, wire_4344, wire_4300, wire_13379, wire_13281, wire_13280, wire_13271, wire_13270, wire_13261, wire_13260, wire_13250, wire_7860, wire_4344, wire_4300, wire_13743, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13634, wire_8039, wire_4344, wire_13745, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13626, wire_8037, wire_4344, wire_13747, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13618, wire_8035, wire_4344, wire_13749, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13610, wire_8033, wire_4304, wire_13751, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13602, wire_8031, wire_4304, wire_13753, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13594, wire_8029, wire_4304, wire_13755, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13586, wire_8027, wire_4348, wire_4304, wire_13757, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13578, wire_8025, wire_4348, wire_4304, wire_13759, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13570, wire_8023, wire_4348, wire_4304, wire_13761, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13562, wire_8021, wire_4348, wire_4300, wire_13763, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13554, wire_8019, wire_4348, wire_4300, wire_13765, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13546, wire_8017, wire_4348, wire_4300, wire_13767, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13538, wire_8015, wire_4344, wire_4300, wire_13769, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13530, wire_8013, wire_4344, wire_4300, wire_13741, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13642, wire_8011, wire_4344, wire_4300};
    // CHNAXY TOTAL: 636
    assign wire_7891 = lut_tile_4_8_chanxy_out[0];
    assign wire_7893 = lut_tile_4_8_chanxy_out[1];
    assign wire_7895 = lut_tile_4_8_chanxy_out[2];
    assign wire_7897 = lut_tile_4_8_chanxy_out[3];
    assign wire_7899 = lut_tile_4_8_chanxy_out[4];
    assign wire_7901 = lut_tile_4_8_chanxy_out[5];
    assign wire_7903 = lut_tile_4_8_chanxy_out[6];
    assign wire_7905 = lut_tile_4_8_chanxy_out[7];
    assign wire_7907 = lut_tile_4_8_chanxy_out[8];
    assign wire_7909 = lut_tile_4_8_chanxy_out[9];
    assign wire_7911 = lut_tile_4_8_chanxy_out[10];
    assign wire_7913 = lut_tile_4_8_chanxy_out[11];
    assign wire_7915 = lut_tile_4_8_chanxy_out[12];
    assign wire_7917 = lut_tile_4_8_chanxy_out[13];
    assign wire_7919 = lut_tile_4_8_chanxy_out[14];
    assign wire_7980 = lut_tile_4_8_chanxy_out[15];
    assign wire_7982 = lut_tile_4_8_chanxy_out[16];
    assign wire_7984 = lut_tile_4_8_chanxy_out[17];
    assign wire_7986 = lut_tile_4_8_chanxy_out[18];
    assign wire_7988 = lut_tile_4_8_chanxy_out[19];
    assign wire_7990 = lut_tile_4_8_chanxy_out[20];
    assign wire_7992 = lut_tile_4_8_chanxy_out[21];
    assign wire_7994 = lut_tile_4_8_chanxy_out[22];
    assign wire_7996 = lut_tile_4_8_chanxy_out[23];
    assign wire_7998 = lut_tile_4_8_chanxy_out[24];
    assign wire_8000 = lut_tile_4_8_chanxy_out[25];
    assign wire_8002 = lut_tile_4_8_chanxy_out[26];
    assign wire_8004 = lut_tile_4_8_chanxy_out[27];
    assign wire_8006 = lut_tile_4_8_chanxy_out[28];
    assign wire_8008 = lut_tile_4_8_chanxy_out[29];
    assign wire_13531 = lut_tile_4_8_chanxy_out[30];
    assign wire_13539 = lut_tile_4_8_chanxy_out[31];
    assign wire_13547 = lut_tile_4_8_chanxy_out[32];
    assign wire_13555 = lut_tile_4_8_chanxy_out[33];
    assign wire_13563 = lut_tile_4_8_chanxy_out[34];
    assign wire_13571 = lut_tile_4_8_chanxy_out[35];
    assign wire_13579 = lut_tile_4_8_chanxy_out[36];
    assign wire_13587 = lut_tile_4_8_chanxy_out[37];
    assign wire_13595 = lut_tile_4_8_chanxy_out[38];
    assign wire_13603 = lut_tile_4_8_chanxy_out[39];
    assign wire_13611 = lut_tile_4_8_chanxy_out[40];
    assign wire_13619 = lut_tile_4_8_chanxy_out[41];
    assign wire_13627 = lut_tile_4_8_chanxy_out[42];
    assign wire_13635 = lut_tile_4_8_chanxy_out[43];
    assign wire_13643 = lut_tile_4_8_chanxy_out[44];
    assign wire_13710 = lut_tile_4_8_chanxy_out[45];
    assign wire_13712 = lut_tile_4_8_chanxy_out[46];
    assign wire_13714 = lut_tile_4_8_chanxy_out[47];
    assign wire_13716 = lut_tile_4_8_chanxy_out[48];
    assign wire_13718 = lut_tile_4_8_chanxy_out[49];
    assign wire_13720 = lut_tile_4_8_chanxy_out[50];
    assign wire_13722 = lut_tile_4_8_chanxy_out[51];
    assign wire_13724 = lut_tile_4_8_chanxy_out[52];
    assign wire_13726 = lut_tile_4_8_chanxy_out[53];
    assign wire_13728 = lut_tile_4_8_chanxy_out[54];
    assign wire_13730 = lut_tile_4_8_chanxy_out[55];
    assign wire_13732 = lut_tile_4_8_chanxy_out[56];
    assign wire_13734 = lut_tile_4_8_chanxy_out[57];
    assign wire_13736 = lut_tile_4_8_chanxy_out[58];
    assign wire_13738 = lut_tile_4_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_9_chanxy_in = {wire_14032, wire_7651, wire_7649, wire_7648, wire_7639, wire_7638, wire_7629, wire_7628, wire_7532, wire_5331, wire_14024, wire_7679, wire_7619, wire_7618, wire_7609, wire_7608, wire_7599, wire_7598, wire_7534, wire_5331, wire_14016, wire_7677, wire_7589, wire_7588, wire_7579, wire_7578, wire_7569, wire_7568, wire_7536, wire_5331, wire_14008, wire_7675, wire_7647, wire_7646, wire_7637, wire_7636, wire_7627, wire_7626, wire_7538, wire_4821, wire_14000, wire_7673, wire_7617, wire_7616, wire_7607, wire_7606, wire_7597, wire_7596, wire_7540, wire_4821, wire_13992, wire_7671, wire_7587, wire_7586, wire_7577, wire_7576, wire_7567, wire_7566, wire_7542, wire_4821, wire_13984, wire_7669, wire_7645, wire_7644, wire_7635, wire_7634, wire_7625, wire_7624, wire_7544, wire_5335, wire_4821, wire_13976, wire_7667, wire_7615, wire_7614, wire_7605, wire_7604, wire_7595, wire_7594, wire_7546, wire_5335, wire_4821, wire_13968, wire_7665, wire_7585, wire_7584, wire_7575, wire_7574, wire_7565, wire_7564, wire_7548, wire_5335, wire_4821, wire_13960, wire_7663, wire_7643, wire_7642, wire_7633, wire_7632, wire_7623, wire_7622, wire_7550, wire_5335, wire_4817, wire_13952, wire_7661, wire_7613, wire_7612, wire_7603, wire_7602, wire_7593, wire_7592, wire_7552, wire_5335, wire_4817, wire_13944, wire_7659, wire_7583, wire_7582, wire_7573, wire_7572, wire_7563, wire_7562, wire_7554, wire_5335, wire_4817, wire_13936, wire_7657, wire_7641, wire_7640, wire_7631, wire_7630, wire_7621, wire_7620, wire_7556, wire_5331, wire_4817, wire_13928, wire_7655, wire_7611, wire_7610, wire_7601, wire_7600, wire_7591, wire_7590, wire_7558, wire_5331, wire_4817, wire_13920, wire_7653, wire_7581, wire_7580, wire_7571, wire_7570, wire_7561, wire_7560, wire_7530, wire_5331, wire_4817, wire_14159, wire_8069, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7920, wire_5331, wire_14157, wire_8041, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7948, wire_5331, wire_14155, wire_8043, wire_8039, wire_8038, wire_8029, wire_8028, wire_8019, wire_8018, wire_7946, wire_5331, wire_14153, wire_8045, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7944, wire_4821, wire_14151, wire_8047, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7942, wire_4821, wire_14149, wire_8049, wire_8037, wire_8036, wire_8027, wire_8026, wire_8017, wire_8016, wire_7940, wire_4821, wire_14147, wire_8051, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7938, wire_5335, wire_4821, wire_14145, wire_8053, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7936, wire_5335, wire_4821, wire_14143, wire_8055, wire_8035, wire_8034, wire_8025, wire_8024, wire_8015, wire_8014, wire_7934, wire_5335, wire_4821, wire_14141, wire_8057, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7932, wire_5335, wire_4817, wire_14139, wire_8059, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7930, wire_5335, wire_4817, wire_14137, wire_8061, wire_8033, wire_8032, wire_8023, wire_8022, wire_8013, wire_8012, wire_7928, wire_5335, wire_4817, wire_14135, wire_8063, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7926, wire_5331, wire_4817, wire_14133, wire_8065, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7924, wire_5331, wire_4817, wire_14131, wire_8067, wire_8031, wire_8030, wire_8021, wire_8020, wire_8011, wire_8010, wire_7922, wire_5331, wire_4817, wire_13767, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13642, wire_7918, wire_4860, wire_13765, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13530, wire_7916, wire_4860, wire_13763, wire_13679, wire_13678, wire_13669, wire_13668, wire_13659, wire_13658, wire_13538, wire_7914, wire_4860, wire_13761, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13546, wire_7912, wire_4820, wire_13759, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13554, wire_7910, wire_4820, wire_13757, wire_13677, wire_13676, wire_13667, wire_13666, wire_13657, wire_13656, wire_13562, wire_7908, wire_4820, wire_13755, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13570, wire_7906, wire_4864, wire_4820, wire_13753, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13578, wire_7904, wire_4864, wire_4820, wire_13751, wire_13675, wire_13674, wire_13665, wire_13664, wire_13655, wire_13654, wire_13586, wire_7902, wire_4864, wire_4820, wire_13749, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13594, wire_7900, wire_4864, wire_4816, wire_13747, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13602, wire_7898, wire_4864, wire_4816, wire_13745, wire_13673, wire_13672, wire_13663, wire_13662, wire_13653, wire_13652, wire_13610, wire_7896, wire_4864, wire_4816, wire_13743, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13618, wire_7894, wire_4860, wire_4816, wire_13741, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13626, wire_7892, wire_4860, wire_4816, wire_13769, wire_13671, wire_13670, wire_13661, wire_13660, wire_13651, wire_13650, wire_13634, wire_7890, wire_4860, wire_4816, wire_14133, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14026, wire_8069, wire_4860, wire_14135, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_14018, wire_8067, wire_4860, wire_14137, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14010, wire_8065, wire_4860, wire_14139, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14002, wire_8063, wire_4820, wire_14141, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_13994, wire_8061, wire_4820, wire_14143, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_13986, wire_8059, wire_4820, wire_14145, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_13978, wire_8057, wire_4864, wire_4820, wire_14147, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13970, wire_8055, wire_4864, wire_4820, wire_14149, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_13962, wire_8053, wire_4864, wire_4820, wire_14151, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_13954, wire_8051, wire_4864, wire_4816, wire_14153, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13946, wire_8049, wire_4864, wire_4816, wire_14155, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_13938, wire_8047, wire_4864, wire_4816, wire_14157, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_13930, wire_8045, wire_4860, wire_4816, wire_14159, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_13922, wire_8043, wire_4860, wire_4816, wire_14131, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14034, wire_8041, wire_4860, wire_4816};
    // CHNAXY TOTAL: 636
    assign wire_7921 = lut_tile_4_9_chanxy_out[0];
    assign wire_7923 = lut_tile_4_9_chanxy_out[1];
    assign wire_7925 = lut_tile_4_9_chanxy_out[2];
    assign wire_7927 = lut_tile_4_9_chanxy_out[3];
    assign wire_7929 = lut_tile_4_9_chanxy_out[4];
    assign wire_7931 = lut_tile_4_9_chanxy_out[5];
    assign wire_7933 = lut_tile_4_9_chanxy_out[6];
    assign wire_7935 = lut_tile_4_9_chanxy_out[7];
    assign wire_7937 = lut_tile_4_9_chanxy_out[8];
    assign wire_7939 = lut_tile_4_9_chanxy_out[9];
    assign wire_7941 = lut_tile_4_9_chanxy_out[10];
    assign wire_7943 = lut_tile_4_9_chanxy_out[11];
    assign wire_7945 = lut_tile_4_9_chanxy_out[12];
    assign wire_7947 = lut_tile_4_9_chanxy_out[13];
    assign wire_7949 = lut_tile_4_9_chanxy_out[14];
    assign wire_8010 = lut_tile_4_9_chanxy_out[15];
    assign wire_8012 = lut_tile_4_9_chanxy_out[16];
    assign wire_8014 = lut_tile_4_9_chanxy_out[17];
    assign wire_8016 = lut_tile_4_9_chanxy_out[18];
    assign wire_8018 = lut_tile_4_9_chanxy_out[19];
    assign wire_8020 = lut_tile_4_9_chanxy_out[20];
    assign wire_8022 = lut_tile_4_9_chanxy_out[21];
    assign wire_8024 = lut_tile_4_9_chanxy_out[22];
    assign wire_8026 = lut_tile_4_9_chanxy_out[23];
    assign wire_8028 = lut_tile_4_9_chanxy_out[24];
    assign wire_8030 = lut_tile_4_9_chanxy_out[25];
    assign wire_8032 = lut_tile_4_9_chanxy_out[26];
    assign wire_8034 = lut_tile_4_9_chanxy_out[27];
    assign wire_8036 = lut_tile_4_9_chanxy_out[28];
    assign wire_8038 = lut_tile_4_9_chanxy_out[29];
    assign wire_13923 = lut_tile_4_9_chanxy_out[30];
    assign wire_13931 = lut_tile_4_9_chanxy_out[31];
    assign wire_13939 = lut_tile_4_9_chanxy_out[32];
    assign wire_13947 = lut_tile_4_9_chanxy_out[33];
    assign wire_13955 = lut_tile_4_9_chanxy_out[34];
    assign wire_13963 = lut_tile_4_9_chanxy_out[35];
    assign wire_13971 = lut_tile_4_9_chanxy_out[36];
    assign wire_13979 = lut_tile_4_9_chanxy_out[37];
    assign wire_13987 = lut_tile_4_9_chanxy_out[38];
    assign wire_13995 = lut_tile_4_9_chanxy_out[39];
    assign wire_14003 = lut_tile_4_9_chanxy_out[40];
    assign wire_14011 = lut_tile_4_9_chanxy_out[41];
    assign wire_14019 = lut_tile_4_9_chanxy_out[42];
    assign wire_14027 = lut_tile_4_9_chanxy_out[43];
    assign wire_14035 = lut_tile_4_9_chanxy_out[44];
    assign wire_14100 = lut_tile_4_9_chanxy_out[45];
    assign wire_14102 = lut_tile_4_9_chanxy_out[46];
    assign wire_14104 = lut_tile_4_9_chanxy_out[47];
    assign wire_14106 = lut_tile_4_9_chanxy_out[48];
    assign wire_14108 = lut_tile_4_9_chanxy_out[49];
    assign wire_14110 = lut_tile_4_9_chanxy_out[50];
    assign wire_14112 = lut_tile_4_9_chanxy_out[51];
    assign wire_14114 = lut_tile_4_9_chanxy_out[52];
    assign wire_14116 = lut_tile_4_9_chanxy_out[53];
    assign wire_14118 = lut_tile_4_9_chanxy_out[54];
    assign wire_14120 = lut_tile_4_9_chanxy_out[55];
    assign wire_14122 = lut_tile_4_9_chanxy_out[56];
    assign wire_14124 = lut_tile_4_9_chanxy_out[57];
    assign wire_14126 = lut_tile_4_9_chanxy_out[58];
    assign wire_14128 = lut_tile_4_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_4_10_chanxy_in = {wire_14424, wire_7672, wire_7648, wire_7596, wire_7574, wire_5830, wire_5824, wire_5815, wire_5809, wire_14416, wire_7664, wire_7640, wire_7618, wire_7566, wire_5830, wire_5824, wire_5815, wire_5809, wire_14408, wire_7656, wire_7632, wire_7610, wire_7588, wire_5830, wire_5824, wire_5815, wire_5809, wire_14400, wire_7678, wire_7624, wire_7602, wire_7580, wire_5830, wire_5821, wire_5815, wire_5337, wire_14392, wire_7670, wire_7646, wire_7594, wire_7572, wire_5830, wire_5821, wire_5815, wire_5337, wire_14384, wire_7662, wire_7638, wire_7616, wire_7564, wire_5830, wire_5821, wire_5815, wire_5337, wire_14376, wire_7654, wire_7630, wire_7608, wire_7586, wire_5827, wire_5821, wire_5812, wire_5337, wire_14368, wire_7676, wire_7622, wire_7600, wire_7578, wire_5827, wire_5821, wire_5812, wire_5337, wire_14360, wire_7668, wire_7644, wire_7592, wire_7570, wire_5827, wire_5821, wire_5812, wire_5337, wire_14352, wire_7660, wire_7636, wire_7614, wire_7562, wire_5827, wire_5818, wire_5812, wire_5333, wire_14344, wire_7652, wire_7628, wire_7606, wire_7584, wire_5827, wire_5818, wire_5812, wire_5333, wire_14336, wire_7674, wire_7620, wire_7598, wire_7576, wire_5827, wire_5818, wire_5812, wire_5333, wire_14328, wire_7666, wire_7642, wire_7590, wire_7568, wire_5824, wire_5818, wire_5809, wire_5333, wire_14320, wire_7658, wire_7634, wire_7612, wire_7560, wire_5824, wire_5818, wire_5809, wire_5333, wire_14312, wire_7650, wire_7626, wire_7604, wire_7582, wire_5824, wire_5818, wire_5809, wire_5333, wire_14549, wire_8054, wire_8032, wire_8008, wire_7956, wire_5830, wire_5824, wire_5815, wire_5809, wire_14547, wire_8046, wire_8024, wire_8000, wire_7978, wire_5830, wire_5824, wire_5815, wire_5809, wire_14545, wire_8068, wire_8016, wire_7992, wire_7970, wire_5830, wire_5824, wire_5815, wire_5809, wire_14543, wire_8060, wire_8038, wire_7984, wire_7962, wire_5830, wire_5821, wire_5815, wire_5337, wire_14541, wire_8052, wire_8030, wire_8006, wire_7954, wire_5830, wire_5821, wire_5815, wire_5337, wire_14539, wire_8044, wire_8022, wire_7998, wire_7976, wire_5830, wire_5821, wire_5815, wire_5337, wire_14537, wire_8066, wire_8014, wire_7990, wire_7968, wire_5827, wire_5821, wire_5812, wire_5337, wire_14535, wire_8058, wire_8036, wire_7982, wire_7960, wire_5827, wire_5821, wire_5812, wire_5337, wire_14533, wire_8050, wire_8028, wire_8004, wire_7952, wire_5827, wire_5821, wire_5812, wire_5337, wire_14531, wire_8042, wire_8020, wire_7996, wire_7974, wire_5827, wire_5818, wire_5812, wire_5333, wire_14529, wire_8064, wire_8012, wire_7988, wire_7966, wire_5827, wire_5818, wire_5812, wire_5333, wire_14527, wire_8056, wire_8034, wire_7980, wire_7958, wire_5827, wire_5818, wire_5812, wire_5333, wire_14525, wire_8048, wire_8026, wire_8002, wire_7950, wire_5824, wire_5818, wire_5809, wire_5333, wire_14523, wire_8040, wire_8018, wire_7994, wire_7972, wire_5824, wire_5818, wire_5809, wire_5333, wire_14521, wire_8062, wire_8010, wire_7986, wire_7964, wire_5824, wire_5818, wire_5809, wire_5333, wire_14443, wire_14442, wire_14157, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14034, wire_7948, wire_5376, wire_14457, wire_14456, wire_14155, wire_14069, wire_14068, wire_14059, wire_14058, wire_14049, wire_14048, wire_13922, wire_7946, wire_5376, wire_14487, wire_14486, wire_14153, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_13930, wire_7944, wire_5376, wire_14455, wire_14454, wire_14151, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_13938, wire_7942, wire_5336, wire_14439, wire_14438, wire_14149, wire_14067, wire_14066, wire_14057, wire_14056, wire_14047, wire_14046, wire_13946, wire_7940, wire_5336, wire_14469, wire_14468, wire_14147, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_13954, wire_7938, wire_5336, wire_14437, wire_14436, wire_14145, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_13962, wire_7936, wire_5380, wire_5336, wire_14451, wire_14450, wire_14143, wire_14065, wire_14064, wire_14055, wire_14054, wire_14045, wire_14044, wire_13970, wire_7934, wire_5380, wire_5336, wire_14481, wire_14480, wire_14141, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_13978, wire_7932, wire_5380, wire_5336, wire_14449, wire_14448, wire_5380, wire_14139, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_13986, wire_7930, wire_5380, wire_5332, wire_14433, wire_14432, wire_5376, wire_14137, wire_14063, wire_14062, wire_14053, wire_14052, wire_14043, wire_14042, wire_13994, wire_7928, wire_5380, wire_5332, wire_14463, wire_14462, wire_5376, wire_14135, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14002, wire_7926, wire_5380, wire_5332, wire_14431, wire_14430, wire_5336, wire_14133, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14010, wire_7924, wire_5376, wire_5332, wire_14445, wire_14444, wire_5332, wire_14131, wire_14061, wire_14060, wire_14051, wire_14050, wire_14041, wire_14040, wire_14018, wire_7922, wire_5376, wire_5332, wire_14475, wire_14474, wire_5332, wire_14159, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14026, wire_7920, wire_5376, wire_5332, wire_14519, wire_14518, wire_14547, wire_14418, wire_14473, wire_14472, wire_14501, wire_14500, wire_14529, wire_14346, wire_14485, wire_14484, wire_14513, wire_14512, wire_14541, wire_14394, wire_14467, wire_14466, wire_14495, wire_14494, wire_5380, wire_14523, wire_14322, wire_5376, wire_14479, wire_14478, wire_5376, wire_14507, wire_14506, wire_5336, wire_14535, wire_14370, wire_5332, wire_14461, wire_14460, wire_5332, wire_14459, wire_14458, wire_14489, wire_14488, wire_14503, wire_14502, wire_14441, wire_14440, wire_14471, wire_14470, wire_14515, wire_14514, wire_14453, wire_14452, wire_14483, wire_14482, wire_14497, wire_14496, wire_14435, wire_14434, wire_5380, wire_14465, wire_14464, wire_5380, wire_14509, wire_14508, wire_5376, wire_14447, wire_14446, wire_5336, wire_14477, wire_14476, wire_5336, wire_14491, wire_14490, wire_5332, wire_14549, wire_14426, wire_14533, wire_14362, wire_14517, wire_14516, wire_14531, wire_14354, wire_14545, wire_14410, wire_14499, wire_14498, wire_14543, wire_14402, wire_14527, wire_14338, wire_14511, wire_14510, wire_14525, wire_14330, wire_5380, wire_14539, wire_14386, wire_5380, wire_14493, wire_14492, wire_5376, wire_14537, wire_14378, wire_5336, wire_14521, wire_14314, wire_5336, wire_14505, wire_14504, wire_5332};
    // CHNAXY TOTAL: 573
    assign wire_7951 = lut_tile_4_10_chanxy_out[0];
    assign wire_7953 = lut_tile_4_10_chanxy_out[1];
    assign wire_7955 = lut_tile_4_10_chanxy_out[2];
    assign wire_7957 = lut_tile_4_10_chanxy_out[3];
    assign wire_7959 = lut_tile_4_10_chanxy_out[4];
    assign wire_7961 = lut_tile_4_10_chanxy_out[5];
    assign wire_7963 = lut_tile_4_10_chanxy_out[6];
    assign wire_7965 = lut_tile_4_10_chanxy_out[7];
    assign wire_7967 = lut_tile_4_10_chanxy_out[8];
    assign wire_7969 = lut_tile_4_10_chanxy_out[9];
    assign wire_7971 = lut_tile_4_10_chanxy_out[10];
    assign wire_7973 = lut_tile_4_10_chanxy_out[11];
    assign wire_7975 = lut_tile_4_10_chanxy_out[12];
    assign wire_7977 = lut_tile_4_10_chanxy_out[13];
    assign wire_7979 = lut_tile_4_10_chanxy_out[14];
    assign wire_7981 = lut_tile_4_10_chanxy_out[15];
    assign wire_7983 = lut_tile_4_10_chanxy_out[16];
    assign wire_7985 = lut_tile_4_10_chanxy_out[17];
    assign wire_7987 = lut_tile_4_10_chanxy_out[18];
    assign wire_7989 = lut_tile_4_10_chanxy_out[19];
    assign wire_7991 = lut_tile_4_10_chanxy_out[20];
    assign wire_7993 = lut_tile_4_10_chanxy_out[21];
    assign wire_7995 = lut_tile_4_10_chanxy_out[22];
    assign wire_7997 = lut_tile_4_10_chanxy_out[23];
    assign wire_7999 = lut_tile_4_10_chanxy_out[24];
    assign wire_8001 = lut_tile_4_10_chanxy_out[25];
    assign wire_8003 = lut_tile_4_10_chanxy_out[26];
    assign wire_8005 = lut_tile_4_10_chanxy_out[27];
    assign wire_8007 = lut_tile_4_10_chanxy_out[28];
    assign wire_8009 = lut_tile_4_10_chanxy_out[29];
    assign wire_8011 = lut_tile_4_10_chanxy_out[30];
    assign wire_8013 = lut_tile_4_10_chanxy_out[31];
    assign wire_8015 = lut_tile_4_10_chanxy_out[32];
    assign wire_8017 = lut_tile_4_10_chanxy_out[33];
    assign wire_8019 = lut_tile_4_10_chanxy_out[34];
    assign wire_8021 = lut_tile_4_10_chanxy_out[35];
    assign wire_8023 = lut_tile_4_10_chanxy_out[36];
    assign wire_8025 = lut_tile_4_10_chanxy_out[37];
    assign wire_8027 = lut_tile_4_10_chanxy_out[38];
    assign wire_8029 = lut_tile_4_10_chanxy_out[39];
    assign wire_8031 = lut_tile_4_10_chanxy_out[40];
    assign wire_8033 = lut_tile_4_10_chanxy_out[41];
    assign wire_8035 = lut_tile_4_10_chanxy_out[42];
    assign wire_8037 = lut_tile_4_10_chanxy_out[43];
    assign wire_8039 = lut_tile_4_10_chanxy_out[44];
    assign wire_8040 = lut_tile_4_10_chanxy_out[45];
    assign wire_8041 = lut_tile_4_10_chanxy_out[46];
    assign wire_8042 = lut_tile_4_10_chanxy_out[47];
    assign wire_8043 = lut_tile_4_10_chanxy_out[48];
    assign wire_8044 = lut_tile_4_10_chanxy_out[49];
    assign wire_8045 = lut_tile_4_10_chanxy_out[50];
    assign wire_8046 = lut_tile_4_10_chanxy_out[51];
    assign wire_8047 = lut_tile_4_10_chanxy_out[52];
    assign wire_8048 = lut_tile_4_10_chanxy_out[53];
    assign wire_8049 = lut_tile_4_10_chanxy_out[54];
    assign wire_8050 = lut_tile_4_10_chanxy_out[55];
    assign wire_8051 = lut_tile_4_10_chanxy_out[56];
    assign wire_8052 = lut_tile_4_10_chanxy_out[57];
    assign wire_8053 = lut_tile_4_10_chanxy_out[58];
    assign wire_8054 = lut_tile_4_10_chanxy_out[59];
    assign wire_8055 = lut_tile_4_10_chanxy_out[60];
    assign wire_8056 = lut_tile_4_10_chanxy_out[61];
    assign wire_8057 = lut_tile_4_10_chanxy_out[62];
    assign wire_8058 = lut_tile_4_10_chanxy_out[63];
    assign wire_8059 = lut_tile_4_10_chanxy_out[64];
    assign wire_8060 = lut_tile_4_10_chanxy_out[65];
    assign wire_8061 = lut_tile_4_10_chanxy_out[66];
    assign wire_8062 = lut_tile_4_10_chanxy_out[67];
    assign wire_8063 = lut_tile_4_10_chanxy_out[68];
    assign wire_8064 = lut_tile_4_10_chanxy_out[69];
    assign wire_8065 = lut_tile_4_10_chanxy_out[70];
    assign wire_8066 = lut_tile_4_10_chanxy_out[71];
    assign wire_8067 = lut_tile_4_10_chanxy_out[72];
    assign wire_8068 = lut_tile_4_10_chanxy_out[73];
    assign wire_8069 = lut_tile_4_10_chanxy_out[74];
    assign wire_14315 = lut_tile_4_10_chanxy_out[75];
    assign wire_14323 = lut_tile_4_10_chanxy_out[76];
    assign wire_14331 = lut_tile_4_10_chanxy_out[77];
    assign wire_14339 = lut_tile_4_10_chanxy_out[78];
    assign wire_14347 = lut_tile_4_10_chanxy_out[79];
    assign wire_14355 = lut_tile_4_10_chanxy_out[80];
    assign wire_14363 = lut_tile_4_10_chanxy_out[81];
    assign wire_14371 = lut_tile_4_10_chanxy_out[82];
    assign wire_14379 = lut_tile_4_10_chanxy_out[83];
    assign wire_14387 = lut_tile_4_10_chanxy_out[84];
    assign wire_14395 = lut_tile_4_10_chanxy_out[85];
    assign wire_14403 = lut_tile_4_10_chanxy_out[86];
    assign wire_14411 = lut_tile_4_10_chanxy_out[87];
    assign wire_14419 = lut_tile_4_10_chanxy_out[88];
    assign wire_14427 = lut_tile_4_10_chanxy_out[89];
    assign wire_14490 = lut_tile_4_10_chanxy_out[90];
    assign wire_14492 = lut_tile_4_10_chanxy_out[91];
    assign wire_14494 = lut_tile_4_10_chanxy_out[92];
    assign wire_14496 = lut_tile_4_10_chanxy_out[93];
    assign wire_14498 = lut_tile_4_10_chanxy_out[94];
    assign wire_14500 = lut_tile_4_10_chanxy_out[95];
    assign wire_14502 = lut_tile_4_10_chanxy_out[96];
    assign wire_14504 = lut_tile_4_10_chanxy_out[97];
    assign wire_14506 = lut_tile_4_10_chanxy_out[98];
    assign wire_14508 = lut_tile_4_10_chanxy_out[99];
    assign wire_14510 = lut_tile_4_10_chanxy_out[100];
    assign wire_14512 = lut_tile_4_10_chanxy_out[101];
    assign wire_14514 = lut_tile_4_10_chanxy_out[102];
    assign wire_14516 = lut_tile_4_10_chanxy_out[103];
    assign wire_14518 = lut_tile_4_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_5_1_chanxy_in = {wire_10914, wire_7801, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_7690, wire_1245, wire_10906, wire_7829, wire_7797, wire_7796, wire_7757, wire_7756, wire_7717, wire_7716, wire_7698, wire_1245, wire_10898, wire_7827, wire_7793, wire_7792, wire_7753, wire_7752, wire_7713, wire_7712, wire_7706, wire_1245, wire_10890, wire_7825, wire_7791, wire_7790, wire_7751, wire_7750, wire_7714, wire_7711, wire_7710, wire_735, wire_10882, wire_7823, wire_7789, wire_7788, wire_7749, wire_7748, wire_7722, wire_7709, wire_7708, wire_735, wire_10874, wire_7821, wire_7785, wire_7784, wire_7745, wire_7744, wire_7730, wire_7705, wire_7704, wire_735, wire_10866, wire_7819, wire_7783, wire_7782, wire_7743, wire_7742, wire_7738, wire_7703, wire_7702, wire_1249, wire_735, wire_10858, wire_7817, wire_7781, wire_7780, wire_7746, wire_7741, wire_7740, wire_7701, wire_7700, wire_1249, wire_735, wire_10850, wire_7815, wire_7777, wire_7776, wire_7754, wire_7737, wire_7736, wire_7697, wire_7696, wire_1249, wire_735, wire_10842, wire_7813, wire_7775, wire_7774, wire_7762, wire_7735, wire_7734, wire_7695, wire_7694, wire_1249, wire_731, wire_10834, wire_7811, wire_7773, wire_7772, wire_7770, wire_7733, wire_7732, wire_7693, wire_7692, wire_1249, wire_731, wire_10826, wire_7809, wire_7778, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_1249, wire_731, wire_10818, wire_7807, wire_7786, wire_7767, wire_7766, wire_7727, wire_7726, wire_7687, wire_7686, wire_1245, wire_731, wire_10810, wire_7805, wire_7794, wire_7765, wire_7764, wire_7725, wire_7724, wire_7685, wire_7684, wire_1245, wire_731, wire_10802, wire_7803, wire_7761, wire_7760, wire_7721, wire_7720, wire_7682, wire_7681, wire_7680, wire_1245, wire_731, wire_11069, wire_8219, wire_8189, wire_8188, wire_8149, wire_8148, wire_8109, wire_8108, wire_8074, wire_1245, wire_11067, wire_8191, wire_8186, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_1245, wire_11065, wire_8193, wire_8183, wire_8182, wire_8178, wire_8143, wire_8142, wire_8103, wire_8102, wire_1245, wire_11063, wire_8195, wire_8181, wire_8180, wire_8170, wire_8141, wire_8140, wire_8101, wire_8100, wire_735, wire_11061, wire_8197, wire_8177, wire_8176, wire_8162, wire_8137, wire_8136, wire_8097, wire_8096, wire_735, wire_11059, wire_8199, wire_8175, wire_8174, wire_8154, wire_8135, wire_8134, wire_8095, wire_8094, wire_735, wire_11057, wire_8201, wire_8173, wire_8172, wire_8146, wire_8133, wire_8132, wire_8093, wire_8092, wire_1249, wire_735, wire_11055, wire_8203, wire_8169, wire_8168, wire_8138, wire_8129, wire_8128, wire_8089, wire_8088, wire_1249, wire_735, wire_11053, wire_8205, wire_8167, wire_8166, wire_8130, wire_8127, wire_8126, wire_8087, wire_8086, wire_1249, wire_735, wire_11051, wire_8207, wire_8165, wire_8164, wire_8125, wire_8124, wire_8122, wire_8085, wire_8084, wire_1249, wire_731, wire_11049, wire_8209, wire_8161, wire_8160, wire_8121, wire_8120, wire_8114, wire_8081, wire_8080, wire_1249, wire_731, wire_11047, wire_8211, wire_8159, wire_8158, wire_8119, wire_8118, wire_8106, wire_8079, wire_8078, wire_1249, wire_731, wire_11045, wire_8213, wire_8157, wire_8156, wire_8117, wire_8116, wire_8098, wire_8077, wire_8076, wire_1245, wire_731, wire_11043, wire_8215, wire_8153, wire_8152, wire_8113, wire_8112, wire_8090, wire_8073, wire_8072, wire_1245, wire_731, wire_11041, wire_8217, wire_8151, wire_8150, wire_8111, wire_8110, wire_8082, wire_8071, wire_8070, wire_1245, wire_731, wire_10603, wire_10602, wire_11043, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10946, wire_8219, wire_774, wire_10619, wire_10618, wire_10589, wire_10588, wire_10573, wire_10572, wire_10679, wire_10558, wire_11045, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10944, wire_8217, wire_774, wire_10649, wire_10648, wire_10663, wire_10542, wire_10617, wire_10616, wire_10587, wire_10586, wire_11047, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10942, wire_8215, wire_774, wire_10633, wire_10632, wire_10677, wire_10556, wire_10647, wire_10646, wire_10615, wire_10614, wire_11049, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10940, wire_8213, wire_734, wire_10601, wire_10600, wire_10571, wire_10570, wire_10585, wire_10584, wire_10661, wire_10540, wire_11051, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10938, wire_8211, wire_734, wire_10631, wire_10630, wire_10675, wire_10554, wire_10599, wire_10598, wire_10569, wire_10568, wire_11053, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10936, wire_8209, wire_734, wire_10645, wire_10644, wire_10659, wire_10538, wire_10629, wire_10628, wire_10597, wire_10596, wire_11055, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10934, wire_8207, wire_778, wire_734, wire_10613, wire_10612, wire_10583, wire_10582, wire_10567, wire_10566, wire_10673, wire_10552, wire_11057, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10932, wire_8205, wire_778, wire_734, wire_10643, wire_10642, wire_10657, wire_10536, wire_10611, wire_10610, wire_10581, wire_10580, wire_11059, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10930, wire_8203, wire_778, wire_734, wire_10627, wire_10626, wire_10671, wire_10550, wire_10641, wire_10640, wire_10609, wire_10608, wire_778, wire_11061, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10928, wire_8201, wire_778, wire_730, wire_10595, wire_10594, wire_778, wire_10565, wire_10564, wire_778, wire_10579, wire_10578, wire_778, wire_10655, wire_10534, wire_778, wire_11063, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10926, wire_8199, wire_778, wire_730, wire_10625, wire_10624, wire_778, wire_10669, wire_10548, wire_774, wire_10593, wire_10592, wire_774, wire_10563, wire_10562, wire_774, wire_11065, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10924, wire_8197, wire_778, wire_730, wire_10639, wire_10638, wire_774, wire_10653, wire_10532, wire_774, wire_10623, wire_10622, wire_774, wire_10591, wire_10590, wire_734, wire_11067, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10922, wire_8195, wire_774, wire_730, wire_10607, wire_10606, wire_734, wire_10577, wire_10576, wire_734, wire_10561, wire_10560, wire_734, wire_10667, wire_10546, wire_734, wire_11069, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10920, wire_8193, wire_774, wire_730, wire_10637, wire_10636, wire_734, wire_10651, wire_10530, wire_730, wire_10605, wire_10604, wire_730, wire_10575, wire_10574, wire_730, wire_11041, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10948, wire_8191, wire_774, wire_730, wire_10621, wire_10620, wire_730, wire_10665, wire_10544, wire_730, wire_10635, wire_10634, wire_730};
    // CHNAXY TOTAL: 621
    assign wire_8070 = lut_tile_5_1_chanxy_out[0];
    assign wire_8072 = lut_tile_5_1_chanxy_out[1];
    assign wire_8074 = lut_tile_5_1_chanxy_out[2];
    assign wire_8075 = lut_tile_5_1_chanxy_out[3];
    assign wire_8076 = lut_tile_5_1_chanxy_out[4];
    assign wire_8078 = lut_tile_5_1_chanxy_out[5];
    assign wire_8080 = lut_tile_5_1_chanxy_out[6];
    assign wire_8082 = lut_tile_5_1_chanxy_out[7];
    assign wire_8083 = lut_tile_5_1_chanxy_out[8];
    assign wire_8084 = lut_tile_5_1_chanxy_out[9];
    assign wire_8086 = lut_tile_5_1_chanxy_out[10];
    assign wire_8088 = lut_tile_5_1_chanxy_out[11];
    assign wire_8090 = lut_tile_5_1_chanxy_out[12];
    assign wire_8091 = lut_tile_5_1_chanxy_out[13];
    assign wire_8092 = lut_tile_5_1_chanxy_out[14];
    assign wire_8094 = lut_tile_5_1_chanxy_out[15];
    assign wire_8096 = lut_tile_5_1_chanxy_out[16];
    assign wire_8098 = lut_tile_5_1_chanxy_out[17];
    assign wire_8099 = lut_tile_5_1_chanxy_out[18];
    assign wire_8100 = lut_tile_5_1_chanxy_out[19];
    assign wire_8102 = lut_tile_5_1_chanxy_out[20];
    assign wire_8104 = lut_tile_5_1_chanxy_out[21];
    assign wire_8106 = lut_tile_5_1_chanxy_out[22];
    assign wire_8107 = lut_tile_5_1_chanxy_out[23];
    assign wire_8108 = lut_tile_5_1_chanxy_out[24];
    assign wire_8110 = lut_tile_5_1_chanxy_out[25];
    assign wire_8112 = lut_tile_5_1_chanxy_out[26];
    assign wire_8114 = lut_tile_5_1_chanxy_out[27];
    assign wire_8115 = lut_tile_5_1_chanxy_out[28];
    assign wire_8116 = lut_tile_5_1_chanxy_out[29];
    assign wire_8118 = lut_tile_5_1_chanxy_out[30];
    assign wire_8120 = lut_tile_5_1_chanxy_out[31];
    assign wire_8122 = lut_tile_5_1_chanxy_out[32];
    assign wire_8123 = lut_tile_5_1_chanxy_out[33];
    assign wire_8124 = lut_tile_5_1_chanxy_out[34];
    assign wire_8126 = lut_tile_5_1_chanxy_out[35];
    assign wire_8128 = lut_tile_5_1_chanxy_out[36];
    assign wire_8130 = lut_tile_5_1_chanxy_out[37];
    assign wire_8131 = lut_tile_5_1_chanxy_out[38];
    assign wire_8132 = lut_tile_5_1_chanxy_out[39];
    assign wire_8134 = lut_tile_5_1_chanxy_out[40];
    assign wire_8136 = lut_tile_5_1_chanxy_out[41];
    assign wire_8138 = lut_tile_5_1_chanxy_out[42];
    assign wire_8139 = lut_tile_5_1_chanxy_out[43];
    assign wire_8140 = lut_tile_5_1_chanxy_out[44];
    assign wire_8142 = lut_tile_5_1_chanxy_out[45];
    assign wire_8144 = lut_tile_5_1_chanxy_out[46];
    assign wire_8146 = lut_tile_5_1_chanxy_out[47];
    assign wire_8147 = lut_tile_5_1_chanxy_out[48];
    assign wire_8148 = lut_tile_5_1_chanxy_out[49];
    assign wire_8150 = lut_tile_5_1_chanxy_out[50];
    assign wire_8152 = lut_tile_5_1_chanxy_out[51];
    assign wire_8154 = lut_tile_5_1_chanxy_out[52];
    assign wire_8155 = lut_tile_5_1_chanxy_out[53];
    assign wire_8156 = lut_tile_5_1_chanxy_out[54];
    assign wire_8158 = lut_tile_5_1_chanxy_out[55];
    assign wire_8160 = lut_tile_5_1_chanxy_out[56];
    assign wire_8162 = lut_tile_5_1_chanxy_out[57];
    assign wire_8163 = lut_tile_5_1_chanxy_out[58];
    assign wire_8164 = lut_tile_5_1_chanxy_out[59];
    assign wire_8166 = lut_tile_5_1_chanxy_out[60];
    assign wire_8168 = lut_tile_5_1_chanxy_out[61];
    assign wire_8170 = lut_tile_5_1_chanxy_out[62];
    assign wire_8171 = lut_tile_5_1_chanxy_out[63];
    assign wire_8172 = lut_tile_5_1_chanxy_out[64];
    assign wire_8174 = lut_tile_5_1_chanxy_out[65];
    assign wire_8176 = lut_tile_5_1_chanxy_out[66];
    assign wire_8178 = lut_tile_5_1_chanxy_out[67];
    assign wire_8179 = lut_tile_5_1_chanxy_out[68];
    assign wire_8180 = lut_tile_5_1_chanxy_out[69];
    assign wire_8182 = lut_tile_5_1_chanxy_out[70];
    assign wire_8184 = lut_tile_5_1_chanxy_out[71];
    assign wire_8186 = lut_tile_5_1_chanxy_out[72];
    assign wire_8187 = lut_tile_5_1_chanxy_out[73];
    assign wire_8188 = lut_tile_5_1_chanxy_out[74];
    assign wire_10921 = lut_tile_5_1_chanxy_out[75];
    assign wire_10923 = lut_tile_5_1_chanxy_out[76];
    assign wire_10925 = lut_tile_5_1_chanxy_out[77];
    assign wire_10927 = lut_tile_5_1_chanxy_out[78];
    assign wire_10929 = lut_tile_5_1_chanxy_out[79];
    assign wire_10931 = lut_tile_5_1_chanxy_out[80];
    assign wire_10933 = lut_tile_5_1_chanxy_out[81];
    assign wire_10935 = lut_tile_5_1_chanxy_out[82];
    assign wire_10937 = lut_tile_5_1_chanxy_out[83];
    assign wire_10939 = lut_tile_5_1_chanxy_out[84];
    assign wire_10941 = lut_tile_5_1_chanxy_out[85];
    assign wire_10943 = lut_tile_5_1_chanxy_out[86];
    assign wire_10945 = lut_tile_5_1_chanxy_out[87];
    assign wire_10947 = lut_tile_5_1_chanxy_out[88];
    assign wire_10949 = lut_tile_5_1_chanxy_out[89];
    assign wire_11010 = lut_tile_5_1_chanxy_out[90];
    assign wire_11012 = lut_tile_5_1_chanxy_out[91];
    assign wire_11014 = lut_tile_5_1_chanxy_out[92];
    assign wire_11016 = lut_tile_5_1_chanxy_out[93];
    assign wire_11018 = lut_tile_5_1_chanxy_out[94];
    assign wire_11020 = lut_tile_5_1_chanxy_out[95];
    assign wire_11022 = lut_tile_5_1_chanxy_out[96];
    assign wire_11024 = lut_tile_5_1_chanxy_out[97];
    assign wire_11026 = lut_tile_5_1_chanxy_out[98];
    assign wire_11028 = lut_tile_5_1_chanxy_out[99];
    assign wire_11030 = lut_tile_5_1_chanxy_out[100];
    assign wire_11032 = lut_tile_5_1_chanxy_out[101];
    assign wire_11034 = lut_tile_5_1_chanxy_out[102];
    assign wire_11036 = lut_tile_5_1_chanxy_out[103];
    assign wire_11038 = lut_tile_5_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_5_2_chanxy_in = {wire_11306, wire_7831, wire_7799, wire_7798, wire_7759, wire_7758, wire_7719, wire_7718, wire_7692, wire_1761, wire_11298, wire_7859, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7700, wire_1761, wire_11290, wire_7857, wire_7793, wire_7792, wire_7753, wire_7752, wire_7713, wire_7712, wire_7708, wire_1761, wire_11282, wire_7855, wire_7791, wire_7790, wire_7751, wire_7750, wire_7716, wire_7711, wire_7710, wire_1251, wire_11274, wire_7853, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7724, wire_1251, wire_11266, wire_7851, wire_7785, wire_7784, wire_7745, wire_7744, wire_7732, wire_7705, wire_7704, wire_1251, wire_11258, wire_7849, wire_7783, wire_7782, wire_7743, wire_7742, wire_7740, wire_7703, wire_7702, wire_1765, wire_1251, wire_11250, wire_7847, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7748, wire_1765, wire_1251, wire_11242, wire_7845, wire_7777, wire_7776, wire_7756, wire_7737, wire_7736, wire_7697, wire_7696, wire_1765, wire_1251, wire_11234, wire_7843, wire_7775, wire_7774, wire_7764, wire_7735, wire_7734, wire_7695, wire_7694, wire_1765, wire_1247, wire_11226, wire_7841, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7772, wire_1765, wire_1247, wire_11218, wire_7839, wire_7780, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_1765, wire_1247, wire_11210, wire_7837, wire_7788, wire_7767, wire_7766, wire_7727, wire_7726, wire_7687, wire_7686, wire_1761, wire_1247, wire_11202, wire_7835, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7796, wire_1761, wire_1247, wire_11194, wire_7833, wire_7761, wire_7760, wire_7721, wire_7720, wire_7684, wire_7681, wire_7680, wire_1761, wire_1247, wire_11459, wire_8249, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8076, wire_1761, wire_11457, wire_8221, wire_8188, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_1761, wire_11455, wire_8223, wire_8183, wire_8182, wire_8180, wire_8143, wire_8142, wire_8103, wire_8102, wire_1761, wire_11453, wire_8225, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8172, wire_1251, wire_11451, wire_8227, wire_8177, wire_8176, wire_8164, wire_8137, wire_8136, wire_8097, wire_8096, wire_1251, wire_11449, wire_8229, wire_8175, wire_8174, wire_8156, wire_8135, wire_8134, wire_8095, wire_8094, wire_1251, wire_11447, wire_8231, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8148, wire_1765, wire_1251, wire_11445, wire_8233, wire_8169, wire_8168, wire_8140, wire_8129, wire_8128, wire_8089, wire_8088, wire_1765, wire_1251, wire_11443, wire_8235, wire_8167, wire_8166, wire_8132, wire_8127, wire_8126, wire_8087, wire_8086, wire_1765, wire_1251, wire_11441, wire_8237, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8124, wire_1765, wire_1247, wire_11439, wire_8239, wire_8161, wire_8160, wire_8121, wire_8120, wire_8116, wire_8081, wire_8080, wire_1765, wire_1247, wire_11437, wire_8241, wire_8159, wire_8158, wire_8119, wire_8118, wire_8108, wire_8079, wire_8078, wire_1765, wire_1247, wire_11435, wire_8243, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8100, wire_1761, wire_1247, wire_11433, wire_8245, wire_8153, wire_8152, wire_8113, wire_8112, wire_8092, wire_8073, wire_8072, wire_1761, wire_1247, wire_11431, wire_8247, wire_8151, wire_8150, wire_8111, wire_8110, wire_8084, wire_8071, wire_8070, wire_1761, wire_1247, wire_11067, wire_10979, wire_10978, wire_10969, wire_10968, wire_10959, wire_10958, wire_10948, wire_8186, wire_1290, wire_11065, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10920, wire_8178, wire_1290, wire_11063, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10922, wire_8170, wire_1290, wire_11061, wire_10977, wire_10976, wire_10967, wire_10966, wire_10957, wire_10956, wire_10924, wire_8162, wire_1250, wire_11059, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10926, wire_8154, wire_1250, wire_11057, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10928, wire_8146, wire_1250, wire_11055, wire_10975, wire_10974, wire_10965, wire_10964, wire_10955, wire_10954, wire_10930, wire_8138, wire_1294, wire_1250, wire_11053, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10932, wire_8130, wire_1294, wire_1250, wire_11051, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10934, wire_8122, wire_1294, wire_1250, wire_11049, wire_10973, wire_10972, wire_10963, wire_10962, wire_10953, wire_10952, wire_10936, wire_8114, wire_1294, wire_1246, wire_11047, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10938, wire_8106, wire_1294, wire_1246, wire_11045, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10940, wire_8098, wire_1294, wire_1246, wire_11043, wire_10971, wire_10970, wire_10961, wire_10960, wire_10951, wire_10950, wire_10942, wire_8090, wire_1290, wire_1246, wire_11041, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10944, wire_8082, wire_1290, wire_1246, wire_11069, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10946, wire_8074, wire_1290, wire_1246, wire_11433, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11336, wire_8249, wire_1290, wire_11435, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11334, wire_8247, wire_1290, wire_11437, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11332, wire_8245, wire_1290, wire_11439, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11330, wire_8243, wire_1250, wire_11441, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11328, wire_8241, wire_1250, wire_11443, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11326, wire_8239, wire_1250, wire_11445, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11324, wire_8237, wire_1294, wire_1250, wire_11447, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11322, wire_8235, wire_1294, wire_1250, wire_11449, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11320, wire_8233, wire_1294, wire_1250, wire_11451, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11318, wire_8231, wire_1294, wire_1246, wire_11453, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11316, wire_8229, wire_1294, wire_1246, wire_11455, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11314, wire_8227, wire_1294, wire_1246, wire_11457, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11312, wire_8225, wire_1290, wire_1246, wire_11459, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11310, wire_8223, wire_1290, wire_1246, wire_11431, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11338, wire_8221, wire_1290, wire_1246};
    // CHNAXY TOTAL: 636
    assign wire_8077 = lut_tile_5_2_chanxy_out[0];
    assign wire_8085 = lut_tile_5_2_chanxy_out[1];
    assign wire_8093 = lut_tile_5_2_chanxy_out[2];
    assign wire_8101 = lut_tile_5_2_chanxy_out[3];
    assign wire_8109 = lut_tile_5_2_chanxy_out[4];
    assign wire_8117 = lut_tile_5_2_chanxy_out[5];
    assign wire_8125 = lut_tile_5_2_chanxy_out[6];
    assign wire_8133 = lut_tile_5_2_chanxy_out[7];
    assign wire_8141 = lut_tile_5_2_chanxy_out[8];
    assign wire_8149 = lut_tile_5_2_chanxy_out[9];
    assign wire_8157 = lut_tile_5_2_chanxy_out[10];
    assign wire_8165 = lut_tile_5_2_chanxy_out[11];
    assign wire_8173 = lut_tile_5_2_chanxy_out[12];
    assign wire_8181 = lut_tile_5_2_chanxy_out[13];
    assign wire_8189 = lut_tile_5_2_chanxy_out[14];
    assign wire_8190 = lut_tile_5_2_chanxy_out[15];
    assign wire_8192 = lut_tile_5_2_chanxy_out[16];
    assign wire_8194 = lut_tile_5_2_chanxy_out[17];
    assign wire_8196 = lut_tile_5_2_chanxy_out[18];
    assign wire_8198 = lut_tile_5_2_chanxy_out[19];
    assign wire_8200 = lut_tile_5_2_chanxy_out[20];
    assign wire_8202 = lut_tile_5_2_chanxy_out[21];
    assign wire_8204 = lut_tile_5_2_chanxy_out[22];
    assign wire_8206 = lut_tile_5_2_chanxy_out[23];
    assign wire_8208 = lut_tile_5_2_chanxy_out[24];
    assign wire_8210 = lut_tile_5_2_chanxy_out[25];
    assign wire_8212 = lut_tile_5_2_chanxy_out[26];
    assign wire_8214 = lut_tile_5_2_chanxy_out[27];
    assign wire_8216 = lut_tile_5_2_chanxy_out[28];
    assign wire_8218 = lut_tile_5_2_chanxy_out[29];
    assign wire_11311 = lut_tile_5_2_chanxy_out[30];
    assign wire_11313 = lut_tile_5_2_chanxy_out[31];
    assign wire_11315 = lut_tile_5_2_chanxy_out[32];
    assign wire_11317 = lut_tile_5_2_chanxy_out[33];
    assign wire_11319 = lut_tile_5_2_chanxy_out[34];
    assign wire_11321 = lut_tile_5_2_chanxy_out[35];
    assign wire_11323 = lut_tile_5_2_chanxy_out[36];
    assign wire_11325 = lut_tile_5_2_chanxy_out[37];
    assign wire_11327 = lut_tile_5_2_chanxy_out[38];
    assign wire_11329 = lut_tile_5_2_chanxy_out[39];
    assign wire_11331 = lut_tile_5_2_chanxy_out[40];
    assign wire_11333 = lut_tile_5_2_chanxy_out[41];
    assign wire_11335 = lut_tile_5_2_chanxy_out[42];
    assign wire_11337 = lut_tile_5_2_chanxy_out[43];
    assign wire_11339 = lut_tile_5_2_chanxy_out[44];
    assign wire_11400 = lut_tile_5_2_chanxy_out[45];
    assign wire_11402 = lut_tile_5_2_chanxy_out[46];
    assign wire_11404 = lut_tile_5_2_chanxy_out[47];
    assign wire_11406 = lut_tile_5_2_chanxy_out[48];
    assign wire_11408 = lut_tile_5_2_chanxy_out[49];
    assign wire_11410 = lut_tile_5_2_chanxy_out[50];
    assign wire_11412 = lut_tile_5_2_chanxy_out[51];
    assign wire_11414 = lut_tile_5_2_chanxy_out[52];
    assign wire_11416 = lut_tile_5_2_chanxy_out[53];
    assign wire_11418 = lut_tile_5_2_chanxy_out[54];
    assign wire_11420 = lut_tile_5_2_chanxy_out[55];
    assign wire_11422 = lut_tile_5_2_chanxy_out[56];
    assign wire_11424 = lut_tile_5_2_chanxy_out[57];
    assign wire_11426 = lut_tile_5_2_chanxy_out[58];
    assign wire_11428 = lut_tile_5_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_3_chanxy_in = {wire_11698, wire_7861, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7694, wire_2277, wire_11690, wire_7889, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7702, wire_2277, wire_11682, wire_7887, wire_7793, wire_7792, wire_7753, wire_7752, wire_7713, wire_7712, wire_7710, wire_2277, wire_11674, wire_7885, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7718, wire_1767, wire_11666, wire_7883, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7726, wire_1767, wire_11658, wire_7881, wire_7785, wire_7784, wire_7745, wire_7744, wire_7734, wire_7705, wire_7704, wire_1767, wire_11650, wire_7879, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7742, wire_2281, wire_1767, wire_11642, wire_7877, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7750, wire_2281, wire_1767, wire_11634, wire_7875, wire_7777, wire_7776, wire_7758, wire_7737, wire_7736, wire_7697, wire_7696, wire_2281, wire_1767, wire_11626, wire_7873, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7766, wire_2281, wire_1763, wire_11618, wire_7871, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7774, wire_2281, wire_1763, wire_11610, wire_7869, wire_7782, wire_7769, wire_7768, wire_7729, wire_7728, wire_7689, wire_7688, wire_2281, wire_1763, wire_11602, wire_7867, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7790, wire_2277, wire_1763, wire_11594, wire_7865, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7798, wire_2277, wire_1763, wire_11586, wire_7863, wire_7761, wire_7760, wire_7721, wire_7720, wire_7686, wire_7681, wire_7680, wire_2277, wire_1763, wire_11849, wire_8279, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8070, wire_2277, wire_11847, wire_8251, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8182, wire_2277, wire_11845, wire_8253, wire_8185, wire_8184, wire_8174, wire_8145, wire_8144, wire_8105, wire_8104, wire_2277, wire_11843, wire_8255, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8166, wire_1767, wire_11841, wire_8257, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8158, wire_1767, wire_11839, wire_8259, wire_8177, wire_8176, wire_8150, wire_8137, wire_8136, wire_8097, wire_8096, wire_1767, wire_11837, wire_8261, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8142, wire_2281, wire_1767, wire_11835, wire_8263, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8134, wire_2281, wire_1767, wire_11833, wire_8265, wire_8169, wire_8168, wire_8129, wire_8128, wire_8126, wire_8089, wire_8088, wire_2281, wire_1767, wire_11831, wire_8267, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8118, wire_2281, wire_1763, wire_11829, wire_8269, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8110, wire_2281, wire_1763, wire_11827, wire_8271, wire_8161, wire_8160, wire_8121, wire_8120, wire_8102, wire_8081, wire_8080, wire_2281, wire_1763, wire_11825, wire_8273, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8094, wire_2277, wire_1763, wire_11823, wire_8275, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8086, wire_2277, wire_1763, wire_11821, wire_8277, wire_8153, wire_8152, wire_8113, wire_8112, wire_8078, wire_8073, wire_8072, wire_2277, wire_1763, wire_11457, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11338, wire_8188, wire_1806, wire_11455, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11310, wire_8180, wire_1806, wire_11453, wire_11369, wire_11368, wire_11359, wire_11358, wire_11349, wire_11348, wire_11312, wire_8172, wire_1806, wire_11451, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11314, wire_8164, wire_1766, wire_11449, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11316, wire_8156, wire_1766, wire_11447, wire_11367, wire_11366, wire_11357, wire_11356, wire_11347, wire_11346, wire_11318, wire_8148, wire_1766, wire_11445, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11320, wire_8140, wire_1810, wire_1766, wire_11443, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11322, wire_8132, wire_1810, wire_1766, wire_11441, wire_11365, wire_11364, wire_11355, wire_11354, wire_11345, wire_11344, wire_11324, wire_8124, wire_1810, wire_1766, wire_11439, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11326, wire_8116, wire_1810, wire_1762, wire_11437, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11328, wire_8108, wire_1810, wire_1762, wire_11435, wire_11363, wire_11362, wire_11353, wire_11352, wire_11343, wire_11342, wire_11330, wire_8100, wire_1810, wire_1762, wire_11433, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11332, wire_8092, wire_1806, wire_1762, wire_11431, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11334, wire_8084, wire_1806, wire_1762, wire_11459, wire_11361, wire_11360, wire_11351, wire_11350, wire_11341, wire_11340, wire_11336, wire_8076, wire_1806, wire_1762, wire_11823, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11726, wire_8279, wire_1806, wire_11825, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11724, wire_8277, wire_1806, wire_11827, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11722, wire_8275, wire_1806, wire_11829, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11720, wire_8273, wire_1766, wire_11831, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11718, wire_8271, wire_1766, wire_11833, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11716, wire_8269, wire_1766, wire_11835, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11714, wire_8267, wire_1810, wire_1766, wire_11837, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11712, wire_8265, wire_1810, wire_1766, wire_11839, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11710, wire_8263, wire_1810, wire_1766, wire_11841, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11708, wire_8261, wire_1810, wire_1762, wire_11843, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11706, wire_8259, wire_1810, wire_1762, wire_11845, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11704, wire_8257, wire_1810, wire_1762, wire_11847, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11702, wire_8255, wire_1806, wire_1762, wire_11849, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11700, wire_8253, wire_1806, wire_1762, wire_11821, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11728, wire_8251, wire_1806, wire_1762};
    // CHNAXY TOTAL: 636
    assign wire_8071 = lut_tile_5_3_chanxy_out[0];
    assign wire_8079 = lut_tile_5_3_chanxy_out[1];
    assign wire_8087 = lut_tile_5_3_chanxy_out[2];
    assign wire_8095 = lut_tile_5_3_chanxy_out[3];
    assign wire_8103 = lut_tile_5_3_chanxy_out[4];
    assign wire_8111 = lut_tile_5_3_chanxy_out[5];
    assign wire_8119 = lut_tile_5_3_chanxy_out[6];
    assign wire_8127 = lut_tile_5_3_chanxy_out[7];
    assign wire_8135 = lut_tile_5_3_chanxy_out[8];
    assign wire_8143 = lut_tile_5_3_chanxy_out[9];
    assign wire_8151 = lut_tile_5_3_chanxy_out[10];
    assign wire_8159 = lut_tile_5_3_chanxy_out[11];
    assign wire_8167 = lut_tile_5_3_chanxy_out[12];
    assign wire_8175 = lut_tile_5_3_chanxy_out[13];
    assign wire_8183 = lut_tile_5_3_chanxy_out[14];
    assign wire_8220 = lut_tile_5_3_chanxy_out[15];
    assign wire_8222 = lut_tile_5_3_chanxy_out[16];
    assign wire_8224 = lut_tile_5_3_chanxy_out[17];
    assign wire_8226 = lut_tile_5_3_chanxy_out[18];
    assign wire_8228 = lut_tile_5_3_chanxy_out[19];
    assign wire_8230 = lut_tile_5_3_chanxy_out[20];
    assign wire_8232 = lut_tile_5_3_chanxy_out[21];
    assign wire_8234 = lut_tile_5_3_chanxy_out[22];
    assign wire_8236 = lut_tile_5_3_chanxy_out[23];
    assign wire_8238 = lut_tile_5_3_chanxy_out[24];
    assign wire_8240 = lut_tile_5_3_chanxy_out[25];
    assign wire_8242 = lut_tile_5_3_chanxy_out[26];
    assign wire_8244 = lut_tile_5_3_chanxy_out[27];
    assign wire_8246 = lut_tile_5_3_chanxy_out[28];
    assign wire_8248 = lut_tile_5_3_chanxy_out[29];
    assign wire_11701 = lut_tile_5_3_chanxy_out[30];
    assign wire_11703 = lut_tile_5_3_chanxy_out[31];
    assign wire_11705 = lut_tile_5_3_chanxy_out[32];
    assign wire_11707 = lut_tile_5_3_chanxy_out[33];
    assign wire_11709 = lut_tile_5_3_chanxy_out[34];
    assign wire_11711 = lut_tile_5_3_chanxy_out[35];
    assign wire_11713 = lut_tile_5_3_chanxy_out[36];
    assign wire_11715 = lut_tile_5_3_chanxy_out[37];
    assign wire_11717 = lut_tile_5_3_chanxy_out[38];
    assign wire_11719 = lut_tile_5_3_chanxy_out[39];
    assign wire_11721 = lut_tile_5_3_chanxy_out[40];
    assign wire_11723 = lut_tile_5_3_chanxy_out[41];
    assign wire_11725 = lut_tile_5_3_chanxy_out[42];
    assign wire_11727 = lut_tile_5_3_chanxy_out[43];
    assign wire_11729 = lut_tile_5_3_chanxy_out[44];
    assign wire_11790 = lut_tile_5_3_chanxy_out[45];
    assign wire_11792 = lut_tile_5_3_chanxy_out[46];
    assign wire_11794 = lut_tile_5_3_chanxy_out[47];
    assign wire_11796 = lut_tile_5_3_chanxy_out[48];
    assign wire_11798 = lut_tile_5_3_chanxy_out[49];
    assign wire_11800 = lut_tile_5_3_chanxy_out[50];
    assign wire_11802 = lut_tile_5_3_chanxy_out[51];
    assign wire_11804 = lut_tile_5_3_chanxy_out[52];
    assign wire_11806 = lut_tile_5_3_chanxy_out[53];
    assign wire_11808 = lut_tile_5_3_chanxy_out[54];
    assign wire_11810 = lut_tile_5_3_chanxy_out[55];
    assign wire_11812 = lut_tile_5_3_chanxy_out[56];
    assign wire_11814 = lut_tile_5_3_chanxy_out[57];
    assign wire_11816 = lut_tile_5_3_chanxy_out[58];
    assign wire_11818 = lut_tile_5_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_4_chanxy_in = {wire_12082, wire_7891, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7688, wire_2793, wire_12074, wire_7919, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7696, wire_2793, wire_12066, wire_7917, wire_7829, wire_7828, wire_7819, wire_7818, wire_7809, wire_7808, wire_7704, wire_2793, wire_12058, wire_7915, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7712, wire_2283, wire_12050, wire_7913, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7720, wire_2283, wire_12042, wire_7911, wire_7827, wire_7826, wire_7817, wire_7816, wire_7807, wire_7806, wire_7728, wire_2283, wire_12034, wire_7909, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7736, wire_2797, wire_2283, wire_12026, wire_7907, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7744, wire_2797, wire_2283, wire_12018, wire_7905, wire_7825, wire_7824, wire_7815, wire_7814, wire_7805, wire_7804, wire_7752, wire_2797, wire_2283, wire_12010, wire_7903, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7760, wire_2797, wire_2279, wire_12002, wire_7901, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7768, wire_2797, wire_2279, wire_11994, wire_7899, wire_7823, wire_7822, wire_7813, wire_7812, wire_7803, wire_7802, wire_7776, wire_2797, wire_2279, wire_11986, wire_7897, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7784, wire_2793, wire_2279, wire_11978, wire_7895, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7792, wire_2793, wire_2279, wire_11970, wire_7893, wire_7821, wire_7820, wire_7811, wire_7810, wire_7801, wire_7800, wire_7680, wire_2793, wire_2279, wire_12239, wire_8309, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8072, wire_2793, wire_12237, wire_8281, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8184, wire_2793, wire_12235, wire_8283, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8176, wire_2793, wire_12233, wire_8285, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8168, wire_2283, wire_12231, wire_8287, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8160, wire_2283, wire_12229, wire_8289, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8152, wire_2283, wire_12227, wire_8291, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8144, wire_2797, wire_2283, wire_12225, wire_8293, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8136, wire_2797, wire_2283, wire_12223, wire_8295, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8128, wire_2797, wire_2283, wire_12221, wire_8297, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8120, wire_2797, wire_2279, wire_12219, wire_8299, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8112, wire_2797, wire_2279, wire_12217, wire_8301, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8104, wire_2797, wire_2279, wire_12215, wire_8303, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8096, wire_2793, wire_2279, wire_12213, wire_8305, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8088, wire_2793, wire_2279, wire_12211, wire_8307, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8080, wire_2793, wire_2279, wire_11847, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11728, wire_8182, wire_2322, wire_11845, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11700, wire_8174, wire_2322, wire_11843, wire_11759, wire_11758, wire_11749, wire_11748, wire_11739, wire_11738, wire_11702, wire_8166, wire_2322, wire_11841, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11704, wire_8158, wire_2282, wire_11839, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11706, wire_8150, wire_2282, wire_11837, wire_11757, wire_11756, wire_11747, wire_11746, wire_11737, wire_11736, wire_11708, wire_8142, wire_2282, wire_11835, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11710, wire_8134, wire_2326, wire_2282, wire_11833, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11712, wire_8126, wire_2326, wire_2282, wire_11831, wire_11755, wire_11754, wire_11745, wire_11744, wire_11735, wire_11734, wire_11714, wire_8118, wire_2326, wire_2282, wire_11829, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11716, wire_8110, wire_2326, wire_2278, wire_11827, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11718, wire_8102, wire_2326, wire_2278, wire_11825, wire_11753, wire_11752, wire_11743, wire_11742, wire_11733, wire_11732, wire_11720, wire_8094, wire_2326, wire_2278, wire_11823, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11722, wire_8086, wire_2322, wire_2278, wire_11821, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11724, wire_8078, wire_2322, wire_2278, wire_11849, wire_11751, wire_11750, wire_11741, wire_11740, wire_11731, wire_11730, wire_11726, wire_8070, wire_2322, wire_2278, wire_12213, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12116, wire_8309, wire_2322, wire_12215, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12114, wire_8307, wire_2322, wire_12217, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12112, wire_8305, wire_2322, wire_12219, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12110, wire_8303, wire_2282, wire_12221, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12108, wire_8301, wire_2282, wire_12223, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12106, wire_8299, wire_2282, wire_12225, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12104, wire_8297, wire_2326, wire_2282, wire_12227, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12102, wire_8295, wire_2326, wire_2282, wire_12229, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12100, wire_8293, wire_2326, wire_2282, wire_12231, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12098, wire_8291, wire_2326, wire_2278, wire_12233, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12096, wire_8289, wire_2326, wire_2278, wire_12235, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12094, wire_8287, wire_2326, wire_2278, wire_12237, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12092, wire_8285, wire_2322, wire_2278, wire_12239, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12090, wire_8283, wire_2322, wire_2278, wire_12211, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12118, wire_8281, wire_2322, wire_2278};
    // CHNAXY TOTAL: 636
    assign wire_8073 = lut_tile_5_4_chanxy_out[0];
    assign wire_8081 = lut_tile_5_4_chanxy_out[1];
    assign wire_8089 = lut_tile_5_4_chanxy_out[2];
    assign wire_8097 = lut_tile_5_4_chanxy_out[3];
    assign wire_8105 = lut_tile_5_4_chanxy_out[4];
    assign wire_8113 = lut_tile_5_4_chanxy_out[5];
    assign wire_8121 = lut_tile_5_4_chanxy_out[6];
    assign wire_8129 = lut_tile_5_4_chanxy_out[7];
    assign wire_8137 = lut_tile_5_4_chanxy_out[8];
    assign wire_8145 = lut_tile_5_4_chanxy_out[9];
    assign wire_8153 = lut_tile_5_4_chanxy_out[10];
    assign wire_8161 = lut_tile_5_4_chanxy_out[11];
    assign wire_8169 = lut_tile_5_4_chanxy_out[12];
    assign wire_8177 = lut_tile_5_4_chanxy_out[13];
    assign wire_8185 = lut_tile_5_4_chanxy_out[14];
    assign wire_8250 = lut_tile_5_4_chanxy_out[15];
    assign wire_8252 = lut_tile_5_4_chanxy_out[16];
    assign wire_8254 = lut_tile_5_4_chanxy_out[17];
    assign wire_8256 = lut_tile_5_4_chanxy_out[18];
    assign wire_8258 = lut_tile_5_4_chanxy_out[19];
    assign wire_8260 = lut_tile_5_4_chanxy_out[20];
    assign wire_8262 = lut_tile_5_4_chanxy_out[21];
    assign wire_8264 = lut_tile_5_4_chanxy_out[22];
    assign wire_8266 = lut_tile_5_4_chanxy_out[23];
    assign wire_8268 = lut_tile_5_4_chanxy_out[24];
    assign wire_8270 = lut_tile_5_4_chanxy_out[25];
    assign wire_8272 = lut_tile_5_4_chanxy_out[26];
    assign wire_8274 = lut_tile_5_4_chanxy_out[27];
    assign wire_8276 = lut_tile_5_4_chanxy_out[28];
    assign wire_8278 = lut_tile_5_4_chanxy_out[29];
    assign wire_12091 = lut_tile_5_4_chanxy_out[30];
    assign wire_12093 = lut_tile_5_4_chanxy_out[31];
    assign wire_12095 = lut_tile_5_4_chanxy_out[32];
    assign wire_12097 = lut_tile_5_4_chanxy_out[33];
    assign wire_12099 = lut_tile_5_4_chanxy_out[34];
    assign wire_12101 = lut_tile_5_4_chanxy_out[35];
    assign wire_12103 = lut_tile_5_4_chanxy_out[36];
    assign wire_12105 = lut_tile_5_4_chanxy_out[37];
    assign wire_12107 = lut_tile_5_4_chanxy_out[38];
    assign wire_12109 = lut_tile_5_4_chanxy_out[39];
    assign wire_12111 = lut_tile_5_4_chanxy_out[40];
    assign wire_12113 = lut_tile_5_4_chanxy_out[41];
    assign wire_12115 = lut_tile_5_4_chanxy_out[42];
    assign wire_12117 = lut_tile_5_4_chanxy_out[43];
    assign wire_12119 = lut_tile_5_4_chanxy_out[44];
    assign wire_12180 = lut_tile_5_4_chanxy_out[45];
    assign wire_12182 = lut_tile_5_4_chanxy_out[46];
    assign wire_12184 = lut_tile_5_4_chanxy_out[47];
    assign wire_12186 = lut_tile_5_4_chanxy_out[48];
    assign wire_12188 = lut_tile_5_4_chanxy_out[49];
    assign wire_12190 = lut_tile_5_4_chanxy_out[50];
    assign wire_12192 = lut_tile_5_4_chanxy_out[51];
    assign wire_12194 = lut_tile_5_4_chanxy_out[52];
    assign wire_12196 = lut_tile_5_4_chanxy_out[53];
    assign wire_12198 = lut_tile_5_4_chanxy_out[54];
    assign wire_12200 = lut_tile_5_4_chanxy_out[55];
    assign wire_12202 = lut_tile_5_4_chanxy_out[56];
    assign wire_12204 = lut_tile_5_4_chanxy_out[57];
    assign wire_12206 = lut_tile_5_4_chanxy_out[58];
    assign wire_12208 = lut_tile_5_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_5_chanxy_in = {wire_12474, wire_7921, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7802, wire_3309, wire_12466, wire_7949, wire_7859, wire_7858, wire_7849, wire_7848, wire_7839, wire_7838, wire_7804, wire_3309, wire_12458, wire_7947, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7806, wire_3309, wire_12450, wire_7945, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7808, wire_2799, wire_12442, wire_7943, wire_7857, wire_7856, wire_7847, wire_7846, wire_7837, wire_7836, wire_7810, wire_2799, wire_12434, wire_7941, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7812, wire_2799, wire_12426, wire_7939, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7814, wire_3313, wire_2799, wire_12418, wire_7937, wire_7855, wire_7854, wire_7845, wire_7844, wire_7835, wire_7834, wire_7816, wire_3313, wire_2799, wire_12410, wire_7935, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7818, wire_3313, wire_2799, wire_12402, wire_7933, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7820, wire_3313, wire_2795, wire_12394, wire_7931, wire_7853, wire_7852, wire_7843, wire_7842, wire_7833, wire_7832, wire_7822, wire_3313, wire_2795, wire_12386, wire_7929, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7824, wire_3313, wire_2795, wire_12378, wire_7927, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7826, wire_3309, wire_2795, wire_12370, wire_7925, wire_7851, wire_7850, wire_7841, wire_7840, wire_7831, wire_7830, wire_7828, wire_3309, wire_2795, wire_12362, wire_7923, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7800, wire_3309, wire_2795, wire_12629, wire_8339, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8190, wire_3309, wire_12627, wire_8311, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8218, wire_3309, wire_12625, wire_8313, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8216, wire_3309, wire_12623, wire_8315, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8214, wire_2799, wire_12621, wire_8317, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8212, wire_2799, wire_12619, wire_8319, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8210, wire_2799, wire_12617, wire_8321, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8208, wire_3313, wire_2799, wire_12615, wire_8323, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8206, wire_3313, wire_2799, wire_12613, wire_8325, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8204, wire_3313, wire_2799, wire_12611, wire_8327, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8202, wire_3313, wire_2795, wire_12609, wire_8329, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8200, wire_3313, wire_2795, wire_12607, wire_8331, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8198, wire_3313, wire_2795, wire_12605, wire_8333, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8196, wire_3309, wire_2795, wire_12603, wire_8335, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8194, wire_3309, wire_2795, wire_12601, wire_8337, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8192, wire_3309, wire_2795, wire_12237, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12118, wire_8184, wire_2838, wire_12235, wire_12149, wire_12148, wire_12139, wire_12138, wire_12129, wire_12128, wire_12090, wire_8176, wire_2838, wire_12233, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12092, wire_8168, wire_2838, wire_12231, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12094, wire_8160, wire_2798, wire_12229, wire_12147, wire_12146, wire_12137, wire_12136, wire_12127, wire_12126, wire_12096, wire_8152, wire_2798, wire_12227, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12098, wire_8144, wire_2798, wire_12225, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12100, wire_8136, wire_2842, wire_2798, wire_12223, wire_12145, wire_12144, wire_12135, wire_12134, wire_12125, wire_12124, wire_12102, wire_8128, wire_2842, wire_2798, wire_12221, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12104, wire_8120, wire_2842, wire_2798, wire_12219, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12106, wire_8112, wire_2842, wire_2794, wire_12217, wire_12143, wire_12142, wire_12133, wire_12132, wire_12123, wire_12122, wire_12108, wire_8104, wire_2842, wire_2794, wire_12215, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12110, wire_8096, wire_2842, wire_2794, wire_12213, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12112, wire_8088, wire_2838, wire_2794, wire_12211, wire_12141, wire_12140, wire_12131, wire_12130, wire_12121, wire_12120, wire_12114, wire_8080, wire_2838, wire_2794, wire_12239, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12116, wire_8072, wire_2838, wire_2794, wire_12603, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12506, wire_8339, wire_2838, wire_12605, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12504, wire_8337, wire_2838, wire_12607, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12502, wire_8335, wire_2838, wire_12609, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12500, wire_8333, wire_2798, wire_12611, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12498, wire_8331, wire_2798, wire_12613, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12496, wire_8329, wire_2798, wire_12615, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12494, wire_8327, wire_2842, wire_2798, wire_12617, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12492, wire_8325, wire_2842, wire_2798, wire_12619, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12490, wire_8323, wire_2842, wire_2798, wire_12621, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12488, wire_8321, wire_2842, wire_2794, wire_12623, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12486, wire_8319, wire_2842, wire_2794, wire_12625, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12484, wire_8317, wire_2842, wire_2794, wire_12627, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12482, wire_8315, wire_2838, wire_2794, wire_12629, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12480, wire_8313, wire_2838, wire_2794, wire_12601, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12508, wire_8311, wire_2838, wire_2794};
    // CHNAXY TOTAL: 636
    assign wire_8191 = lut_tile_5_5_chanxy_out[0];
    assign wire_8193 = lut_tile_5_5_chanxy_out[1];
    assign wire_8195 = lut_tile_5_5_chanxy_out[2];
    assign wire_8197 = lut_tile_5_5_chanxy_out[3];
    assign wire_8199 = lut_tile_5_5_chanxy_out[4];
    assign wire_8201 = lut_tile_5_5_chanxy_out[5];
    assign wire_8203 = lut_tile_5_5_chanxy_out[6];
    assign wire_8205 = lut_tile_5_5_chanxy_out[7];
    assign wire_8207 = lut_tile_5_5_chanxy_out[8];
    assign wire_8209 = lut_tile_5_5_chanxy_out[9];
    assign wire_8211 = lut_tile_5_5_chanxy_out[10];
    assign wire_8213 = lut_tile_5_5_chanxy_out[11];
    assign wire_8215 = lut_tile_5_5_chanxy_out[12];
    assign wire_8217 = lut_tile_5_5_chanxy_out[13];
    assign wire_8219 = lut_tile_5_5_chanxy_out[14];
    assign wire_8280 = lut_tile_5_5_chanxy_out[15];
    assign wire_8282 = lut_tile_5_5_chanxy_out[16];
    assign wire_8284 = lut_tile_5_5_chanxy_out[17];
    assign wire_8286 = lut_tile_5_5_chanxy_out[18];
    assign wire_8288 = lut_tile_5_5_chanxy_out[19];
    assign wire_8290 = lut_tile_5_5_chanxy_out[20];
    assign wire_8292 = lut_tile_5_5_chanxy_out[21];
    assign wire_8294 = lut_tile_5_5_chanxy_out[22];
    assign wire_8296 = lut_tile_5_5_chanxy_out[23];
    assign wire_8298 = lut_tile_5_5_chanxy_out[24];
    assign wire_8300 = lut_tile_5_5_chanxy_out[25];
    assign wire_8302 = lut_tile_5_5_chanxy_out[26];
    assign wire_8304 = lut_tile_5_5_chanxy_out[27];
    assign wire_8306 = lut_tile_5_5_chanxy_out[28];
    assign wire_8308 = lut_tile_5_5_chanxy_out[29];
    assign wire_12481 = lut_tile_5_5_chanxy_out[30];
    assign wire_12483 = lut_tile_5_5_chanxy_out[31];
    assign wire_12485 = lut_tile_5_5_chanxy_out[32];
    assign wire_12487 = lut_tile_5_5_chanxy_out[33];
    assign wire_12489 = lut_tile_5_5_chanxy_out[34];
    assign wire_12491 = lut_tile_5_5_chanxy_out[35];
    assign wire_12493 = lut_tile_5_5_chanxy_out[36];
    assign wire_12495 = lut_tile_5_5_chanxy_out[37];
    assign wire_12497 = lut_tile_5_5_chanxy_out[38];
    assign wire_12499 = lut_tile_5_5_chanxy_out[39];
    assign wire_12501 = lut_tile_5_5_chanxy_out[40];
    assign wire_12503 = lut_tile_5_5_chanxy_out[41];
    assign wire_12505 = lut_tile_5_5_chanxy_out[42];
    assign wire_12507 = lut_tile_5_5_chanxy_out[43];
    assign wire_12509 = lut_tile_5_5_chanxy_out[44];
    assign wire_12570 = lut_tile_5_5_chanxy_out[45];
    assign wire_12572 = lut_tile_5_5_chanxy_out[46];
    assign wire_12574 = lut_tile_5_5_chanxy_out[47];
    assign wire_12576 = lut_tile_5_5_chanxy_out[48];
    assign wire_12578 = lut_tile_5_5_chanxy_out[49];
    assign wire_12580 = lut_tile_5_5_chanxy_out[50];
    assign wire_12582 = lut_tile_5_5_chanxy_out[51];
    assign wire_12584 = lut_tile_5_5_chanxy_out[52];
    assign wire_12586 = lut_tile_5_5_chanxy_out[53];
    assign wire_12588 = lut_tile_5_5_chanxy_out[54];
    assign wire_12590 = lut_tile_5_5_chanxy_out[55];
    assign wire_12592 = lut_tile_5_5_chanxy_out[56];
    assign wire_12594 = lut_tile_5_5_chanxy_out[57];
    assign wire_12596 = lut_tile_5_5_chanxy_out[58];
    assign wire_12598 = lut_tile_5_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_6_chanxy_in = {wire_12866, wire_7951, wire_7889, wire_7888, wire_7879, wire_7878, wire_7869, wire_7868, wire_7832, wire_3825, wire_12858, wire_7979, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7834, wire_3825, wire_12850, wire_7977, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7836, wire_3825, wire_12842, wire_7975, wire_7887, wire_7886, wire_7877, wire_7876, wire_7867, wire_7866, wire_7838, wire_3315, wire_12834, wire_7973, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7840, wire_3315, wire_12826, wire_7971, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7842, wire_3315, wire_12818, wire_7969, wire_7885, wire_7884, wire_7875, wire_7874, wire_7865, wire_7864, wire_7844, wire_3829, wire_3315, wire_12810, wire_7967, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7846, wire_3829, wire_3315, wire_12802, wire_7965, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7848, wire_3829, wire_3315, wire_12794, wire_7963, wire_7883, wire_7882, wire_7873, wire_7872, wire_7863, wire_7862, wire_7850, wire_3829, wire_3311, wire_12786, wire_7961, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7852, wire_3829, wire_3311, wire_12778, wire_7959, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7854, wire_3829, wire_3311, wire_12770, wire_7957, wire_7881, wire_7880, wire_7871, wire_7870, wire_7861, wire_7860, wire_7856, wire_3825, wire_3311, wire_12762, wire_7955, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7858, wire_3825, wire_3311, wire_12754, wire_7953, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7830, wire_3825, wire_3311, wire_13019, wire_8369, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8220, wire_3825, wire_13017, wire_8341, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8248, wire_3825, wire_13015, wire_8343, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8246, wire_3825, wire_13013, wire_8345, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8244, wire_3315, wire_13011, wire_8347, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8242, wire_3315, wire_13009, wire_8349, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8240, wire_3315, wire_13007, wire_8351, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8238, wire_3829, wire_3315, wire_13005, wire_8353, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8236, wire_3829, wire_3315, wire_13003, wire_8355, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8234, wire_3829, wire_3315, wire_13001, wire_8357, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8232, wire_3829, wire_3311, wire_12999, wire_8359, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8230, wire_3829, wire_3311, wire_12997, wire_8361, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8228, wire_3829, wire_3311, wire_12995, wire_8363, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8226, wire_3825, wire_3311, wire_12993, wire_8365, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8224, wire_3825, wire_3311, wire_12991, wire_8367, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8222, wire_3825, wire_3311, wire_12627, wire_12539, wire_12538, wire_12529, wire_12528, wire_12519, wire_12518, wire_12508, wire_8218, wire_3354, wire_12625, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12480, wire_8216, wire_3354, wire_12623, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12482, wire_8214, wire_3354, wire_12621, wire_12537, wire_12536, wire_12527, wire_12526, wire_12517, wire_12516, wire_12484, wire_8212, wire_3314, wire_12619, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12486, wire_8210, wire_3314, wire_12617, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12488, wire_8208, wire_3314, wire_12615, wire_12535, wire_12534, wire_12525, wire_12524, wire_12515, wire_12514, wire_12490, wire_8206, wire_3358, wire_3314, wire_12613, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12492, wire_8204, wire_3358, wire_3314, wire_12611, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12494, wire_8202, wire_3358, wire_3314, wire_12609, wire_12533, wire_12532, wire_12523, wire_12522, wire_12513, wire_12512, wire_12496, wire_8200, wire_3358, wire_3310, wire_12607, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12498, wire_8198, wire_3358, wire_3310, wire_12605, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12500, wire_8196, wire_3358, wire_3310, wire_12603, wire_12531, wire_12530, wire_12521, wire_12520, wire_12511, wire_12510, wire_12502, wire_8194, wire_3354, wire_3310, wire_12601, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12504, wire_8192, wire_3354, wire_3310, wire_12629, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12506, wire_8190, wire_3354, wire_3310, wire_12993, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12896, wire_8369, wire_3354, wire_12995, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12894, wire_8367, wire_3354, wire_12997, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12892, wire_8365, wire_3354, wire_12999, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12890, wire_8363, wire_3314, wire_13001, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12888, wire_8361, wire_3314, wire_13003, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12886, wire_8359, wire_3314, wire_13005, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12884, wire_8357, wire_3358, wire_3314, wire_13007, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12882, wire_8355, wire_3358, wire_3314, wire_13009, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12880, wire_8353, wire_3358, wire_3314, wire_13011, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12878, wire_8351, wire_3358, wire_3310, wire_13013, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12876, wire_8349, wire_3358, wire_3310, wire_13015, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12874, wire_8347, wire_3358, wire_3310, wire_13017, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12872, wire_8345, wire_3354, wire_3310, wire_13019, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12870, wire_8343, wire_3354, wire_3310, wire_12991, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12898, wire_8341, wire_3354, wire_3310};
    // CHNAXY TOTAL: 636
    assign wire_8221 = lut_tile_5_6_chanxy_out[0];
    assign wire_8223 = lut_tile_5_6_chanxy_out[1];
    assign wire_8225 = lut_tile_5_6_chanxy_out[2];
    assign wire_8227 = lut_tile_5_6_chanxy_out[3];
    assign wire_8229 = lut_tile_5_6_chanxy_out[4];
    assign wire_8231 = lut_tile_5_6_chanxy_out[5];
    assign wire_8233 = lut_tile_5_6_chanxy_out[6];
    assign wire_8235 = lut_tile_5_6_chanxy_out[7];
    assign wire_8237 = lut_tile_5_6_chanxy_out[8];
    assign wire_8239 = lut_tile_5_6_chanxy_out[9];
    assign wire_8241 = lut_tile_5_6_chanxy_out[10];
    assign wire_8243 = lut_tile_5_6_chanxy_out[11];
    assign wire_8245 = lut_tile_5_6_chanxy_out[12];
    assign wire_8247 = lut_tile_5_6_chanxy_out[13];
    assign wire_8249 = lut_tile_5_6_chanxy_out[14];
    assign wire_8310 = lut_tile_5_6_chanxy_out[15];
    assign wire_8312 = lut_tile_5_6_chanxy_out[16];
    assign wire_8314 = lut_tile_5_6_chanxy_out[17];
    assign wire_8316 = lut_tile_5_6_chanxy_out[18];
    assign wire_8318 = lut_tile_5_6_chanxy_out[19];
    assign wire_8320 = lut_tile_5_6_chanxy_out[20];
    assign wire_8322 = lut_tile_5_6_chanxy_out[21];
    assign wire_8324 = lut_tile_5_6_chanxy_out[22];
    assign wire_8326 = lut_tile_5_6_chanxy_out[23];
    assign wire_8328 = lut_tile_5_6_chanxy_out[24];
    assign wire_8330 = lut_tile_5_6_chanxy_out[25];
    assign wire_8332 = lut_tile_5_6_chanxy_out[26];
    assign wire_8334 = lut_tile_5_6_chanxy_out[27];
    assign wire_8336 = lut_tile_5_6_chanxy_out[28];
    assign wire_8338 = lut_tile_5_6_chanxy_out[29];
    assign wire_12871 = lut_tile_5_6_chanxy_out[30];
    assign wire_12873 = lut_tile_5_6_chanxy_out[31];
    assign wire_12875 = lut_tile_5_6_chanxy_out[32];
    assign wire_12877 = lut_tile_5_6_chanxy_out[33];
    assign wire_12879 = lut_tile_5_6_chanxy_out[34];
    assign wire_12881 = lut_tile_5_6_chanxy_out[35];
    assign wire_12883 = lut_tile_5_6_chanxy_out[36];
    assign wire_12885 = lut_tile_5_6_chanxy_out[37];
    assign wire_12887 = lut_tile_5_6_chanxy_out[38];
    assign wire_12889 = lut_tile_5_6_chanxy_out[39];
    assign wire_12891 = lut_tile_5_6_chanxy_out[40];
    assign wire_12893 = lut_tile_5_6_chanxy_out[41];
    assign wire_12895 = lut_tile_5_6_chanxy_out[42];
    assign wire_12897 = lut_tile_5_6_chanxy_out[43];
    assign wire_12899 = lut_tile_5_6_chanxy_out[44];
    assign wire_12960 = lut_tile_5_6_chanxy_out[45];
    assign wire_12962 = lut_tile_5_6_chanxy_out[46];
    assign wire_12964 = lut_tile_5_6_chanxy_out[47];
    assign wire_12966 = lut_tile_5_6_chanxy_out[48];
    assign wire_12968 = lut_tile_5_6_chanxy_out[49];
    assign wire_12970 = lut_tile_5_6_chanxy_out[50];
    assign wire_12972 = lut_tile_5_6_chanxy_out[51];
    assign wire_12974 = lut_tile_5_6_chanxy_out[52];
    assign wire_12976 = lut_tile_5_6_chanxy_out[53];
    assign wire_12978 = lut_tile_5_6_chanxy_out[54];
    assign wire_12980 = lut_tile_5_6_chanxy_out[55];
    assign wire_12982 = lut_tile_5_6_chanxy_out[56];
    assign wire_12984 = lut_tile_5_6_chanxy_out[57];
    assign wire_12986 = lut_tile_5_6_chanxy_out[58];
    assign wire_12988 = lut_tile_5_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_7_chanxy_in = {wire_13258, wire_7981, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7862, wire_4341, wire_13250, wire_8009, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7864, wire_4341, wire_13242, wire_8007, wire_7919, wire_7918, wire_7909, wire_7908, wire_7899, wire_7898, wire_7866, wire_4341, wire_13234, wire_8005, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7868, wire_3831, wire_13226, wire_8003, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7870, wire_3831, wire_13218, wire_8001, wire_7917, wire_7916, wire_7907, wire_7906, wire_7897, wire_7896, wire_7872, wire_3831, wire_13210, wire_7999, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7874, wire_4345, wire_3831, wire_13202, wire_7997, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7876, wire_4345, wire_3831, wire_13194, wire_7995, wire_7915, wire_7914, wire_7905, wire_7904, wire_7895, wire_7894, wire_7878, wire_4345, wire_3831, wire_13186, wire_7993, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7880, wire_4345, wire_3827, wire_13178, wire_7991, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7882, wire_4345, wire_3827, wire_13170, wire_7989, wire_7913, wire_7912, wire_7903, wire_7902, wire_7893, wire_7892, wire_7884, wire_4345, wire_3827, wire_13162, wire_7987, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7886, wire_4341, wire_3827, wire_13154, wire_7985, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7888, wire_4341, wire_3827, wire_13146, wire_7983, wire_7911, wire_7910, wire_7901, wire_7900, wire_7891, wire_7890, wire_7860, wire_4341, wire_3827, wire_13409, wire_8399, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8250, wire_4341, wire_13407, wire_8371, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8278, wire_4341, wire_13405, wire_8373, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8276, wire_4341, wire_13403, wire_8375, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8274, wire_3831, wire_13401, wire_8377, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8272, wire_3831, wire_13399, wire_8379, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8270, wire_3831, wire_13397, wire_8381, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8268, wire_4345, wire_3831, wire_13395, wire_8383, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8266, wire_4345, wire_3831, wire_13393, wire_8385, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8264, wire_4345, wire_3831, wire_13391, wire_8387, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8262, wire_4345, wire_3827, wire_13389, wire_8389, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8260, wire_4345, wire_3827, wire_13387, wire_8391, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8258, wire_4345, wire_3827, wire_13385, wire_8393, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8256, wire_4341, wire_3827, wire_13383, wire_8395, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8254, wire_4341, wire_3827, wire_13381, wire_8397, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8252, wire_4341, wire_3827, wire_13017, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12898, wire_8248, wire_3870, wire_13015, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12870, wire_8246, wire_3870, wire_13013, wire_12929, wire_12928, wire_12919, wire_12918, wire_12909, wire_12908, wire_12872, wire_8244, wire_3870, wire_13011, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12874, wire_8242, wire_3830, wire_13009, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12876, wire_8240, wire_3830, wire_13007, wire_12927, wire_12926, wire_12917, wire_12916, wire_12907, wire_12906, wire_12878, wire_8238, wire_3830, wire_13005, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12880, wire_8236, wire_3874, wire_3830, wire_13003, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12882, wire_8234, wire_3874, wire_3830, wire_13001, wire_12925, wire_12924, wire_12915, wire_12914, wire_12905, wire_12904, wire_12884, wire_8232, wire_3874, wire_3830, wire_12999, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12886, wire_8230, wire_3874, wire_3826, wire_12997, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12888, wire_8228, wire_3874, wire_3826, wire_12995, wire_12923, wire_12922, wire_12913, wire_12912, wire_12903, wire_12902, wire_12890, wire_8226, wire_3874, wire_3826, wire_12993, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12892, wire_8224, wire_3870, wire_3826, wire_12991, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12894, wire_8222, wire_3870, wire_3826, wire_13019, wire_12921, wire_12920, wire_12911, wire_12910, wire_12901, wire_12900, wire_12896, wire_8220, wire_3870, wire_3826, wire_13383, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13286, wire_8399, wire_3870, wire_13385, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13284, wire_8397, wire_3870, wire_13387, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13282, wire_8395, wire_3870, wire_13389, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13280, wire_8393, wire_3830, wire_13391, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13278, wire_8391, wire_3830, wire_13393, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13276, wire_8389, wire_3830, wire_13395, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13274, wire_8387, wire_3874, wire_3830, wire_13397, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13272, wire_8385, wire_3874, wire_3830, wire_13399, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13270, wire_8383, wire_3874, wire_3830, wire_13401, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13268, wire_8381, wire_3874, wire_3826, wire_13403, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13266, wire_8379, wire_3874, wire_3826, wire_13405, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13264, wire_8377, wire_3874, wire_3826, wire_13407, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13262, wire_8375, wire_3870, wire_3826, wire_13409, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13260, wire_8373, wire_3870, wire_3826, wire_13381, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13288, wire_8371, wire_3870, wire_3826};
    // CHNAXY TOTAL: 636
    assign wire_8251 = lut_tile_5_7_chanxy_out[0];
    assign wire_8253 = lut_tile_5_7_chanxy_out[1];
    assign wire_8255 = lut_tile_5_7_chanxy_out[2];
    assign wire_8257 = lut_tile_5_7_chanxy_out[3];
    assign wire_8259 = lut_tile_5_7_chanxy_out[4];
    assign wire_8261 = lut_tile_5_7_chanxy_out[5];
    assign wire_8263 = lut_tile_5_7_chanxy_out[6];
    assign wire_8265 = lut_tile_5_7_chanxy_out[7];
    assign wire_8267 = lut_tile_5_7_chanxy_out[8];
    assign wire_8269 = lut_tile_5_7_chanxy_out[9];
    assign wire_8271 = lut_tile_5_7_chanxy_out[10];
    assign wire_8273 = lut_tile_5_7_chanxy_out[11];
    assign wire_8275 = lut_tile_5_7_chanxy_out[12];
    assign wire_8277 = lut_tile_5_7_chanxy_out[13];
    assign wire_8279 = lut_tile_5_7_chanxy_out[14];
    assign wire_8340 = lut_tile_5_7_chanxy_out[15];
    assign wire_8342 = lut_tile_5_7_chanxy_out[16];
    assign wire_8344 = lut_tile_5_7_chanxy_out[17];
    assign wire_8346 = lut_tile_5_7_chanxy_out[18];
    assign wire_8348 = lut_tile_5_7_chanxy_out[19];
    assign wire_8350 = lut_tile_5_7_chanxy_out[20];
    assign wire_8352 = lut_tile_5_7_chanxy_out[21];
    assign wire_8354 = lut_tile_5_7_chanxy_out[22];
    assign wire_8356 = lut_tile_5_7_chanxy_out[23];
    assign wire_8358 = lut_tile_5_7_chanxy_out[24];
    assign wire_8360 = lut_tile_5_7_chanxy_out[25];
    assign wire_8362 = lut_tile_5_7_chanxy_out[26];
    assign wire_8364 = lut_tile_5_7_chanxy_out[27];
    assign wire_8366 = lut_tile_5_7_chanxy_out[28];
    assign wire_8368 = lut_tile_5_7_chanxy_out[29];
    assign wire_13261 = lut_tile_5_7_chanxy_out[30];
    assign wire_13263 = lut_tile_5_7_chanxy_out[31];
    assign wire_13265 = lut_tile_5_7_chanxy_out[32];
    assign wire_13267 = lut_tile_5_7_chanxy_out[33];
    assign wire_13269 = lut_tile_5_7_chanxy_out[34];
    assign wire_13271 = lut_tile_5_7_chanxy_out[35];
    assign wire_13273 = lut_tile_5_7_chanxy_out[36];
    assign wire_13275 = lut_tile_5_7_chanxy_out[37];
    assign wire_13277 = lut_tile_5_7_chanxy_out[38];
    assign wire_13279 = lut_tile_5_7_chanxy_out[39];
    assign wire_13281 = lut_tile_5_7_chanxy_out[40];
    assign wire_13283 = lut_tile_5_7_chanxy_out[41];
    assign wire_13285 = lut_tile_5_7_chanxy_out[42];
    assign wire_13287 = lut_tile_5_7_chanxy_out[43];
    assign wire_13289 = lut_tile_5_7_chanxy_out[44];
    assign wire_13350 = lut_tile_5_7_chanxy_out[45];
    assign wire_13352 = lut_tile_5_7_chanxy_out[46];
    assign wire_13354 = lut_tile_5_7_chanxy_out[47];
    assign wire_13356 = lut_tile_5_7_chanxy_out[48];
    assign wire_13358 = lut_tile_5_7_chanxy_out[49];
    assign wire_13360 = lut_tile_5_7_chanxy_out[50];
    assign wire_13362 = lut_tile_5_7_chanxy_out[51];
    assign wire_13364 = lut_tile_5_7_chanxy_out[52];
    assign wire_13366 = lut_tile_5_7_chanxy_out[53];
    assign wire_13368 = lut_tile_5_7_chanxy_out[54];
    assign wire_13370 = lut_tile_5_7_chanxy_out[55];
    assign wire_13372 = lut_tile_5_7_chanxy_out[56];
    assign wire_13374 = lut_tile_5_7_chanxy_out[57];
    assign wire_13376 = lut_tile_5_7_chanxy_out[58];
    assign wire_13378 = lut_tile_5_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_8_chanxy_in = {wire_13642, wire_8011, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7892, wire_4857, wire_13634, wire_8039, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7894, wire_4857, wire_13626, wire_8037, wire_7949, wire_7948, wire_7939, wire_7938, wire_7929, wire_7928, wire_7896, wire_4857, wire_13618, wire_8035, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7898, wire_4347, wire_13610, wire_8033, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7900, wire_4347, wire_13602, wire_8031, wire_7947, wire_7946, wire_7937, wire_7936, wire_7927, wire_7926, wire_7902, wire_4347, wire_13594, wire_8029, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7904, wire_4861, wire_4347, wire_13586, wire_8027, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7906, wire_4861, wire_4347, wire_13578, wire_8025, wire_7945, wire_7944, wire_7935, wire_7934, wire_7925, wire_7924, wire_7908, wire_4861, wire_4347, wire_13570, wire_8023, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7910, wire_4861, wire_4343, wire_13562, wire_8021, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7912, wire_4861, wire_4343, wire_13554, wire_8019, wire_7943, wire_7942, wire_7933, wire_7932, wire_7923, wire_7922, wire_7914, wire_4861, wire_4343, wire_13546, wire_8017, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7916, wire_4857, wire_4343, wire_13538, wire_8015, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7918, wire_4857, wire_4343, wire_13530, wire_8013, wire_7941, wire_7940, wire_7931, wire_7930, wire_7921, wire_7920, wire_7890, wire_4857, wire_4343, wire_13799, wire_8429, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8280, wire_4857, wire_13797, wire_8401, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8308, wire_4857, wire_13795, wire_8403, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8306, wire_4857, wire_13793, wire_8405, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8304, wire_4347, wire_13791, wire_8407, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8302, wire_4347, wire_13789, wire_8409, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8300, wire_4347, wire_13787, wire_8411, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8298, wire_4861, wire_4347, wire_13785, wire_8413, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8296, wire_4861, wire_4347, wire_13783, wire_8415, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8294, wire_4861, wire_4347, wire_13781, wire_8417, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8292, wire_4861, wire_4343, wire_13779, wire_8419, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8290, wire_4861, wire_4343, wire_13777, wire_8421, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8288, wire_4861, wire_4343, wire_13775, wire_8423, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8286, wire_4857, wire_4343, wire_13773, wire_8425, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8284, wire_4857, wire_4343, wire_13771, wire_8427, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8282, wire_4857, wire_4343, wire_13407, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13288, wire_8278, wire_4386, wire_13405, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13260, wire_8276, wire_4386, wire_13403, wire_13319, wire_13318, wire_13309, wire_13308, wire_13299, wire_13298, wire_13262, wire_8274, wire_4386, wire_13401, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13264, wire_8272, wire_4346, wire_13399, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13266, wire_8270, wire_4346, wire_13397, wire_13317, wire_13316, wire_13307, wire_13306, wire_13297, wire_13296, wire_13268, wire_8268, wire_4346, wire_13395, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13270, wire_8266, wire_4390, wire_4346, wire_13393, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13272, wire_8264, wire_4390, wire_4346, wire_13391, wire_13315, wire_13314, wire_13305, wire_13304, wire_13295, wire_13294, wire_13274, wire_8262, wire_4390, wire_4346, wire_13389, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13276, wire_8260, wire_4390, wire_4342, wire_13387, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13278, wire_8258, wire_4390, wire_4342, wire_13385, wire_13313, wire_13312, wire_13303, wire_13302, wire_13293, wire_13292, wire_13280, wire_8256, wire_4390, wire_4342, wire_13383, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13282, wire_8254, wire_4386, wire_4342, wire_13381, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13284, wire_8252, wire_4386, wire_4342, wire_13409, wire_13311, wire_13310, wire_13301, wire_13300, wire_13291, wire_13290, wire_13286, wire_8250, wire_4386, wire_4342, wire_13773, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13676, wire_8429, wire_4386, wire_13775, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13674, wire_8427, wire_4386, wire_13777, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13672, wire_8425, wire_4386, wire_13779, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13670, wire_8423, wire_4346, wire_13781, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13668, wire_8421, wire_4346, wire_13783, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13666, wire_8419, wire_4346, wire_13785, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13664, wire_8417, wire_4390, wire_4346, wire_13787, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13662, wire_8415, wire_4390, wire_4346, wire_13789, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13660, wire_8413, wire_4390, wire_4346, wire_13791, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13658, wire_8411, wire_4390, wire_4342, wire_13793, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13656, wire_8409, wire_4390, wire_4342, wire_13795, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13654, wire_8407, wire_4390, wire_4342, wire_13797, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13652, wire_8405, wire_4386, wire_4342, wire_13799, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13650, wire_8403, wire_4386, wire_4342, wire_13771, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13678, wire_8401, wire_4386, wire_4342};
    // CHNAXY TOTAL: 636
    assign wire_8281 = lut_tile_5_8_chanxy_out[0];
    assign wire_8283 = lut_tile_5_8_chanxy_out[1];
    assign wire_8285 = lut_tile_5_8_chanxy_out[2];
    assign wire_8287 = lut_tile_5_8_chanxy_out[3];
    assign wire_8289 = lut_tile_5_8_chanxy_out[4];
    assign wire_8291 = lut_tile_5_8_chanxy_out[5];
    assign wire_8293 = lut_tile_5_8_chanxy_out[6];
    assign wire_8295 = lut_tile_5_8_chanxy_out[7];
    assign wire_8297 = lut_tile_5_8_chanxy_out[8];
    assign wire_8299 = lut_tile_5_8_chanxy_out[9];
    assign wire_8301 = lut_tile_5_8_chanxy_out[10];
    assign wire_8303 = lut_tile_5_8_chanxy_out[11];
    assign wire_8305 = lut_tile_5_8_chanxy_out[12];
    assign wire_8307 = lut_tile_5_8_chanxy_out[13];
    assign wire_8309 = lut_tile_5_8_chanxy_out[14];
    assign wire_8370 = lut_tile_5_8_chanxy_out[15];
    assign wire_8372 = lut_tile_5_8_chanxy_out[16];
    assign wire_8374 = lut_tile_5_8_chanxy_out[17];
    assign wire_8376 = lut_tile_5_8_chanxy_out[18];
    assign wire_8378 = lut_tile_5_8_chanxy_out[19];
    assign wire_8380 = lut_tile_5_8_chanxy_out[20];
    assign wire_8382 = lut_tile_5_8_chanxy_out[21];
    assign wire_8384 = lut_tile_5_8_chanxy_out[22];
    assign wire_8386 = lut_tile_5_8_chanxy_out[23];
    assign wire_8388 = lut_tile_5_8_chanxy_out[24];
    assign wire_8390 = lut_tile_5_8_chanxy_out[25];
    assign wire_8392 = lut_tile_5_8_chanxy_out[26];
    assign wire_8394 = lut_tile_5_8_chanxy_out[27];
    assign wire_8396 = lut_tile_5_8_chanxy_out[28];
    assign wire_8398 = lut_tile_5_8_chanxy_out[29];
    assign wire_13651 = lut_tile_5_8_chanxy_out[30];
    assign wire_13653 = lut_tile_5_8_chanxy_out[31];
    assign wire_13655 = lut_tile_5_8_chanxy_out[32];
    assign wire_13657 = lut_tile_5_8_chanxy_out[33];
    assign wire_13659 = lut_tile_5_8_chanxy_out[34];
    assign wire_13661 = lut_tile_5_8_chanxy_out[35];
    assign wire_13663 = lut_tile_5_8_chanxy_out[36];
    assign wire_13665 = lut_tile_5_8_chanxy_out[37];
    assign wire_13667 = lut_tile_5_8_chanxy_out[38];
    assign wire_13669 = lut_tile_5_8_chanxy_out[39];
    assign wire_13671 = lut_tile_5_8_chanxy_out[40];
    assign wire_13673 = lut_tile_5_8_chanxy_out[41];
    assign wire_13675 = lut_tile_5_8_chanxy_out[42];
    assign wire_13677 = lut_tile_5_8_chanxy_out[43];
    assign wire_13679 = lut_tile_5_8_chanxy_out[44];
    assign wire_13740 = lut_tile_5_8_chanxy_out[45];
    assign wire_13742 = lut_tile_5_8_chanxy_out[46];
    assign wire_13744 = lut_tile_5_8_chanxy_out[47];
    assign wire_13746 = lut_tile_5_8_chanxy_out[48];
    assign wire_13748 = lut_tile_5_8_chanxy_out[49];
    assign wire_13750 = lut_tile_5_8_chanxy_out[50];
    assign wire_13752 = lut_tile_5_8_chanxy_out[51];
    assign wire_13754 = lut_tile_5_8_chanxy_out[52];
    assign wire_13756 = lut_tile_5_8_chanxy_out[53];
    assign wire_13758 = lut_tile_5_8_chanxy_out[54];
    assign wire_13760 = lut_tile_5_8_chanxy_out[55];
    assign wire_13762 = lut_tile_5_8_chanxy_out[56];
    assign wire_13764 = lut_tile_5_8_chanxy_out[57];
    assign wire_13766 = lut_tile_5_8_chanxy_out[58];
    assign wire_13768 = lut_tile_5_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_9_chanxy_in = {wire_14034, wire_8041, wire_8009, wire_8008, wire_7999, wire_7998, wire_7989, wire_7988, wire_7922, wire_5373, wire_14026, wire_8069, wire_7979, wire_7978, wire_7969, wire_7968, wire_7959, wire_7958, wire_7924, wire_5373, wire_14018, wire_8067, wire_8039, wire_8038, wire_8029, wire_8028, wire_8019, wire_8018, wire_7926, wire_5373, wire_14010, wire_8065, wire_8007, wire_8006, wire_7997, wire_7996, wire_7987, wire_7986, wire_7928, wire_4863, wire_14002, wire_8063, wire_7977, wire_7976, wire_7967, wire_7966, wire_7957, wire_7956, wire_7930, wire_4863, wire_13994, wire_8061, wire_8037, wire_8036, wire_8027, wire_8026, wire_8017, wire_8016, wire_7932, wire_4863, wire_13986, wire_8059, wire_8005, wire_8004, wire_7995, wire_7994, wire_7985, wire_7984, wire_7934, wire_5377, wire_4863, wire_13978, wire_8057, wire_7975, wire_7974, wire_7965, wire_7964, wire_7955, wire_7954, wire_7936, wire_5377, wire_4863, wire_13970, wire_8055, wire_8035, wire_8034, wire_8025, wire_8024, wire_8015, wire_8014, wire_7938, wire_5377, wire_4863, wire_13962, wire_8053, wire_8003, wire_8002, wire_7993, wire_7992, wire_7983, wire_7982, wire_7940, wire_5377, wire_4859, wire_13954, wire_8051, wire_7973, wire_7972, wire_7963, wire_7962, wire_7953, wire_7952, wire_7942, wire_5377, wire_4859, wire_13946, wire_8049, wire_8033, wire_8032, wire_8023, wire_8022, wire_8013, wire_8012, wire_7944, wire_5377, wire_4859, wire_13938, wire_8047, wire_8001, wire_8000, wire_7991, wire_7990, wire_7981, wire_7980, wire_7946, wire_5373, wire_4859, wire_13930, wire_8045, wire_7971, wire_7970, wire_7961, wire_7960, wire_7951, wire_7950, wire_7948, wire_5373, wire_4859, wire_13922, wire_8043, wire_8031, wire_8030, wire_8021, wire_8020, wire_8011, wire_8010, wire_7920, wire_5373, wire_4859, wire_14189, wire_8459, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8310, wire_5373, wire_14187, wire_8431, wire_8429, wire_8428, wire_8419, wire_8418, wire_8409, wire_8408, wire_8338, wire_5373, wire_14185, wire_8433, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8336, wire_5373, wire_14183, wire_8435, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8334, wire_4863, wire_14181, wire_8437, wire_8427, wire_8426, wire_8417, wire_8416, wire_8407, wire_8406, wire_8332, wire_4863, wire_14179, wire_8439, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8330, wire_4863, wire_14177, wire_8441, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8328, wire_5377, wire_4863, wire_14175, wire_8443, wire_8425, wire_8424, wire_8415, wire_8414, wire_8405, wire_8404, wire_8326, wire_5377, wire_4863, wire_14173, wire_8445, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8324, wire_5377, wire_4863, wire_14171, wire_8447, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8322, wire_5377, wire_4859, wire_14169, wire_8449, wire_8423, wire_8422, wire_8413, wire_8412, wire_8403, wire_8402, wire_8320, wire_5377, wire_4859, wire_14167, wire_8451, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8318, wire_5377, wire_4859, wire_14165, wire_8453, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8316, wire_5373, wire_4859, wire_14163, wire_8455, wire_8421, wire_8420, wire_8411, wire_8410, wire_8401, wire_8400, wire_8314, wire_5373, wire_4859, wire_14161, wire_8457, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8312, wire_5373, wire_4859, wire_13797, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13678, wire_8308, wire_4902, wire_13795, wire_13709, wire_13708, wire_13699, wire_13698, wire_13689, wire_13688, wire_13650, wire_8306, wire_4902, wire_13793, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13652, wire_8304, wire_4902, wire_13791, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13654, wire_8302, wire_4862, wire_13789, wire_13707, wire_13706, wire_13697, wire_13696, wire_13687, wire_13686, wire_13656, wire_8300, wire_4862, wire_13787, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13658, wire_8298, wire_4862, wire_13785, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13660, wire_8296, wire_4906, wire_4862, wire_13783, wire_13705, wire_13704, wire_13695, wire_13694, wire_13685, wire_13684, wire_13662, wire_8294, wire_4906, wire_4862, wire_13781, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13664, wire_8292, wire_4906, wire_4862, wire_13779, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13666, wire_8290, wire_4906, wire_4858, wire_13777, wire_13703, wire_13702, wire_13693, wire_13692, wire_13683, wire_13682, wire_13668, wire_8288, wire_4906, wire_4858, wire_13775, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13670, wire_8286, wire_4906, wire_4858, wire_13773, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13672, wire_8284, wire_4902, wire_4858, wire_13771, wire_13701, wire_13700, wire_13691, wire_13690, wire_13681, wire_13680, wire_13674, wire_8282, wire_4902, wire_4858, wire_13799, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13676, wire_8280, wire_4902, wire_4858, wire_14163, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14066, wire_8459, wire_4902, wire_14165, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14064, wire_8457, wire_4902, wire_14167, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14062, wire_8455, wire_4902, wire_14169, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14060, wire_8453, wire_4862, wire_14171, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14058, wire_8451, wire_4862, wire_14173, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14056, wire_8449, wire_4862, wire_14175, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_14054, wire_8447, wire_4906, wire_4862, wire_14177, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14052, wire_8445, wire_4906, wire_4862, wire_14179, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14050, wire_8443, wire_4906, wire_4862, wire_14181, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_14048, wire_8441, wire_4906, wire_4858, wire_14183, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14046, wire_8439, wire_4906, wire_4858, wire_14185, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14044, wire_8437, wire_4906, wire_4858, wire_14187, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14042, wire_8435, wire_4902, wire_4858, wire_14189, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14040, wire_8433, wire_4902, wire_4858, wire_14161, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14068, wire_8431, wire_4902, wire_4858};
    // CHNAXY TOTAL: 636
    assign wire_8311 = lut_tile_5_9_chanxy_out[0];
    assign wire_8313 = lut_tile_5_9_chanxy_out[1];
    assign wire_8315 = lut_tile_5_9_chanxy_out[2];
    assign wire_8317 = lut_tile_5_9_chanxy_out[3];
    assign wire_8319 = lut_tile_5_9_chanxy_out[4];
    assign wire_8321 = lut_tile_5_9_chanxy_out[5];
    assign wire_8323 = lut_tile_5_9_chanxy_out[6];
    assign wire_8325 = lut_tile_5_9_chanxy_out[7];
    assign wire_8327 = lut_tile_5_9_chanxy_out[8];
    assign wire_8329 = lut_tile_5_9_chanxy_out[9];
    assign wire_8331 = lut_tile_5_9_chanxy_out[10];
    assign wire_8333 = lut_tile_5_9_chanxy_out[11];
    assign wire_8335 = lut_tile_5_9_chanxy_out[12];
    assign wire_8337 = lut_tile_5_9_chanxy_out[13];
    assign wire_8339 = lut_tile_5_9_chanxy_out[14];
    assign wire_8400 = lut_tile_5_9_chanxy_out[15];
    assign wire_8402 = lut_tile_5_9_chanxy_out[16];
    assign wire_8404 = lut_tile_5_9_chanxy_out[17];
    assign wire_8406 = lut_tile_5_9_chanxy_out[18];
    assign wire_8408 = lut_tile_5_9_chanxy_out[19];
    assign wire_8410 = lut_tile_5_9_chanxy_out[20];
    assign wire_8412 = lut_tile_5_9_chanxy_out[21];
    assign wire_8414 = lut_tile_5_9_chanxy_out[22];
    assign wire_8416 = lut_tile_5_9_chanxy_out[23];
    assign wire_8418 = lut_tile_5_9_chanxy_out[24];
    assign wire_8420 = lut_tile_5_9_chanxy_out[25];
    assign wire_8422 = lut_tile_5_9_chanxy_out[26];
    assign wire_8424 = lut_tile_5_9_chanxy_out[27];
    assign wire_8426 = lut_tile_5_9_chanxy_out[28];
    assign wire_8428 = lut_tile_5_9_chanxy_out[29];
    assign wire_14041 = lut_tile_5_9_chanxy_out[30];
    assign wire_14043 = lut_tile_5_9_chanxy_out[31];
    assign wire_14045 = lut_tile_5_9_chanxy_out[32];
    assign wire_14047 = lut_tile_5_9_chanxy_out[33];
    assign wire_14049 = lut_tile_5_9_chanxy_out[34];
    assign wire_14051 = lut_tile_5_9_chanxy_out[35];
    assign wire_14053 = lut_tile_5_9_chanxy_out[36];
    assign wire_14055 = lut_tile_5_9_chanxy_out[37];
    assign wire_14057 = lut_tile_5_9_chanxy_out[38];
    assign wire_14059 = lut_tile_5_9_chanxy_out[39];
    assign wire_14061 = lut_tile_5_9_chanxy_out[40];
    assign wire_14063 = lut_tile_5_9_chanxy_out[41];
    assign wire_14065 = lut_tile_5_9_chanxy_out[42];
    assign wire_14067 = lut_tile_5_9_chanxy_out[43];
    assign wire_14069 = lut_tile_5_9_chanxy_out[44];
    assign wire_14130 = lut_tile_5_9_chanxy_out[45];
    assign wire_14132 = lut_tile_5_9_chanxy_out[46];
    assign wire_14134 = lut_tile_5_9_chanxy_out[47];
    assign wire_14136 = lut_tile_5_9_chanxy_out[48];
    assign wire_14138 = lut_tile_5_9_chanxy_out[49];
    assign wire_14140 = lut_tile_5_9_chanxy_out[50];
    assign wire_14142 = lut_tile_5_9_chanxy_out[51];
    assign wire_14144 = lut_tile_5_9_chanxy_out[52];
    assign wire_14146 = lut_tile_5_9_chanxy_out[53];
    assign wire_14148 = lut_tile_5_9_chanxy_out[54];
    assign wire_14150 = lut_tile_5_9_chanxy_out[55];
    assign wire_14152 = lut_tile_5_9_chanxy_out[56];
    assign wire_14154 = lut_tile_5_9_chanxy_out[57];
    assign wire_14156 = lut_tile_5_9_chanxy_out[58];
    assign wire_14158 = lut_tile_5_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_5_10_chanxy_in = {wire_14426, wire_8054, wire_8032, wire_8008, wire_7956, wire_5878, wire_5872, wire_5863, wire_5857, wire_14418, wire_8046, wire_8024, wire_8000, wire_7978, wire_5878, wire_5872, wire_5863, wire_5857, wire_14410, wire_8068, wire_8016, wire_7992, wire_7970, wire_5878, wire_5872, wire_5863, wire_5857, wire_14402, wire_8060, wire_8038, wire_7984, wire_7962, wire_5878, wire_5869, wire_5863, wire_5379, wire_14394, wire_8052, wire_8030, wire_8006, wire_7954, wire_5878, wire_5869, wire_5863, wire_5379, wire_14386, wire_8044, wire_8022, wire_7998, wire_7976, wire_5878, wire_5869, wire_5863, wire_5379, wire_14378, wire_8066, wire_8014, wire_7990, wire_7968, wire_5875, wire_5869, wire_5860, wire_5379, wire_14370, wire_8058, wire_8036, wire_7982, wire_7960, wire_5875, wire_5869, wire_5860, wire_5379, wire_14362, wire_8050, wire_8028, wire_8004, wire_7952, wire_5875, wire_5869, wire_5860, wire_5379, wire_14354, wire_8042, wire_8020, wire_7996, wire_7974, wire_5875, wire_5866, wire_5860, wire_5375, wire_14346, wire_8064, wire_8012, wire_7988, wire_7966, wire_5875, wire_5866, wire_5860, wire_5375, wire_14338, wire_8056, wire_8034, wire_7980, wire_7958, wire_5875, wire_5866, wire_5860, wire_5375, wire_14330, wire_8048, wire_8026, wire_8002, wire_7950, wire_5872, wire_5866, wire_5857, wire_5375, wire_14322, wire_8040, wire_8018, wire_7994, wire_7972, wire_5872, wire_5866, wire_5857, wire_5375, wire_14314, wire_8062, wire_8010, wire_7986, wire_7964, wire_5872, wire_5866, wire_5857, wire_5375, wire_14579, wire_8436, wire_8414, wire_8392, wire_8368, wire_5878, wire_5872, wire_5863, wire_5857, wire_14577, wire_8458, wire_8406, wire_8384, wire_8360, wire_5878, wire_5872, wire_5863, wire_5857, wire_14575, wire_8450, wire_8428, wire_8376, wire_8352, wire_5878, wire_5872, wire_5863, wire_5857, wire_14573, wire_8442, wire_8420, wire_8398, wire_8344, wire_5878, wire_5869, wire_5863, wire_5379, wire_14571, wire_8434, wire_8412, wire_8390, wire_8366, wire_5878, wire_5869, wire_5863, wire_5379, wire_14569, wire_8456, wire_8404, wire_8382, wire_8358, wire_5878, wire_5869, wire_5863, wire_5379, wire_14567, wire_8448, wire_8426, wire_8374, wire_8350, wire_5875, wire_5869, wire_5860, wire_5379, wire_14565, wire_8440, wire_8418, wire_8396, wire_8342, wire_5875, wire_5869, wire_5860, wire_5379, wire_14563, wire_8432, wire_8410, wire_8388, wire_8364, wire_5875, wire_5869, wire_5860, wire_5379, wire_14561, wire_8454, wire_8402, wire_8380, wire_8356, wire_5875, wire_5866, wire_5860, wire_5375, wire_14559, wire_8446, wire_8424, wire_8372, wire_8348, wire_5875, wire_5866, wire_5860, wire_5375, wire_14557, wire_8438, wire_8416, wire_8394, wire_8340, wire_5875, wire_5866, wire_5860, wire_5375, wire_14555, wire_8430, wire_8408, wire_8386, wire_8362, wire_5872, wire_5866, wire_5857, wire_5375, wire_14553, wire_8452, wire_8400, wire_8378, wire_8354, wire_5872, wire_5866, wire_5857, wire_5375, wire_14551, wire_8444, wire_8422, wire_8370, wire_8346, wire_5872, wire_5866, wire_5857, wire_5375, wire_14549, wire_14548, wire_14187, wire_14099, wire_14098, wire_14089, wire_14088, wire_14079, wire_14078, wire_14068, wire_8338, wire_5418, wire_14533, wire_14532, wire_14185, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14040, wire_8336, wire_5418, wire_14517, wire_14516, wire_14183, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14042, wire_8334, wire_5418, wire_14531, wire_14530, wire_14181, wire_14097, wire_14096, wire_14087, wire_14086, wire_14077, wire_14076, wire_14044, wire_8332, wire_5378, wire_14545, wire_14544, wire_14179, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14046, wire_8330, wire_5378, wire_14499, wire_14498, wire_14177, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14048, wire_8328, wire_5378, wire_14543, wire_14542, wire_14175, wire_14095, wire_14094, wire_14085, wire_14084, wire_14075, wire_14074, wire_14050, wire_8326, wire_5422, wire_5378, wire_14527, wire_14526, wire_14173, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14052, wire_8324, wire_5422, wire_5378, wire_14511, wire_14510, wire_14171, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14054, wire_8322, wire_5422, wire_5378, wire_14525, wire_14524, wire_5422, wire_14169, wire_14093, wire_14092, wire_14083, wire_14082, wire_14073, wire_14072, wire_14056, wire_8320, wire_5422, wire_5374, wire_14539, wire_14538, wire_5422, wire_14167, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14058, wire_8318, wire_5422, wire_5374, wire_14493, wire_14492, wire_5418, wire_14165, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14060, wire_8316, wire_5422, wire_5374, wire_14537, wire_14536, wire_5378, wire_14163, wire_14091, wire_14090, wire_14081, wire_14080, wire_14071, wire_14070, wire_14062, wire_8314, wire_5418, wire_5374, wire_14521, wire_14520, wire_5378, wire_14161, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14064, wire_8312, wire_5418, wire_5374, wire_14505, wire_14504, wire_5374, wire_14189, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14066, wire_8310, wire_5418, wire_5374, wire_14563, wire_14442, wire_14577, wire_14456, wire_14487, wire_14486, wire_14575, wire_14454, wire_14559, wire_14438, wire_14469, wire_14468, wire_14557, wire_14436, wire_14571, wire_14450, wire_14481, wire_14480, wire_14569, wire_14448, wire_5422, wire_14553, wire_14432, wire_5418, wire_14463, wire_14462, wire_5418, wire_14551, wire_14430, wire_5378, wire_14565, wire_14444, wire_5374, wire_14475, wire_14474, wire_5374, wire_14519, wire_14518, wire_14547, wire_14546, wire_14473, wire_14472, wire_14501, wire_14500, wire_14529, wire_14528, wire_14485, wire_14484, wire_14513, wire_14512, wire_14541, wire_14540, wire_14467, wire_14466, wire_14495, wire_14494, wire_5422, wire_14523, wire_14522, wire_5418, wire_14479, wire_14478, wire_5418, wire_14507, wire_14506, wire_5378, wire_14535, wire_14534, wire_5374, wire_14461, wire_14460, wire_5374, wire_14579, wire_14458, wire_14489, wire_14488, wire_14503, wire_14502, wire_14561, wire_14440, wire_14471, wire_14470, wire_14515, wire_14514, wire_14573, wire_14452, wire_14483, wire_14482, wire_14497, wire_14496, wire_14555, wire_14434, wire_5422, wire_14465, wire_14464, wire_5422, wire_14509, wire_14508, wire_5418, wire_14567, wire_14446, wire_5378, wire_14477, wire_14476, wire_5378, wire_14491, wire_14490, wire_5374};
    // CHNAXY TOTAL: 573
    assign wire_8341 = lut_tile_5_10_chanxy_out[0];
    assign wire_8343 = lut_tile_5_10_chanxy_out[1];
    assign wire_8345 = lut_tile_5_10_chanxy_out[2];
    assign wire_8347 = lut_tile_5_10_chanxy_out[3];
    assign wire_8349 = lut_tile_5_10_chanxy_out[4];
    assign wire_8351 = lut_tile_5_10_chanxy_out[5];
    assign wire_8353 = lut_tile_5_10_chanxy_out[6];
    assign wire_8355 = lut_tile_5_10_chanxy_out[7];
    assign wire_8357 = lut_tile_5_10_chanxy_out[8];
    assign wire_8359 = lut_tile_5_10_chanxy_out[9];
    assign wire_8361 = lut_tile_5_10_chanxy_out[10];
    assign wire_8363 = lut_tile_5_10_chanxy_out[11];
    assign wire_8365 = lut_tile_5_10_chanxy_out[12];
    assign wire_8367 = lut_tile_5_10_chanxy_out[13];
    assign wire_8369 = lut_tile_5_10_chanxy_out[14];
    assign wire_8371 = lut_tile_5_10_chanxy_out[15];
    assign wire_8373 = lut_tile_5_10_chanxy_out[16];
    assign wire_8375 = lut_tile_5_10_chanxy_out[17];
    assign wire_8377 = lut_tile_5_10_chanxy_out[18];
    assign wire_8379 = lut_tile_5_10_chanxy_out[19];
    assign wire_8381 = lut_tile_5_10_chanxy_out[20];
    assign wire_8383 = lut_tile_5_10_chanxy_out[21];
    assign wire_8385 = lut_tile_5_10_chanxy_out[22];
    assign wire_8387 = lut_tile_5_10_chanxy_out[23];
    assign wire_8389 = lut_tile_5_10_chanxy_out[24];
    assign wire_8391 = lut_tile_5_10_chanxy_out[25];
    assign wire_8393 = lut_tile_5_10_chanxy_out[26];
    assign wire_8395 = lut_tile_5_10_chanxy_out[27];
    assign wire_8397 = lut_tile_5_10_chanxy_out[28];
    assign wire_8399 = lut_tile_5_10_chanxy_out[29];
    assign wire_8401 = lut_tile_5_10_chanxy_out[30];
    assign wire_8403 = lut_tile_5_10_chanxy_out[31];
    assign wire_8405 = lut_tile_5_10_chanxy_out[32];
    assign wire_8407 = lut_tile_5_10_chanxy_out[33];
    assign wire_8409 = lut_tile_5_10_chanxy_out[34];
    assign wire_8411 = lut_tile_5_10_chanxy_out[35];
    assign wire_8413 = lut_tile_5_10_chanxy_out[36];
    assign wire_8415 = lut_tile_5_10_chanxy_out[37];
    assign wire_8417 = lut_tile_5_10_chanxy_out[38];
    assign wire_8419 = lut_tile_5_10_chanxy_out[39];
    assign wire_8421 = lut_tile_5_10_chanxy_out[40];
    assign wire_8423 = lut_tile_5_10_chanxy_out[41];
    assign wire_8425 = lut_tile_5_10_chanxy_out[42];
    assign wire_8427 = lut_tile_5_10_chanxy_out[43];
    assign wire_8429 = lut_tile_5_10_chanxy_out[44];
    assign wire_8430 = lut_tile_5_10_chanxy_out[45];
    assign wire_8431 = lut_tile_5_10_chanxy_out[46];
    assign wire_8432 = lut_tile_5_10_chanxy_out[47];
    assign wire_8433 = lut_tile_5_10_chanxy_out[48];
    assign wire_8434 = lut_tile_5_10_chanxy_out[49];
    assign wire_8435 = lut_tile_5_10_chanxy_out[50];
    assign wire_8436 = lut_tile_5_10_chanxy_out[51];
    assign wire_8437 = lut_tile_5_10_chanxy_out[52];
    assign wire_8438 = lut_tile_5_10_chanxy_out[53];
    assign wire_8439 = lut_tile_5_10_chanxy_out[54];
    assign wire_8440 = lut_tile_5_10_chanxy_out[55];
    assign wire_8441 = lut_tile_5_10_chanxy_out[56];
    assign wire_8442 = lut_tile_5_10_chanxy_out[57];
    assign wire_8443 = lut_tile_5_10_chanxy_out[58];
    assign wire_8444 = lut_tile_5_10_chanxy_out[59];
    assign wire_8445 = lut_tile_5_10_chanxy_out[60];
    assign wire_8446 = lut_tile_5_10_chanxy_out[61];
    assign wire_8447 = lut_tile_5_10_chanxy_out[62];
    assign wire_8448 = lut_tile_5_10_chanxy_out[63];
    assign wire_8449 = lut_tile_5_10_chanxy_out[64];
    assign wire_8450 = lut_tile_5_10_chanxy_out[65];
    assign wire_8451 = lut_tile_5_10_chanxy_out[66];
    assign wire_8452 = lut_tile_5_10_chanxy_out[67];
    assign wire_8453 = lut_tile_5_10_chanxy_out[68];
    assign wire_8454 = lut_tile_5_10_chanxy_out[69];
    assign wire_8455 = lut_tile_5_10_chanxy_out[70];
    assign wire_8456 = lut_tile_5_10_chanxy_out[71];
    assign wire_8457 = lut_tile_5_10_chanxy_out[72];
    assign wire_8458 = lut_tile_5_10_chanxy_out[73];
    assign wire_8459 = lut_tile_5_10_chanxy_out[74];
    assign wire_14431 = lut_tile_5_10_chanxy_out[75];
    assign wire_14433 = lut_tile_5_10_chanxy_out[76];
    assign wire_14435 = lut_tile_5_10_chanxy_out[77];
    assign wire_14437 = lut_tile_5_10_chanxy_out[78];
    assign wire_14439 = lut_tile_5_10_chanxy_out[79];
    assign wire_14441 = lut_tile_5_10_chanxy_out[80];
    assign wire_14443 = lut_tile_5_10_chanxy_out[81];
    assign wire_14445 = lut_tile_5_10_chanxy_out[82];
    assign wire_14447 = lut_tile_5_10_chanxy_out[83];
    assign wire_14449 = lut_tile_5_10_chanxy_out[84];
    assign wire_14451 = lut_tile_5_10_chanxy_out[85];
    assign wire_14453 = lut_tile_5_10_chanxy_out[86];
    assign wire_14455 = lut_tile_5_10_chanxy_out[87];
    assign wire_14457 = lut_tile_5_10_chanxy_out[88];
    assign wire_14459 = lut_tile_5_10_chanxy_out[89];
    assign wire_14520 = lut_tile_5_10_chanxy_out[90];
    assign wire_14522 = lut_tile_5_10_chanxy_out[91];
    assign wire_14524 = lut_tile_5_10_chanxy_out[92];
    assign wire_14526 = lut_tile_5_10_chanxy_out[93];
    assign wire_14528 = lut_tile_5_10_chanxy_out[94];
    assign wire_14530 = lut_tile_5_10_chanxy_out[95];
    assign wire_14532 = lut_tile_5_10_chanxy_out[96];
    assign wire_14534 = lut_tile_5_10_chanxy_out[97];
    assign wire_14536 = lut_tile_5_10_chanxy_out[98];
    assign wire_14538 = lut_tile_5_10_chanxy_out[99];
    assign wire_14540 = lut_tile_5_10_chanxy_out[100];
    assign wire_14542 = lut_tile_5_10_chanxy_out[101];
    assign wire_14544 = lut_tile_5_10_chanxy_out[102];
    assign wire_14546 = lut_tile_5_10_chanxy_out[103];
    assign wire_14548 = lut_tile_5_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_6_1_chanxy_in = {wire_10948, wire_8191, wire_8189, wire_8188, wire_8149, wire_8148, wire_8109, wire_8108, wire_8082, wire_1287, wire_10946, wire_8219, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_8090, wire_1287, wire_10944, wire_8217, wire_8183, wire_8182, wire_8143, wire_8142, wire_8103, wire_8102, wire_8098, wire_1287, wire_10942, wire_8215, wire_8181, wire_8180, wire_8141, wire_8140, wire_8106, wire_8101, wire_8100, wire_777, wire_10940, wire_8213, wire_8177, wire_8176, wire_8137, wire_8136, wire_8114, wire_8097, wire_8096, wire_777, wire_10938, wire_8211, wire_8175, wire_8174, wire_8135, wire_8134, wire_8122, wire_8095, wire_8094, wire_777, wire_10936, wire_8209, wire_8173, wire_8172, wire_8133, wire_8132, wire_8130, wire_8093, wire_8092, wire_1291, wire_777, wire_10934, wire_8207, wire_8169, wire_8168, wire_8138, wire_8129, wire_8128, wire_8089, wire_8088, wire_1291, wire_777, wire_10932, wire_8205, wire_8167, wire_8166, wire_8146, wire_8127, wire_8126, wire_8087, wire_8086, wire_1291, wire_777, wire_10930, wire_8203, wire_8165, wire_8164, wire_8154, wire_8125, wire_8124, wire_8085, wire_8084, wire_1291, wire_773, wire_10928, wire_8201, wire_8162, wire_8161, wire_8160, wire_8121, wire_8120, wire_8081, wire_8080, wire_1291, wire_773, wire_10926, wire_8199, wire_8170, wire_8159, wire_8158, wire_8119, wire_8118, wire_8079, wire_8078, wire_1291, wire_773, wire_10924, wire_8197, wire_8178, wire_8157, wire_8156, wire_8117, wire_8116, wire_8077, wire_8076, wire_1287, wire_773, wire_10922, wire_8195, wire_8186, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072, wire_1287, wire_773, wire_10920, wire_8193, wire_8151, wire_8150, wire_8111, wire_8110, wire_8074, wire_8071, wire_8070, wire_1287, wire_773, wire_11099, wire_8609, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_8466, wire_1287, wire_11097, wire_8581, wire_8578, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_1287, wire_11095, wire_8583, wire_8573, wire_8572, wire_8570, wire_8533, wire_8532, wire_8493, wire_8492, wire_1287, wire_11093, wire_8585, wire_8569, wire_8568, wire_8562, wire_8529, wire_8528, wire_8489, wire_8488, wire_777, wire_11091, wire_8587, wire_8567, wire_8566, wire_8554, wire_8527, wire_8526, wire_8487, wire_8486, wire_777, wire_11089, wire_8589, wire_8565, wire_8564, wire_8546, wire_8525, wire_8524, wire_8485, wire_8484, wire_777, wire_11087, wire_8591, wire_8561, wire_8560, wire_8538, wire_8521, wire_8520, wire_8481, wire_8480, wire_1291, wire_777, wire_11085, wire_8593, wire_8559, wire_8558, wire_8530, wire_8519, wire_8518, wire_8479, wire_8478, wire_1291, wire_777, wire_11083, wire_8595, wire_8557, wire_8556, wire_8522, wire_8517, wire_8516, wire_8477, wire_8476, wire_1291, wire_777, wire_11081, wire_8597, wire_8553, wire_8552, wire_8514, wire_8513, wire_8512, wire_8473, wire_8472, wire_1291, wire_773, wire_11079, wire_8599, wire_8551, wire_8550, wire_8511, wire_8510, wire_8506, wire_8471, wire_8470, wire_1291, wire_773, wire_11077, wire_8601, wire_8549, wire_8548, wire_8509, wire_8508, wire_8498, wire_8469, wire_8468, wire_1291, wire_773, wire_11075, wire_8603, wire_8545, wire_8544, wire_8505, wire_8504, wire_8490, wire_8465, wire_8464, wire_1287, wire_773, wire_11073, wire_8605, wire_8543, wire_8542, wire_8503, wire_8502, wire_8482, wire_8463, wire_8462, wire_1287, wire_773, wire_11071, wire_8607, wire_8541, wire_8540, wire_8501, wire_8500, wire_8474, wire_8461, wire_8460, wire_1287, wire_773, wire_11073, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_10976, wire_8609, wire_816, wire_10603, wire_10602, wire_10619, wire_10618, wire_10709, wire_10588, wire_10693, wire_10572, wire_11075, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10974, wire_8607, wire_816, wire_10679, wire_10678, wire_10649, wire_10648, wire_10663, wire_10662, wire_10617, wire_10616, wire_11077, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10972, wire_8605, wire_816, wire_10707, wire_10586, wire_10633, wire_10632, wire_10677, wire_10676, wire_10647, wire_10646, wire_11079, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_10970, wire_8603, wire_776, wire_10615, wire_10614, wire_10601, wire_10600, wire_10691, wire_10570, wire_10705, wire_10584, wire_11081, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10968, wire_8601, wire_776, wire_10661, wire_10660, wire_10631, wire_10630, wire_10675, wire_10674, wire_10599, wire_10598, wire_11083, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10966, wire_8599, wire_776, wire_10689, wire_10568, wire_10645, wire_10644, wire_10659, wire_10658, wire_10629, wire_10628, wire_11085, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_10964, wire_8597, wire_820, wire_776, wire_10597, wire_10596, wire_10613, wire_10612, wire_10703, wire_10582, wire_10687, wire_10566, wire_11087, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10962, wire_8595, wire_820, wire_776, wire_10673, wire_10672, wire_10643, wire_10642, wire_10657, wire_10656, wire_10611, wire_10610, wire_11089, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10960, wire_8593, wire_820, wire_776, wire_10701, wire_10580, wire_10627, wire_10626, wire_10671, wire_10670, wire_10641, wire_10640, wire_11091, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_10958, wire_8591, wire_820, wire_772, wire_10609, wire_10608, wire_820, wire_10595, wire_10594, wire_820, wire_10685, wire_10564, wire_820, wire_10699, wire_10578, wire_820, wire_11093, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10956, wire_8589, wire_820, wire_772, wire_10655, wire_10654, wire_820, wire_10625, wire_10624, wire_820, wire_10669, wire_10668, wire_816, wire_10593, wire_10592, wire_816, wire_11095, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10954, wire_8587, wire_820, wire_772, wire_10683, wire_10562, wire_816, wire_10639, wire_10638, wire_816, wire_10653, wire_10652, wire_816, wire_10623, wire_10622, wire_816, wire_11097, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_10952, wire_8585, wire_816, wire_772, wire_10591, wire_10590, wire_776, wire_10607, wire_10606, wire_776, wire_10697, wire_10576, wire_776, wire_10681, wire_10560, wire_776, wire_11099, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10950, wire_8583, wire_816, wire_772, wire_10667, wire_10666, wire_776, wire_10637, wire_10636, wire_776, wire_10651, wire_10650, wire_772, wire_10605, wire_10604, wire_772, wire_11071, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10978, wire_8581, wire_816, wire_772, wire_10695, wire_10574, wire_772, wire_10621, wire_10620, wire_772, wire_10665, wire_10664, wire_772, wire_10635, wire_10634, wire_772};
    // CHNAXY TOTAL: 621
    assign wire_8460 = lut_tile_6_1_chanxy_out[0];
    assign wire_8462 = lut_tile_6_1_chanxy_out[1];
    assign wire_8464 = lut_tile_6_1_chanxy_out[2];
    assign wire_8466 = lut_tile_6_1_chanxy_out[3];
    assign wire_8467 = lut_tile_6_1_chanxy_out[4];
    assign wire_8468 = lut_tile_6_1_chanxy_out[5];
    assign wire_8470 = lut_tile_6_1_chanxy_out[6];
    assign wire_8472 = lut_tile_6_1_chanxy_out[7];
    assign wire_8474 = lut_tile_6_1_chanxy_out[8];
    assign wire_8475 = lut_tile_6_1_chanxy_out[9];
    assign wire_8476 = lut_tile_6_1_chanxy_out[10];
    assign wire_8478 = lut_tile_6_1_chanxy_out[11];
    assign wire_8480 = lut_tile_6_1_chanxy_out[12];
    assign wire_8482 = lut_tile_6_1_chanxy_out[13];
    assign wire_8483 = lut_tile_6_1_chanxy_out[14];
    assign wire_8484 = lut_tile_6_1_chanxy_out[15];
    assign wire_8486 = lut_tile_6_1_chanxy_out[16];
    assign wire_8488 = lut_tile_6_1_chanxy_out[17];
    assign wire_8490 = lut_tile_6_1_chanxy_out[18];
    assign wire_8491 = lut_tile_6_1_chanxy_out[19];
    assign wire_8492 = lut_tile_6_1_chanxy_out[20];
    assign wire_8494 = lut_tile_6_1_chanxy_out[21];
    assign wire_8496 = lut_tile_6_1_chanxy_out[22];
    assign wire_8498 = lut_tile_6_1_chanxy_out[23];
    assign wire_8499 = lut_tile_6_1_chanxy_out[24];
    assign wire_8500 = lut_tile_6_1_chanxy_out[25];
    assign wire_8502 = lut_tile_6_1_chanxy_out[26];
    assign wire_8504 = lut_tile_6_1_chanxy_out[27];
    assign wire_8506 = lut_tile_6_1_chanxy_out[28];
    assign wire_8507 = lut_tile_6_1_chanxy_out[29];
    assign wire_8508 = lut_tile_6_1_chanxy_out[30];
    assign wire_8510 = lut_tile_6_1_chanxy_out[31];
    assign wire_8512 = lut_tile_6_1_chanxy_out[32];
    assign wire_8514 = lut_tile_6_1_chanxy_out[33];
    assign wire_8515 = lut_tile_6_1_chanxy_out[34];
    assign wire_8516 = lut_tile_6_1_chanxy_out[35];
    assign wire_8518 = lut_tile_6_1_chanxy_out[36];
    assign wire_8520 = lut_tile_6_1_chanxy_out[37];
    assign wire_8522 = lut_tile_6_1_chanxy_out[38];
    assign wire_8523 = lut_tile_6_1_chanxy_out[39];
    assign wire_8524 = lut_tile_6_1_chanxy_out[40];
    assign wire_8526 = lut_tile_6_1_chanxy_out[41];
    assign wire_8528 = lut_tile_6_1_chanxy_out[42];
    assign wire_8530 = lut_tile_6_1_chanxy_out[43];
    assign wire_8531 = lut_tile_6_1_chanxy_out[44];
    assign wire_8532 = lut_tile_6_1_chanxy_out[45];
    assign wire_8534 = lut_tile_6_1_chanxy_out[46];
    assign wire_8536 = lut_tile_6_1_chanxy_out[47];
    assign wire_8538 = lut_tile_6_1_chanxy_out[48];
    assign wire_8539 = lut_tile_6_1_chanxy_out[49];
    assign wire_8540 = lut_tile_6_1_chanxy_out[50];
    assign wire_8542 = lut_tile_6_1_chanxy_out[51];
    assign wire_8544 = lut_tile_6_1_chanxy_out[52];
    assign wire_8546 = lut_tile_6_1_chanxy_out[53];
    assign wire_8547 = lut_tile_6_1_chanxy_out[54];
    assign wire_8548 = lut_tile_6_1_chanxy_out[55];
    assign wire_8550 = lut_tile_6_1_chanxy_out[56];
    assign wire_8552 = lut_tile_6_1_chanxy_out[57];
    assign wire_8554 = lut_tile_6_1_chanxy_out[58];
    assign wire_8555 = lut_tile_6_1_chanxy_out[59];
    assign wire_8556 = lut_tile_6_1_chanxy_out[60];
    assign wire_8558 = lut_tile_6_1_chanxy_out[61];
    assign wire_8560 = lut_tile_6_1_chanxy_out[62];
    assign wire_8562 = lut_tile_6_1_chanxy_out[63];
    assign wire_8563 = lut_tile_6_1_chanxy_out[64];
    assign wire_8564 = lut_tile_6_1_chanxy_out[65];
    assign wire_8566 = lut_tile_6_1_chanxy_out[66];
    assign wire_8568 = lut_tile_6_1_chanxy_out[67];
    assign wire_8570 = lut_tile_6_1_chanxy_out[68];
    assign wire_8571 = lut_tile_6_1_chanxy_out[69];
    assign wire_8572 = lut_tile_6_1_chanxy_out[70];
    assign wire_8574 = lut_tile_6_1_chanxy_out[71];
    assign wire_8576 = lut_tile_6_1_chanxy_out[72];
    assign wire_8578 = lut_tile_6_1_chanxy_out[73];
    assign wire_8579 = lut_tile_6_1_chanxy_out[74];
    assign wire_10951 = lut_tile_6_1_chanxy_out[75];
    assign wire_10953 = lut_tile_6_1_chanxy_out[76];
    assign wire_10955 = lut_tile_6_1_chanxy_out[77];
    assign wire_10957 = lut_tile_6_1_chanxy_out[78];
    assign wire_10959 = lut_tile_6_1_chanxy_out[79];
    assign wire_10961 = lut_tile_6_1_chanxy_out[80];
    assign wire_10963 = lut_tile_6_1_chanxy_out[81];
    assign wire_10965 = lut_tile_6_1_chanxy_out[82];
    assign wire_10967 = lut_tile_6_1_chanxy_out[83];
    assign wire_10969 = lut_tile_6_1_chanxy_out[84];
    assign wire_10971 = lut_tile_6_1_chanxy_out[85];
    assign wire_10973 = lut_tile_6_1_chanxy_out[86];
    assign wire_10975 = lut_tile_6_1_chanxy_out[87];
    assign wire_10977 = lut_tile_6_1_chanxy_out[88];
    assign wire_10979 = lut_tile_6_1_chanxy_out[89];
    assign wire_11040 = lut_tile_6_1_chanxy_out[90];
    assign wire_11042 = lut_tile_6_1_chanxy_out[91];
    assign wire_11044 = lut_tile_6_1_chanxy_out[92];
    assign wire_11046 = lut_tile_6_1_chanxy_out[93];
    assign wire_11048 = lut_tile_6_1_chanxy_out[94];
    assign wire_11050 = lut_tile_6_1_chanxy_out[95];
    assign wire_11052 = lut_tile_6_1_chanxy_out[96];
    assign wire_11054 = lut_tile_6_1_chanxy_out[97];
    assign wire_11056 = lut_tile_6_1_chanxy_out[98];
    assign wire_11058 = lut_tile_6_1_chanxy_out[99];
    assign wire_11060 = lut_tile_6_1_chanxy_out[100];
    assign wire_11062 = lut_tile_6_1_chanxy_out[101];
    assign wire_11064 = lut_tile_6_1_chanxy_out[102];
    assign wire_11066 = lut_tile_6_1_chanxy_out[103];
    assign wire_11068 = lut_tile_6_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_6_2_chanxy_in = {wire_11338, wire_8221, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8084, wire_1803, wire_11336, wire_8249, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_8092, wire_1803, wire_11334, wire_8247, wire_8183, wire_8182, wire_8143, wire_8142, wire_8103, wire_8102, wire_8100, wire_1803, wire_11332, wire_8245, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8108, wire_1293, wire_11330, wire_8243, wire_8177, wire_8176, wire_8137, wire_8136, wire_8116, wire_8097, wire_8096, wire_1293, wire_11328, wire_8241, wire_8175, wire_8174, wire_8135, wire_8134, wire_8124, wire_8095, wire_8094, wire_1293, wire_11326, wire_8239, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8132, wire_1807, wire_1293, wire_11324, wire_8237, wire_8169, wire_8168, wire_8140, wire_8129, wire_8128, wire_8089, wire_8088, wire_1807, wire_1293, wire_11322, wire_8235, wire_8167, wire_8166, wire_8148, wire_8127, wire_8126, wire_8087, wire_8086, wire_1807, wire_1293, wire_11320, wire_8233, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8156, wire_1807, wire_1289, wire_11318, wire_8231, wire_8164, wire_8161, wire_8160, wire_8121, wire_8120, wire_8081, wire_8080, wire_1807, wire_1289, wire_11316, wire_8229, wire_8172, wire_8159, wire_8158, wire_8119, wire_8118, wire_8079, wire_8078, wire_1807, wire_1289, wire_11314, wire_8227, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8180, wire_1803, wire_1289, wire_11312, wire_8225, wire_8188, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072, wire_1803, wire_1289, wire_11310, wire_8223, wire_8151, wire_8150, wire_8111, wire_8110, wire_8076, wire_8071, wire_8070, wire_1803, wire_1289, wire_11489, wire_8639, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8460, wire_1803, wire_11487, wire_8611, wire_8577, wire_8576, wire_8572, wire_8537, wire_8536, wire_8497, wire_8496, wire_1803, wire_11485, wire_8613, wire_8575, wire_8574, wire_8564, wire_8535, wire_8534, wire_8495, wire_8494, wire_1803, wire_11483, wire_8615, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8556, wire_1293, wire_11481, wire_8617, wire_8569, wire_8568, wire_8548, wire_8529, wire_8528, wire_8489, wire_8488, wire_1293, wire_11479, wire_8619, wire_8567, wire_8566, wire_8540, wire_8527, wire_8526, wire_8487, wire_8486, wire_1293, wire_11477, wire_8621, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8532, wire_1807, wire_1293, wire_11475, wire_8623, wire_8561, wire_8560, wire_8524, wire_8521, wire_8520, wire_8481, wire_8480, wire_1807, wire_1293, wire_11473, wire_8625, wire_8559, wire_8558, wire_8519, wire_8518, wire_8516, wire_8479, wire_8478, wire_1807, wire_1293, wire_11471, wire_8627, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8508, wire_1807, wire_1289, wire_11469, wire_8629, wire_8553, wire_8552, wire_8513, wire_8512, wire_8500, wire_8473, wire_8472, wire_1807, wire_1289, wire_11467, wire_8631, wire_8551, wire_8550, wire_8511, wire_8510, wire_8492, wire_8471, wire_8470, wire_1807, wire_1289, wire_11465, wire_8633, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8484, wire_1803, wire_1289, wire_11463, wire_8635, wire_8545, wire_8544, wire_8505, wire_8504, wire_8476, wire_8465, wire_8464, wire_1803, wire_1289, wire_11461, wire_8637, wire_8543, wire_8542, wire_8503, wire_8502, wire_8468, wire_8463, wire_8462, wire_1803, wire_1289, wire_11097, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_10978, wire_8578, wire_1332, wire_11095, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10950, wire_8570, wire_1332, wire_11093, wire_11009, wire_11008, wire_10999, wire_10998, wire_10989, wire_10988, wire_10952, wire_8562, wire_1332, wire_11091, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_10954, wire_8554, wire_1292, wire_11089, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10956, wire_8546, wire_1292, wire_11087, wire_11007, wire_11006, wire_10997, wire_10996, wire_10987, wire_10986, wire_10958, wire_8538, wire_1292, wire_11085, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_10960, wire_8530, wire_1336, wire_1292, wire_11083, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10962, wire_8522, wire_1336, wire_1292, wire_11081, wire_11005, wire_11004, wire_10995, wire_10994, wire_10985, wire_10984, wire_10964, wire_8514, wire_1336, wire_1292, wire_11079, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_10966, wire_8506, wire_1336, wire_1288, wire_11077, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10968, wire_8498, wire_1336, wire_1288, wire_11075, wire_11003, wire_11002, wire_10993, wire_10992, wire_10983, wire_10982, wire_10970, wire_8490, wire_1336, wire_1288, wire_11073, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_10972, wire_8482, wire_1332, wire_1288, wire_11071, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_10974, wire_8474, wire_1332, wire_1288, wire_11099, wire_11001, wire_11000, wire_10991, wire_10990, wire_10981, wire_10980, wire_10976, wire_8466, wire_1332, wire_1288, wire_11463, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11366, wire_8639, wire_1332, wire_11465, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11364, wire_8637, wire_1332, wire_11467, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11362, wire_8635, wire_1332, wire_11469, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11360, wire_8633, wire_1292, wire_11471, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11358, wire_8631, wire_1292, wire_11473, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11356, wire_8629, wire_1292, wire_11475, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11354, wire_8627, wire_1336, wire_1292, wire_11477, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11352, wire_8625, wire_1336, wire_1292, wire_11479, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11350, wire_8623, wire_1336, wire_1292, wire_11481, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11348, wire_8621, wire_1336, wire_1288, wire_11483, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11346, wire_8619, wire_1336, wire_1288, wire_11485, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11344, wire_8617, wire_1336, wire_1288, wire_11487, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11342, wire_8615, wire_1332, wire_1288, wire_11489, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11340, wire_8613, wire_1332, wire_1288, wire_11461, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11368, wire_8611, wire_1332, wire_1288};
    // CHNAXY TOTAL: 636
    assign wire_8461 = lut_tile_6_2_chanxy_out[0];
    assign wire_8469 = lut_tile_6_2_chanxy_out[1];
    assign wire_8477 = lut_tile_6_2_chanxy_out[2];
    assign wire_8485 = lut_tile_6_2_chanxy_out[3];
    assign wire_8493 = lut_tile_6_2_chanxy_out[4];
    assign wire_8501 = lut_tile_6_2_chanxy_out[5];
    assign wire_8509 = lut_tile_6_2_chanxy_out[6];
    assign wire_8517 = lut_tile_6_2_chanxy_out[7];
    assign wire_8525 = lut_tile_6_2_chanxy_out[8];
    assign wire_8533 = lut_tile_6_2_chanxy_out[9];
    assign wire_8541 = lut_tile_6_2_chanxy_out[10];
    assign wire_8549 = lut_tile_6_2_chanxy_out[11];
    assign wire_8557 = lut_tile_6_2_chanxy_out[12];
    assign wire_8565 = lut_tile_6_2_chanxy_out[13];
    assign wire_8573 = lut_tile_6_2_chanxy_out[14];
    assign wire_8580 = lut_tile_6_2_chanxy_out[15];
    assign wire_8582 = lut_tile_6_2_chanxy_out[16];
    assign wire_8584 = lut_tile_6_2_chanxy_out[17];
    assign wire_8586 = lut_tile_6_2_chanxy_out[18];
    assign wire_8588 = lut_tile_6_2_chanxy_out[19];
    assign wire_8590 = lut_tile_6_2_chanxy_out[20];
    assign wire_8592 = lut_tile_6_2_chanxy_out[21];
    assign wire_8594 = lut_tile_6_2_chanxy_out[22];
    assign wire_8596 = lut_tile_6_2_chanxy_out[23];
    assign wire_8598 = lut_tile_6_2_chanxy_out[24];
    assign wire_8600 = lut_tile_6_2_chanxy_out[25];
    assign wire_8602 = lut_tile_6_2_chanxy_out[26];
    assign wire_8604 = lut_tile_6_2_chanxy_out[27];
    assign wire_8606 = lut_tile_6_2_chanxy_out[28];
    assign wire_8608 = lut_tile_6_2_chanxy_out[29];
    assign wire_11341 = lut_tile_6_2_chanxy_out[30];
    assign wire_11343 = lut_tile_6_2_chanxy_out[31];
    assign wire_11345 = lut_tile_6_2_chanxy_out[32];
    assign wire_11347 = lut_tile_6_2_chanxy_out[33];
    assign wire_11349 = lut_tile_6_2_chanxy_out[34];
    assign wire_11351 = lut_tile_6_2_chanxy_out[35];
    assign wire_11353 = lut_tile_6_2_chanxy_out[36];
    assign wire_11355 = lut_tile_6_2_chanxy_out[37];
    assign wire_11357 = lut_tile_6_2_chanxy_out[38];
    assign wire_11359 = lut_tile_6_2_chanxy_out[39];
    assign wire_11361 = lut_tile_6_2_chanxy_out[40];
    assign wire_11363 = lut_tile_6_2_chanxy_out[41];
    assign wire_11365 = lut_tile_6_2_chanxy_out[42];
    assign wire_11367 = lut_tile_6_2_chanxy_out[43];
    assign wire_11369 = lut_tile_6_2_chanxy_out[44];
    assign wire_11430 = lut_tile_6_2_chanxy_out[45];
    assign wire_11432 = lut_tile_6_2_chanxy_out[46];
    assign wire_11434 = lut_tile_6_2_chanxy_out[47];
    assign wire_11436 = lut_tile_6_2_chanxy_out[48];
    assign wire_11438 = lut_tile_6_2_chanxy_out[49];
    assign wire_11440 = lut_tile_6_2_chanxy_out[50];
    assign wire_11442 = lut_tile_6_2_chanxy_out[51];
    assign wire_11444 = lut_tile_6_2_chanxy_out[52];
    assign wire_11446 = lut_tile_6_2_chanxy_out[53];
    assign wire_11448 = lut_tile_6_2_chanxy_out[54];
    assign wire_11450 = lut_tile_6_2_chanxy_out[55];
    assign wire_11452 = lut_tile_6_2_chanxy_out[56];
    assign wire_11454 = lut_tile_6_2_chanxy_out[57];
    assign wire_11456 = lut_tile_6_2_chanxy_out[58];
    assign wire_11458 = lut_tile_6_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_3_chanxy_in = {wire_11728, wire_8251, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8078, wire_2319, wire_11726, wire_8279, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8086, wire_2319, wire_11724, wire_8277, wire_8185, wire_8184, wire_8145, wire_8144, wire_8105, wire_8104, wire_8094, wire_2319, wire_11722, wire_8275, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8102, wire_1809, wire_11720, wire_8273, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8110, wire_1809, wire_11718, wire_8271, wire_8177, wire_8176, wire_8137, wire_8136, wire_8118, wire_8097, wire_8096, wire_1809, wire_11716, wire_8269, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8126, wire_2323, wire_1809, wire_11714, wire_8267, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8134, wire_2323, wire_1809, wire_11712, wire_8265, wire_8169, wire_8168, wire_8142, wire_8129, wire_8128, wire_8089, wire_8088, wire_2323, wire_1809, wire_11710, wire_8263, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8150, wire_2323, wire_1805, wire_11708, wire_8261, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8158, wire_2323, wire_1805, wire_11706, wire_8259, wire_8166, wire_8161, wire_8160, wire_8121, wire_8120, wire_8081, wire_8080, wire_2323, wire_1805, wire_11704, wire_8257, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8174, wire_2319, wire_1805, wire_11702, wire_8255, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8182, wire_2319, wire_1805, wire_11700, wire_8253, wire_8153, wire_8152, wire_8113, wire_8112, wire_8073, wire_8072, wire_8070, wire_2319, wire_1805, wire_11879, wire_8669, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8462, wire_2319, wire_11877, wire_8641, wire_8577, wire_8576, wire_8574, wire_8537, wire_8536, wire_8497, wire_8496, wire_2319, wire_11875, wire_8643, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8566, wire_2319, wire_11873, wire_8645, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8558, wire_1809, wire_11871, wire_8647, wire_8569, wire_8568, wire_8550, wire_8529, wire_8528, wire_8489, wire_8488, wire_1809, wire_11869, wire_8649, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8542, wire_1809, wire_11867, wire_8651, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8534, wire_2323, wire_1809, wire_11865, wire_8653, wire_8561, wire_8560, wire_8526, wire_8521, wire_8520, wire_8481, wire_8480, wire_2323, wire_1809, wire_11863, wire_8655, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8518, wire_2323, wire_1809, wire_11861, wire_8657, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8510, wire_2323, wire_1805, wire_11859, wire_8659, wire_8553, wire_8552, wire_8513, wire_8512, wire_8502, wire_8473, wire_8472, wire_2323, wire_1805, wire_11857, wire_8661, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8494, wire_2323, wire_1805, wire_11855, wire_8663, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8486, wire_2319, wire_1805, wire_11853, wire_8665, wire_8545, wire_8544, wire_8505, wire_8504, wire_8478, wire_8465, wire_8464, wire_2319, wire_1805, wire_11851, wire_8667, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8470, wire_2319, wire_1805, wire_11487, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11368, wire_8572, wire_1848, wire_11485, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11340, wire_8564, wire_1848, wire_11483, wire_11399, wire_11398, wire_11389, wire_11388, wire_11379, wire_11378, wire_11342, wire_8556, wire_1848, wire_11481, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11344, wire_8548, wire_1808, wire_11479, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11346, wire_8540, wire_1808, wire_11477, wire_11397, wire_11396, wire_11387, wire_11386, wire_11377, wire_11376, wire_11348, wire_8532, wire_1808, wire_11475, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11350, wire_8524, wire_1852, wire_1808, wire_11473, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11352, wire_8516, wire_1852, wire_1808, wire_11471, wire_11395, wire_11394, wire_11385, wire_11384, wire_11375, wire_11374, wire_11354, wire_8508, wire_1852, wire_1808, wire_11469, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11356, wire_8500, wire_1852, wire_1804, wire_11467, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11358, wire_8492, wire_1852, wire_1804, wire_11465, wire_11393, wire_11392, wire_11383, wire_11382, wire_11373, wire_11372, wire_11360, wire_8484, wire_1852, wire_1804, wire_11463, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11362, wire_8476, wire_1848, wire_1804, wire_11461, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11364, wire_8468, wire_1848, wire_1804, wire_11489, wire_11391, wire_11390, wire_11381, wire_11380, wire_11371, wire_11370, wire_11366, wire_8460, wire_1848, wire_1804, wire_11853, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11756, wire_8669, wire_1848, wire_11855, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11754, wire_8667, wire_1848, wire_11857, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11752, wire_8665, wire_1848, wire_11859, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11750, wire_8663, wire_1808, wire_11861, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11748, wire_8661, wire_1808, wire_11863, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11746, wire_8659, wire_1808, wire_11865, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11744, wire_8657, wire_1852, wire_1808, wire_11867, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11742, wire_8655, wire_1852, wire_1808, wire_11869, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11740, wire_8653, wire_1852, wire_1808, wire_11871, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11738, wire_8651, wire_1852, wire_1804, wire_11873, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11736, wire_8649, wire_1852, wire_1804, wire_11875, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11734, wire_8647, wire_1852, wire_1804, wire_11877, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11732, wire_8645, wire_1848, wire_1804, wire_11879, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11730, wire_8643, wire_1848, wire_1804, wire_11851, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11758, wire_8641, wire_1848, wire_1804};
    // CHNAXY TOTAL: 636
    assign wire_8463 = lut_tile_6_3_chanxy_out[0];
    assign wire_8471 = lut_tile_6_3_chanxy_out[1];
    assign wire_8479 = lut_tile_6_3_chanxy_out[2];
    assign wire_8487 = lut_tile_6_3_chanxy_out[3];
    assign wire_8495 = lut_tile_6_3_chanxy_out[4];
    assign wire_8503 = lut_tile_6_3_chanxy_out[5];
    assign wire_8511 = lut_tile_6_3_chanxy_out[6];
    assign wire_8519 = lut_tile_6_3_chanxy_out[7];
    assign wire_8527 = lut_tile_6_3_chanxy_out[8];
    assign wire_8535 = lut_tile_6_3_chanxy_out[9];
    assign wire_8543 = lut_tile_6_3_chanxy_out[10];
    assign wire_8551 = lut_tile_6_3_chanxy_out[11];
    assign wire_8559 = lut_tile_6_3_chanxy_out[12];
    assign wire_8567 = lut_tile_6_3_chanxy_out[13];
    assign wire_8575 = lut_tile_6_3_chanxy_out[14];
    assign wire_8610 = lut_tile_6_3_chanxy_out[15];
    assign wire_8612 = lut_tile_6_3_chanxy_out[16];
    assign wire_8614 = lut_tile_6_3_chanxy_out[17];
    assign wire_8616 = lut_tile_6_3_chanxy_out[18];
    assign wire_8618 = lut_tile_6_3_chanxy_out[19];
    assign wire_8620 = lut_tile_6_3_chanxy_out[20];
    assign wire_8622 = lut_tile_6_3_chanxy_out[21];
    assign wire_8624 = lut_tile_6_3_chanxy_out[22];
    assign wire_8626 = lut_tile_6_3_chanxy_out[23];
    assign wire_8628 = lut_tile_6_3_chanxy_out[24];
    assign wire_8630 = lut_tile_6_3_chanxy_out[25];
    assign wire_8632 = lut_tile_6_3_chanxy_out[26];
    assign wire_8634 = lut_tile_6_3_chanxy_out[27];
    assign wire_8636 = lut_tile_6_3_chanxy_out[28];
    assign wire_8638 = lut_tile_6_3_chanxy_out[29];
    assign wire_11731 = lut_tile_6_3_chanxy_out[30];
    assign wire_11733 = lut_tile_6_3_chanxy_out[31];
    assign wire_11735 = lut_tile_6_3_chanxy_out[32];
    assign wire_11737 = lut_tile_6_3_chanxy_out[33];
    assign wire_11739 = lut_tile_6_3_chanxy_out[34];
    assign wire_11741 = lut_tile_6_3_chanxy_out[35];
    assign wire_11743 = lut_tile_6_3_chanxy_out[36];
    assign wire_11745 = lut_tile_6_3_chanxy_out[37];
    assign wire_11747 = lut_tile_6_3_chanxy_out[38];
    assign wire_11749 = lut_tile_6_3_chanxy_out[39];
    assign wire_11751 = lut_tile_6_3_chanxy_out[40];
    assign wire_11753 = lut_tile_6_3_chanxy_out[41];
    assign wire_11755 = lut_tile_6_3_chanxy_out[42];
    assign wire_11757 = lut_tile_6_3_chanxy_out[43];
    assign wire_11759 = lut_tile_6_3_chanxy_out[44];
    assign wire_11820 = lut_tile_6_3_chanxy_out[45];
    assign wire_11822 = lut_tile_6_3_chanxy_out[46];
    assign wire_11824 = lut_tile_6_3_chanxy_out[47];
    assign wire_11826 = lut_tile_6_3_chanxy_out[48];
    assign wire_11828 = lut_tile_6_3_chanxy_out[49];
    assign wire_11830 = lut_tile_6_3_chanxy_out[50];
    assign wire_11832 = lut_tile_6_3_chanxy_out[51];
    assign wire_11834 = lut_tile_6_3_chanxy_out[52];
    assign wire_11836 = lut_tile_6_3_chanxy_out[53];
    assign wire_11838 = lut_tile_6_3_chanxy_out[54];
    assign wire_11840 = lut_tile_6_3_chanxy_out[55];
    assign wire_11842 = lut_tile_6_3_chanxy_out[56];
    assign wire_11844 = lut_tile_6_3_chanxy_out[57];
    assign wire_11846 = lut_tile_6_3_chanxy_out[58];
    assign wire_11848 = lut_tile_6_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_4_chanxy_in = {wire_12118, wire_8281, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8080, wire_2835, wire_12116, wire_8309, wire_8219, wire_8218, wire_8209, wire_8208, wire_8199, wire_8198, wire_8088, wire_2835, wire_12114, wire_8307, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8096, wire_2835, wire_12112, wire_8305, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8104, wire_2325, wire_12110, wire_8303, wire_8217, wire_8216, wire_8207, wire_8206, wire_8197, wire_8196, wire_8112, wire_2325, wire_12108, wire_8301, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8120, wire_2325, wire_12106, wire_8299, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8128, wire_2839, wire_2325, wire_12104, wire_8297, wire_8215, wire_8214, wire_8205, wire_8204, wire_8195, wire_8194, wire_8136, wire_2839, wire_2325, wire_12102, wire_8295, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8144, wire_2839, wire_2325, wire_12100, wire_8293, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8152, wire_2839, wire_2321, wire_12098, wire_8291, wire_8213, wire_8212, wire_8203, wire_8202, wire_8193, wire_8192, wire_8160, wire_2839, wire_2321, wire_12096, wire_8289, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8168, wire_2839, wire_2321, wire_12094, wire_8287, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8176, wire_2835, wire_2321, wire_12092, wire_8285, wire_8211, wire_8210, wire_8201, wire_8200, wire_8191, wire_8190, wire_8184, wire_2835, wire_2321, wire_12090, wire_8283, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8072, wire_2835, wire_2321, wire_12269, wire_8699, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8464, wire_2835, wire_12267, wire_8671, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8576, wire_2835, wire_12265, wire_8673, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8568, wire_2835, wire_12263, wire_8675, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8560, wire_2325, wire_12261, wire_8677, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8552, wire_2325, wire_12259, wire_8679, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8544, wire_2325, wire_12257, wire_8681, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8536, wire_2839, wire_2325, wire_12255, wire_8683, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8528, wire_2839, wire_2325, wire_12253, wire_8685, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8520, wire_2839, wire_2325, wire_12251, wire_8687, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8512, wire_2839, wire_2321, wire_12249, wire_8689, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8504, wire_2839, wire_2321, wire_12247, wire_8691, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8496, wire_2839, wire_2321, wire_12245, wire_8693, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8488, wire_2835, wire_2321, wire_12243, wire_8695, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8480, wire_2835, wire_2321, wire_12241, wire_8697, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8472, wire_2835, wire_2321, wire_11877, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11758, wire_8574, wire_2364, wire_11875, wire_11789, wire_11788, wire_11779, wire_11778, wire_11769, wire_11768, wire_11730, wire_8566, wire_2364, wire_11873, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11732, wire_8558, wire_2364, wire_11871, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11734, wire_8550, wire_2324, wire_11869, wire_11787, wire_11786, wire_11777, wire_11776, wire_11767, wire_11766, wire_11736, wire_8542, wire_2324, wire_11867, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11738, wire_8534, wire_2324, wire_11865, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11740, wire_8526, wire_2368, wire_2324, wire_11863, wire_11785, wire_11784, wire_11775, wire_11774, wire_11765, wire_11764, wire_11742, wire_8518, wire_2368, wire_2324, wire_11861, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11744, wire_8510, wire_2368, wire_2324, wire_11859, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11746, wire_8502, wire_2368, wire_2320, wire_11857, wire_11783, wire_11782, wire_11773, wire_11772, wire_11763, wire_11762, wire_11748, wire_8494, wire_2368, wire_2320, wire_11855, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11750, wire_8486, wire_2368, wire_2320, wire_11853, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11752, wire_8478, wire_2364, wire_2320, wire_11851, wire_11781, wire_11780, wire_11771, wire_11770, wire_11761, wire_11760, wire_11754, wire_8470, wire_2364, wire_2320, wire_11879, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11756, wire_8462, wire_2364, wire_2320, wire_12243, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12146, wire_8699, wire_2364, wire_12245, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12144, wire_8697, wire_2364, wire_12247, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12142, wire_8695, wire_2364, wire_12249, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12140, wire_8693, wire_2324, wire_12251, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12138, wire_8691, wire_2324, wire_12253, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12136, wire_8689, wire_2324, wire_12255, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12134, wire_8687, wire_2368, wire_2324, wire_12257, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12132, wire_8685, wire_2368, wire_2324, wire_12259, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12130, wire_8683, wire_2368, wire_2324, wire_12261, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12128, wire_8681, wire_2368, wire_2320, wire_12263, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12126, wire_8679, wire_2368, wire_2320, wire_12265, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12124, wire_8677, wire_2368, wire_2320, wire_12267, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12122, wire_8675, wire_2364, wire_2320, wire_12269, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12120, wire_8673, wire_2364, wire_2320, wire_12241, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12148, wire_8671, wire_2364, wire_2320};
    // CHNAXY TOTAL: 636
    assign wire_8465 = lut_tile_6_4_chanxy_out[0];
    assign wire_8473 = lut_tile_6_4_chanxy_out[1];
    assign wire_8481 = lut_tile_6_4_chanxy_out[2];
    assign wire_8489 = lut_tile_6_4_chanxy_out[3];
    assign wire_8497 = lut_tile_6_4_chanxy_out[4];
    assign wire_8505 = lut_tile_6_4_chanxy_out[5];
    assign wire_8513 = lut_tile_6_4_chanxy_out[6];
    assign wire_8521 = lut_tile_6_4_chanxy_out[7];
    assign wire_8529 = lut_tile_6_4_chanxy_out[8];
    assign wire_8537 = lut_tile_6_4_chanxy_out[9];
    assign wire_8545 = lut_tile_6_4_chanxy_out[10];
    assign wire_8553 = lut_tile_6_4_chanxy_out[11];
    assign wire_8561 = lut_tile_6_4_chanxy_out[12];
    assign wire_8569 = lut_tile_6_4_chanxy_out[13];
    assign wire_8577 = lut_tile_6_4_chanxy_out[14];
    assign wire_8640 = lut_tile_6_4_chanxy_out[15];
    assign wire_8642 = lut_tile_6_4_chanxy_out[16];
    assign wire_8644 = lut_tile_6_4_chanxy_out[17];
    assign wire_8646 = lut_tile_6_4_chanxy_out[18];
    assign wire_8648 = lut_tile_6_4_chanxy_out[19];
    assign wire_8650 = lut_tile_6_4_chanxy_out[20];
    assign wire_8652 = lut_tile_6_4_chanxy_out[21];
    assign wire_8654 = lut_tile_6_4_chanxy_out[22];
    assign wire_8656 = lut_tile_6_4_chanxy_out[23];
    assign wire_8658 = lut_tile_6_4_chanxy_out[24];
    assign wire_8660 = lut_tile_6_4_chanxy_out[25];
    assign wire_8662 = lut_tile_6_4_chanxy_out[26];
    assign wire_8664 = lut_tile_6_4_chanxy_out[27];
    assign wire_8666 = lut_tile_6_4_chanxy_out[28];
    assign wire_8668 = lut_tile_6_4_chanxy_out[29];
    assign wire_12121 = lut_tile_6_4_chanxy_out[30];
    assign wire_12123 = lut_tile_6_4_chanxy_out[31];
    assign wire_12125 = lut_tile_6_4_chanxy_out[32];
    assign wire_12127 = lut_tile_6_4_chanxy_out[33];
    assign wire_12129 = lut_tile_6_4_chanxy_out[34];
    assign wire_12131 = lut_tile_6_4_chanxy_out[35];
    assign wire_12133 = lut_tile_6_4_chanxy_out[36];
    assign wire_12135 = lut_tile_6_4_chanxy_out[37];
    assign wire_12137 = lut_tile_6_4_chanxy_out[38];
    assign wire_12139 = lut_tile_6_4_chanxy_out[39];
    assign wire_12141 = lut_tile_6_4_chanxy_out[40];
    assign wire_12143 = lut_tile_6_4_chanxy_out[41];
    assign wire_12145 = lut_tile_6_4_chanxy_out[42];
    assign wire_12147 = lut_tile_6_4_chanxy_out[43];
    assign wire_12149 = lut_tile_6_4_chanxy_out[44];
    assign wire_12210 = lut_tile_6_4_chanxy_out[45];
    assign wire_12212 = lut_tile_6_4_chanxy_out[46];
    assign wire_12214 = lut_tile_6_4_chanxy_out[47];
    assign wire_12216 = lut_tile_6_4_chanxy_out[48];
    assign wire_12218 = lut_tile_6_4_chanxy_out[49];
    assign wire_12220 = lut_tile_6_4_chanxy_out[50];
    assign wire_12222 = lut_tile_6_4_chanxy_out[51];
    assign wire_12224 = lut_tile_6_4_chanxy_out[52];
    assign wire_12226 = lut_tile_6_4_chanxy_out[53];
    assign wire_12228 = lut_tile_6_4_chanxy_out[54];
    assign wire_12230 = lut_tile_6_4_chanxy_out[55];
    assign wire_12232 = lut_tile_6_4_chanxy_out[56];
    assign wire_12234 = lut_tile_6_4_chanxy_out[57];
    assign wire_12236 = lut_tile_6_4_chanxy_out[58];
    assign wire_12238 = lut_tile_6_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_5_chanxy_in = {wire_12508, wire_8311, wire_8249, wire_8248, wire_8239, wire_8238, wire_8229, wire_8228, wire_8192, wire_3351, wire_12506, wire_8339, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8194, wire_3351, wire_12504, wire_8337, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8196, wire_3351, wire_12502, wire_8335, wire_8247, wire_8246, wire_8237, wire_8236, wire_8227, wire_8226, wire_8198, wire_2841, wire_12500, wire_8333, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8200, wire_2841, wire_12498, wire_8331, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8202, wire_2841, wire_12496, wire_8329, wire_8245, wire_8244, wire_8235, wire_8234, wire_8225, wire_8224, wire_8204, wire_3355, wire_2841, wire_12494, wire_8327, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8206, wire_3355, wire_2841, wire_12492, wire_8325, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8208, wire_3355, wire_2841, wire_12490, wire_8323, wire_8243, wire_8242, wire_8233, wire_8232, wire_8223, wire_8222, wire_8210, wire_3355, wire_2837, wire_12488, wire_8321, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8212, wire_3355, wire_2837, wire_12486, wire_8319, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8214, wire_3355, wire_2837, wire_12484, wire_8317, wire_8241, wire_8240, wire_8231, wire_8230, wire_8221, wire_8220, wire_8216, wire_3351, wire_2837, wire_12482, wire_8315, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8218, wire_3351, wire_2837, wire_12480, wire_8313, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8190, wire_3351, wire_2837, wire_12659, wire_8729, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8580, wire_3351, wire_12657, wire_8701, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8608, wire_3351, wire_12655, wire_8703, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8606, wire_3351, wire_12653, wire_8705, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8604, wire_2841, wire_12651, wire_8707, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8602, wire_2841, wire_12649, wire_8709, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8600, wire_2841, wire_12647, wire_8711, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8598, wire_3355, wire_2841, wire_12645, wire_8713, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8596, wire_3355, wire_2841, wire_12643, wire_8715, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8594, wire_3355, wire_2841, wire_12641, wire_8717, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8592, wire_3355, wire_2837, wire_12639, wire_8719, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8590, wire_3355, wire_2837, wire_12637, wire_8721, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8588, wire_3355, wire_2837, wire_12635, wire_8723, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8586, wire_3351, wire_2837, wire_12633, wire_8725, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8584, wire_3351, wire_2837, wire_12631, wire_8727, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8582, wire_3351, wire_2837, wire_12267, wire_12179, wire_12178, wire_12169, wire_12168, wire_12159, wire_12158, wire_12148, wire_8576, wire_2880, wire_12265, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12120, wire_8568, wire_2880, wire_12263, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12122, wire_8560, wire_2880, wire_12261, wire_12177, wire_12176, wire_12167, wire_12166, wire_12157, wire_12156, wire_12124, wire_8552, wire_2840, wire_12259, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12126, wire_8544, wire_2840, wire_12257, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12128, wire_8536, wire_2840, wire_12255, wire_12175, wire_12174, wire_12165, wire_12164, wire_12155, wire_12154, wire_12130, wire_8528, wire_2884, wire_2840, wire_12253, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12132, wire_8520, wire_2884, wire_2840, wire_12251, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12134, wire_8512, wire_2884, wire_2840, wire_12249, wire_12173, wire_12172, wire_12163, wire_12162, wire_12153, wire_12152, wire_12136, wire_8504, wire_2884, wire_2836, wire_12247, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12138, wire_8496, wire_2884, wire_2836, wire_12245, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12140, wire_8488, wire_2884, wire_2836, wire_12243, wire_12171, wire_12170, wire_12161, wire_12160, wire_12151, wire_12150, wire_12142, wire_8480, wire_2880, wire_2836, wire_12241, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12144, wire_8472, wire_2880, wire_2836, wire_12269, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12146, wire_8464, wire_2880, wire_2836, wire_12633, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12536, wire_8729, wire_2880, wire_12635, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12534, wire_8727, wire_2880, wire_12637, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12532, wire_8725, wire_2880, wire_12639, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12530, wire_8723, wire_2840, wire_12641, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12528, wire_8721, wire_2840, wire_12643, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12526, wire_8719, wire_2840, wire_12645, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12524, wire_8717, wire_2884, wire_2840, wire_12647, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12522, wire_8715, wire_2884, wire_2840, wire_12649, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12520, wire_8713, wire_2884, wire_2840, wire_12651, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12518, wire_8711, wire_2884, wire_2836, wire_12653, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12516, wire_8709, wire_2884, wire_2836, wire_12655, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12514, wire_8707, wire_2884, wire_2836, wire_12657, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12512, wire_8705, wire_2880, wire_2836, wire_12659, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12510, wire_8703, wire_2880, wire_2836, wire_12631, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12538, wire_8701, wire_2880, wire_2836};
    // CHNAXY TOTAL: 636
    assign wire_8581 = lut_tile_6_5_chanxy_out[0];
    assign wire_8583 = lut_tile_6_5_chanxy_out[1];
    assign wire_8585 = lut_tile_6_5_chanxy_out[2];
    assign wire_8587 = lut_tile_6_5_chanxy_out[3];
    assign wire_8589 = lut_tile_6_5_chanxy_out[4];
    assign wire_8591 = lut_tile_6_5_chanxy_out[5];
    assign wire_8593 = lut_tile_6_5_chanxy_out[6];
    assign wire_8595 = lut_tile_6_5_chanxy_out[7];
    assign wire_8597 = lut_tile_6_5_chanxy_out[8];
    assign wire_8599 = lut_tile_6_5_chanxy_out[9];
    assign wire_8601 = lut_tile_6_5_chanxy_out[10];
    assign wire_8603 = lut_tile_6_5_chanxy_out[11];
    assign wire_8605 = lut_tile_6_5_chanxy_out[12];
    assign wire_8607 = lut_tile_6_5_chanxy_out[13];
    assign wire_8609 = lut_tile_6_5_chanxy_out[14];
    assign wire_8670 = lut_tile_6_5_chanxy_out[15];
    assign wire_8672 = lut_tile_6_5_chanxy_out[16];
    assign wire_8674 = lut_tile_6_5_chanxy_out[17];
    assign wire_8676 = lut_tile_6_5_chanxy_out[18];
    assign wire_8678 = lut_tile_6_5_chanxy_out[19];
    assign wire_8680 = lut_tile_6_5_chanxy_out[20];
    assign wire_8682 = lut_tile_6_5_chanxy_out[21];
    assign wire_8684 = lut_tile_6_5_chanxy_out[22];
    assign wire_8686 = lut_tile_6_5_chanxy_out[23];
    assign wire_8688 = lut_tile_6_5_chanxy_out[24];
    assign wire_8690 = lut_tile_6_5_chanxy_out[25];
    assign wire_8692 = lut_tile_6_5_chanxy_out[26];
    assign wire_8694 = lut_tile_6_5_chanxy_out[27];
    assign wire_8696 = lut_tile_6_5_chanxy_out[28];
    assign wire_8698 = lut_tile_6_5_chanxy_out[29];
    assign wire_12511 = lut_tile_6_5_chanxy_out[30];
    assign wire_12513 = lut_tile_6_5_chanxy_out[31];
    assign wire_12515 = lut_tile_6_5_chanxy_out[32];
    assign wire_12517 = lut_tile_6_5_chanxy_out[33];
    assign wire_12519 = lut_tile_6_5_chanxy_out[34];
    assign wire_12521 = lut_tile_6_5_chanxy_out[35];
    assign wire_12523 = lut_tile_6_5_chanxy_out[36];
    assign wire_12525 = lut_tile_6_5_chanxy_out[37];
    assign wire_12527 = lut_tile_6_5_chanxy_out[38];
    assign wire_12529 = lut_tile_6_5_chanxy_out[39];
    assign wire_12531 = lut_tile_6_5_chanxy_out[40];
    assign wire_12533 = lut_tile_6_5_chanxy_out[41];
    assign wire_12535 = lut_tile_6_5_chanxy_out[42];
    assign wire_12537 = lut_tile_6_5_chanxy_out[43];
    assign wire_12539 = lut_tile_6_5_chanxy_out[44];
    assign wire_12600 = lut_tile_6_5_chanxy_out[45];
    assign wire_12602 = lut_tile_6_5_chanxy_out[46];
    assign wire_12604 = lut_tile_6_5_chanxy_out[47];
    assign wire_12606 = lut_tile_6_5_chanxy_out[48];
    assign wire_12608 = lut_tile_6_5_chanxy_out[49];
    assign wire_12610 = lut_tile_6_5_chanxy_out[50];
    assign wire_12612 = lut_tile_6_5_chanxy_out[51];
    assign wire_12614 = lut_tile_6_5_chanxy_out[52];
    assign wire_12616 = lut_tile_6_5_chanxy_out[53];
    assign wire_12618 = lut_tile_6_5_chanxy_out[54];
    assign wire_12620 = lut_tile_6_5_chanxy_out[55];
    assign wire_12622 = lut_tile_6_5_chanxy_out[56];
    assign wire_12624 = lut_tile_6_5_chanxy_out[57];
    assign wire_12626 = lut_tile_6_5_chanxy_out[58];
    assign wire_12628 = lut_tile_6_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_6_chanxy_in = {wire_12898, wire_8341, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8222, wire_3867, wire_12896, wire_8369, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8224, wire_3867, wire_12894, wire_8367, wire_8279, wire_8278, wire_8269, wire_8268, wire_8259, wire_8258, wire_8226, wire_3867, wire_12892, wire_8365, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8228, wire_3357, wire_12890, wire_8363, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8230, wire_3357, wire_12888, wire_8361, wire_8277, wire_8276, wire_8267, wire_8266, wire_8257, wire_8256, wire_8232, wire_3357, wire_12886, wire_8359, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8234, wire_3871, wire_3357, wire_12884, wire_8357, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8236, wire_3871, wire_3357, wire_12882, wire_8355, wire_8275, wire_8274, wire_8265, wire_8264, wire_8255, wire_8254, wire_8238, wire_3871, wire_3357, wire_12880, wire_8353, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8240, wire_3871, wire_3353, wire_12878, wire_8351, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8242, wire_3871, wire_3353, wire_12876, wire_8349, wire_8273, wire_8272, wire_8263, wire_8262, wire_8253, wire_8252, wire_8244, wire_3871, wire_3353, wire_12874, wire_8347, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8246, wire_3867, wire_3353, wire_12872, wire_8345, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8248, wire_3867, wire_3353, wire_12870, wire_8343, wire_8271, wire_8270, wire_8261, wire_8260, wire_8251, wire_8250, wire_8220, wire_3867, wire_3353, wire_13049, wire_8759, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8610, wire_3867, wire_13047, wire_8731, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8638, wire_3867, wire_13045, wire_8733, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8636, wire_3867, wire_13043, wire_8735, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8634, wire_3357, wire_13041, wire_8737, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8632, wire_3357, wire_13039, wire_8739, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8630, wire_3357, wire_13037, wire_8741, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8628, wire_3871, wire_3357, wire_13035, wire_8743, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8626, wire_3871, wire_3357, wire_13033, wire_8745, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8624, wire_3871, wire_3357, wire_13031, wire_8747, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8622, wire_3871, wire_3353, wire_13029, wire_8749, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8620, wire_3871, wire_3353, wire_13027, wire_8751, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8618, wire_3871, wire_3353, wire_13025, wire_8753, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8616, wire_3867, wire_3353, wire_13023, wire_8755, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8614, wire_3867, wire_3353, wire_13021, wire_8757, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8612, wire_3867, wire_3353, wire_12657, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12538, wire_8608, wire_3396, wire_12655, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12510, wire_8606, wire_3396, wire_12653, wire_12569, wire_12568, wire_12559, wire_12558, wire_12549, wire_12548, wire_12512, wire_8604, wire_3396, wire_12651, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12514, wire_8602, wire_3356, wire_12649, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12516, wire_8600, wire_3356, wire_12647, wire_12567, wire_12566, wire_12557, wire_12556, wire_12547, wire_12546, wire_12518, wire_8598, wire_3356, wire_12645, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12520, wire_8596, wire_3400, wire_3356, wire_12643, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12522, wire_8594, wire_3400, wire_3356, wire_12641, wire_12565, wire_12564, wire_12555, wire_12554, wire_12545, wire_12544, wire_12524, wire_8592, wire_3400, wire_3356, wire_12639, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12526, wire_8590, wire_3400, wire_3352, wire_12637, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12528, wire_8588, wire_3400, wire_3352, wire_12635, wire_12563, wire_12562, wire_12553, wire_12552, wire_12543, wire_12542, wire_12530, wire_8586, wire_3400, wire_3352, wire_12633, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12532, wire_8584, wire_3396, wire_3352, wire_12631, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12534, wire_8582, wire_3396, wire_3352, wire_12659, wire_12561, wire_12560, wire_12551, wire_12550, wire_12541, wire_12540, wire_12536, wire_8580, wire_3396, wire_3352, wire_13023, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12926, wire_8759, wire_3396, wire_13025, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12924, wire_8757, wire_3396, wire_13027, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12922, wire_8755, wire_3396, wire_13029, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12920, wire_8753, wire_3356, wire_13031, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12918, wire_8751, wire_3356, wire_13033, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12916, wire_8749, wire_3356, wire_13035, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12914, wire_8747, wire_3400, wire_3356, wire_13037, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12912, wire_8745, wire_3400, wire_3356, wire_13039, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12910, wire_8743, wire_3400, wire_3356, wire_13041, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12908, wire_8741, wire_3400, wire_3352, wire_13043, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12906, wire_8739, wire_3400, wire_3352, wire_13045, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12904, wire_8737, wire_3400, wire_3352, wire_13047, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12902, wire_8735, wire_3396, wire_3352, wire_13049, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12900, wire_8733, wire_3396, wire_3352, wire_13021, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12928, wire_8731, wire_3396, wire_3352};
    // CHNAXY TOTAL: 636
    assign wire_8611 = lut_tile_6_6_chanxy_out[0];
    assign wire_8613 = lut_tile_6_6_chanxy_out[1];
    assign wire_8615 = lut_tile_6_6_chanxy_out[2];
    assign wire_8617 = lut_tile_6_6_chanxy_out[3];
    assign wire_8619 = lut_tile_6_6_chanxy_out[4];
    assign wire_8621 = lut_tile_6_6_chanxy_out[5];
    assign wire_8623 = lut_tile_6_6_chanxy_out[6];
    assign wire_8625 = lut_tile_6_6_chanxy_out[7];
    assign wire_8627 = lut_tile_6_6_chanxy_out[8];
    assign wire_8629 = lut_tile_6_6_chanxy_out[9];
    assign wire_8631 = lut_tile_6_6_chanxy_out[10];
    assign wire_8633 = lut_tile_6_6_chanxy_out[11];
    assign wire_8635 = lut_tile_6_6_chanxy_out[12];
    assign wire_8637 = lut_tile_6_6_chanxy_out[13];
    assign wire_8639 = lut_tile_6_6_chanxy_out[14];
    assign wire_8700 = lut_tile_6_6_chanxy_out[15];
    assign wire_8702 = lut_tile_6_6_chanxy_out[16];
    assign wire_8704 = lut_tile_6_6_chanxy_out[17];
    assign wire_8706 = lut_tile_6_6_chanxy_out[18];
    assign wire_8708 = lut_tile_6_6_chanxy_out[19];
    assign wire_8710 = lut_tile_6_6_chanxy_out[20];
    assign wire_8712 = lut_tile_6_6_chanxy_out[21];
    assign wire_8714 = lut_tile_6_6_chanxy_out[22];
    assign wire_8716 = lut_tile_6_6_chanxy_out[23];
    assign wire_8718 = lut_tile_6_6_chanxy_out[24];
    assign wire_8720 = lut_tile_6_6_chanxy_out[25];
    assign wire_8722 = lut_tile_6_6_chanxy_out[26];
    assign wire_8724 = lut_tile_6_6_chanxy_out[27];
    assign wire_8726 = lut_tile_6_6_chanxy_out[28];
    assign wire_8728 = lut_tile_6_6_chanxy_out[29];
    assign wire_12901 = lut_tile_6_6_chanxy_out[30];
    assign wire_12903 = lut_tile_6_6_chanxy_out[31];
    assign wire_12905 = lut_tile_6_6_chanxy_out[32];
    assign wire_12907 = lut_tile_6_6_chanxy_out[33];
    assign wire_12909 = lut_tile_6_6_chanxy_out[34];
    assign wire_12911 = lut_tile_6_6_chanxy_out[35];
    assign wire_12913 = lut_tile_6_6_chanxy_out[36];
    assign wire_12915 = lut_tile_6_6_chanxy_out[37];
    assign wire_12917 = lut_tile_6_6_chanxy_out[38];
    assign wire_12919 = lut_tile_6_6_chanxy_out[39];
    assign wire_12921 = lut_tile_6_6_chanxy_out[40];
    assign wire_12923 = lut_tile_6_6_chanxy_out[41];
    assign wire_12925 = lut_tile_6_6_chanxy_out[42];
    assign wire_12927 = lut_tile_6_6_chanxy_out[43];
    assign wire_12929 = lut_tile_6_6_chanxy_out[44];
    assign wire_12990 = lut_tile_6_6_chanxy_out[45];
    assign wire_12992 = lut_tile_6_6_chanxy_out[46];
    assign wire_12994 = lut_tile_6_6_chanxy_out[47];
    assign wire_12996 = lut_tile_6_6_chanxy_out[48];
    assign wire_12998 = lut_tile_6_6_chanxy_out[49];
    assign wire_13000 = lut_tile_6_6_chanxy_out[50];
    assign wire_13002 = lut_tile_6_6_chanxy_out[51];
    assign wire_13004 = lut_tile_6_6_chanxy_out[52];
    assign wire_13006 = lut_tile_6_6_chanxy_out[53];
    assign wire_13008 = lut_tile_6_6_chanxy_out[54];
    assign wire_13010 = lut_tile_6_6_chanxy_out[55];
    assign wire_13012 = lut_tile_6_6_chanxy_out[56];
    assign wire_13014 = lut_tile_6_6_chanxy_out[57];
    assign wire_13016 = lut_tile_6_6_chanxy_out[58];
    assign wire_13018 = lut_tile_6_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_7_chanxy_in = {wire_13288, wire_8371, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8252, wire_4383, wire_13286, wire_8399, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8254, wire_4383, wire_13284, wire_8397, wire_8309, wire_8308, wire_8299, wire_8298, wire_8289, wire_8288, wire_8256, wire_4383, wire_13282, wire_8395, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8258, wire_3873, wire_13280, wire_8393, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8260, wire_3873, wire_13278, wire_8391, wire_8307, wire_8306, wire_8297, wire_8296, wire_8287, wire_8286, wire_8262, wire_3873, wire_13276, wire_8389, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8264, wire_4387, wire_3873, wire_13274, wire_8387, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8266, wire_4387, wire_3873, wire_13272, wire_8385, wire_8305, wire_8304, wire_8295, wire_8294, wire_8285, wire_8284, wire_8268, wire_4387, wire_3873, wire_13270, wire_8383, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8270, wire_4387, wire_3869, wire_13268, wire_8381, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8272, wire_4387, wire_3869, wire_13266, wire_8379, wire_8303, wire_8302, wire_8293, wire_8292, wire_8283, wire_8282, wire_8274, wire_4387, wire_3869, wire_13264, wire_8377, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8276, wire_4383, wire_3869, wire_13262, wire_8375, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8278, wire_4383, wire_3869, wire_13260, wire_8373, wire_8301, wire_8300, wire_8291, wire_8290, wire_8281, wire_8280, wire_8250, wire_4383, wire_3869, wire_13439, wire_8789, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8640, wire_4383, wire_13437, wire_8761, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8668, wire_4383, wire_13435, wire_8763, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8666, wire_4383, wire_13433, wire_8765, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8664, wire_3873, wire_13431, wire_8767, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8662, wire_3873, wire_13429, wire_8769, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8660, wire_3873, wire_13427, wire_8771, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8658, wire_4387, wire_3873, wire_13425, wire_8773, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8656, wire_4387, wire_3873, wire_13423, wire_8775, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8654, wire_4387, wire_3873, wire_13421, wire_8777, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8652, wire_4387, wire_3869, wire_13419, wire_8779, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8650, wire_4387, wire_3869, wire_13417, wire_8781, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8648, wire_4387, wire_3869, wire_13415, wire_8783, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8646, wire_4383, wire_3869, wire_13413, wire_8785, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8644, wire_4383, wire_3869, wire_13411, wire_8787, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8642, wire_4383, wire_3869, wire_13047, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12928, wire_8638, wire_3912, wire_13045, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12900, wire_8636, wire_3912, wire_13043, wire_12959, wire_12958, wire_12949, wire_12948, wire_12939, wire_12938, wire_12902, wire_8634, wire_3912, wire_13041, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12904, wire_8632, wire_3872, wire_13039, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12906, wire_8630, wire_3872, wire_13037, wire_12957, wire_12956, wire_12947, wire_12946, wire_12937, wire_12936, wire_12908, wire_8628, wire_3872, wire_13035, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12910, wire_8626, wire_3916, wire_3872, wire_13033, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12912, wire_8624, wire_3916, wire_3872, wire_13031, wire_12955, wire_12954, wire_12945, wire_12944, wire_12935, wire_12934, wire_12914, wire_8622, wire_3916, wire_3872, wire_13029, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12916, wire_8620, wire_3916, wire_3868, wire_13027, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12918, wire_8618, wire_3916, wire_3868, wire_13025, wire_12953, wire_12952, wire_12943, wire_12942, wire_12933, wire_12932, wire_12920, wire_8616, wire_3916, wire_3868, wire_13023, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12922, wire_8614, wire_3912, wire_3868, wire_13021, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12924, wire_8612, wire_3912, wire_3868, wire_13049, wire_12951, wire_12950, wire_12941, wire_12940, wire_12931, wire_12930, wire_12926, wire_8610, wire_3912, wire_3868, wire_13413, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13316, wire_8789, wire_3912, wire_13415, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13314, wire_8787, wire_3912, wire_13417, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13312, wire_8785, wire_3912, wire_13419, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13310, wire_8783, wire_3872, wire_13421, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13308, wire_8781, wire_3872, wire_13423, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13306, wire_8779, wire_3872, wire_13425, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13304, wire_8777, wire_3916, wire_3872, wire_13427, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13302, wire_8775, wire_3916, wire_3872, wire_13429, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13300, wire_8773, wire_3916, wire_3872, wire_13431, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13298, wire_8771, wire_3916, wire_3868, wire_13433, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13296, wire_8769, wire_3916, wire_3868, wire_13435, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13294, wire_8767, wire_3916, wire_3868, wire_13437, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13292, wire_8765, wire_3912, wire_3868, wire_13439, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13290, wire_8763, wire_3912, wire_3868, wire_13411, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13318, wire_8761, wire_3912, wire_3868};
    // CHNAXY TOTAL: 636
    assign wire_8641 = lut_tile_6_7_chanxy_out[0];
    assign wire_8643 = lut_tile_6_7_chanxy_out[1];
    assign wire_8645 = lut_tile_6_7_chanxy_out[2];
    assign wire_8647 = lut_tile_6_7_chanxy_out[3];
    assign wire_8649 = lut_tile_6_7_chanxy_out[4];
    assign wire_8651 = lut_tile_6_7_chanxy_out[5];
    assign wire_8653 = lut_tile_6_7_chanxy_out[6];
    assign wire_8655 = lut_tile_6_7_chanxy_out[7];
    assign wire_8657 = lut_tile_6_7_chanxy_out[8];
    assign wire_8659 = lut_tile_6_7_chanxy_out[9];
    assign wire_8661 = lut_tile_6_7_chanxy_out[10];
    assign wire_8663 = lut_tile_6_7_chanxy_out[11];
    assign wire_8665 = lut_tile_6_7_chanxy_out[12];
    assign wire_8667 = lut_tile_6_7_chanxy_out[13];
    assign wire_8669 = lut_tile_6_7_chanxy_out[14];
    assign wire_8730 = lut_tile_6_7_chanxy_out[15];
    assign wire_8732 = lut_tile_6_7_chanxy_out[16];
    assign wire_8734 = lut_tile_6_7_chanxy_out[17];
    assign wire_8736 = lut_tile_6_7_chanxy_out[18];
    assign wire_8738 = lut_tile_6_7_chanxy_out[19];
    assign wire_8740 = lut_tile_6_7_chanxy_out[20];
    assign wire_8742 = lut_tile_6_7_chanxy_out[21];
    assign wire_8744 = lut_tile_6_7_chanxy_out[22];
    assign wire_8746 = lut_tile_6_7_chanxy_out[23];
    assign wire_8748 = lut_tile_6_7_chanxy_out[24];
    assign wire_8750 = lut_tile_6_7_chanxy_out[25];
    assign wire_8752 = lut_tile_6_7_chanxy_out[26];
    assign wire_8754 = lut_tile_6_7_chanxy_out[27];
    assign wire_8756 = lut_tile_6_7_chanxy_out[28];
    assign wire_8758 = lut_tile_6_7_chanxy_out[29];
    assign wire_13291 = lut_tile_6_7_chanxy_out[30];
    assign wire_13293 = lut_tile_6_7_chanxy_out[31];
    assign wire_13295 = lut_tile_6_7_chanxy_out[32];
    assign wire_13297 = lut_tile_6_7_chanxy_out[33];
    assign wire_13299 = lut_tile_6_7_chanxy_out[34];
    assign wire_13301 = lut_tile_6_7_chanxy_out[35];
    assign wire_13303 = lut_tile_6_7_chanxy_out[36];
    assign wire_13305 = lut_tile_6_7_chanxy_out[37];
    assign wire_13307 = lut_tile_6_7_chanxy_out[38];
    assign wire_13309 = lut_tile_6_7_chanxy_out[39];
    assign wire_13311 = lut_tile_6_7_chanxy_out[40];
    assign wire_13313 = lut_tile_6_7_chanxy_out[41];
    assign wire_13315 = lut_tile_6_7_chanxy_out[42];
    assign wire_13317 = lut_tile_6_7_chanxy_out[43];
    assign wire_13319 = lut_tile_6_7_chanxy_out[44];
    assign wire_13380 = lut_tile_6_7_chanxy_out[45];
    assign wire_13382 = lut_tile_6_7_chanxy_out[46];
    assign wire_13384 = lut_tile_6_7_chanxy_out[47];
    assign wire_13386 = lut_tile_6_7_chanxy_out[48];
    assign wire_13388 = lut_tile_6_7_chanxy_out[49];
    assign wire_13390 = lut_tile_6_7_chanxy_out[50];
    assign wire_13392 = lut_tile_6_7_chanxy_out[51];
    assign wire_13394 = lut_tile_6_7_chanxy_out[52];
    assign wire_13396 = lut_tile_6_7_chanxy_out[53];
    assign wire_13398 = lut_tile_6_7_chanxy_out[54];
    assign wire_13400 = lut_tile_6_7_chanxy_out[55];
    assign wire_13402 = lut_tile_6_7_chanxy_out[56];
    assign wire_13404 = lut_tile_6_7_chanxy_out[57];
    assign wire_13406 = lut_tile_6_7_chanxy_out[58];
    assign wire_13408 = lut_tile_6_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_8_chanxy_in = {wire_13678, wire_8401, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8282, wire_4899, wire_13676, wire_8429, wire_8339, wire_8338, wire_8329, wire_8328, wire_8319, wire_8318, wire_8284, wire_4899, wire_13674, wire_8427, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8286, wire_4899, wire_13672, wire_8425, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8288, wire_4389, wire_13670, wire_8423, wire_8337, wire_8336, wire_8327, wire_8326, wire_8317, wire_8316, wire_8290, wire_4389, wire_13668, wire_8421, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8292, wire_4389, wire_13666, wire_8419, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8294, wire_4903, wire_4389, wire_13664, wire_8417, wire_8335, wire_8334, wire_8325, wire_8324, wire_8315, wire_8314, wire_8296, wire_4903, wire_4389, wire_13662, wire_8415, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8298, wire_4903, wire_4389, wire_13660, wire_8413, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8300, wire_4903, wire_4385, wire_13658, wire_8411, wire_8333, wire_8332, wire_8323, wire_8322, wire_8313, wire_8312, wire_8302, wire_4903, wire_4385, wire_13656, wire_8409, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8304, wire_4903, wire_4385, wire_13654, wire_8407, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8306, wire_4899, wire_4385, wire_13652, wire_8405, wire_8331, wire_8330, wire_8321, wire_8320, wire_8311, wire_8310, wire_8308, wire_4899, wire_4385, wire_13650, wire_8403, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8280, wire_4899, wire_4385, wire_13829, wire_8819, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8670, wire_4899, wire_13827, wire_8791, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8698, wire_4899, wire_13825, wire_8793, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8696, wire_4899, wire_13823, wire_8795, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8694, wire_4389, wire_13821, wire_8797, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8692, wire_4389, wire_13819, wire_8799, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8690, wire_4389, wire_13817, wire_8801, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8688, wire_4903, wire_4389, wire_13815, wire_8803, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8686, wire_4903, wire_4389, wire_13813, wire_8805, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8684, wire_4903, wire_4389, wire_13811, wire_8807, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8682, wire_4903, wire_4385, wire_13809, wire_8809, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8680, wire_4903, wire_4385, wire_13807, wire_8811, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8678, wire_4903, wire_4385, wire_13805, wire_8813, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8676, wire_4899, wire_4385, wire_13803, wire_8815, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8674, wire_4899, wire_4385, wire_13801, wire_8817, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8672, wire_4899, wire_4385, wire_13437, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13318, wire_8668, wire_4428, wire_13435, wire_13349, wire_13348, wire_13339, wire_13338, wire_13329, wire_13328, wire_13290, wire_8666, wire_4428, wire_13433, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13292, wire_8664, wire_4428, wire_13431, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13294, wire_8662, wire_4388, wire_13429, wire_13347, wire_13346, wire_13337, wire_13336, wire_13327, wire_13326, wire_13296, wire_8660, wire_4388, wire_13427, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13298, wire_8658, wire_4388, wire_13425, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13300, wire_8656, wire_4432, wire_4388, wire_13423, wire_13345, wire_13344, wire_13335, wire_13334, wire_13325, wire_13324, wire_13302, wire_8654, wire_4432, wire_4388, wire_13421, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13304, wire_8652, wire_4432, wire_4388, wire_13419, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13306, wire_8650, wire_4432, wire_4384, wire_13417, wire_13343, wire_13342, wire_13333, wire_13332, wire_13323, wire_13322, wire_13308, wire_8648, wire_4432, wire_4384, wire_13415, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13310, wire_8646, wire_4432, wire_4384, wire_13413, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13312, wire_8644, wire_4428, wire_4384, wire_13411, wire_13341, wire_13340, wire_13331, wire_13330, wire_13321, wire_13320, wire_13314, wire_8642, wire_4428, wire_4384, wire_13439, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13316, wire_8640, wire_4428, wire_4384, wire_13803, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13706, wire_8819, wire_4428, wire_13805, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13704, wire_8817, wire_4428, wire_13807, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13702, wire_8815, wire_4428, wire_13809, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13700, wire_8813, wire_4388, wire_13811, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13698, wire_8811, wire_4388, wire_13813, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13696, wire_8809, wire_4388, wire_13815, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13694, wire_8807, wire_4432, wire_4388, wire_13817, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13692, wire_8805, wire_4432, wire_4388, wire_13819, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13690, wire_8803, wire_4432, wire_4388, wire_13821, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13688, wire_8801, wire_4432, wire_4384, wire_13823, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13686, wire_8799, wire_4432, wire_4384, wire_13825, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13684, wire_8797, wire_4432, wire_4384, wire_13827, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13682, wire_8795, wire_4428, wire_4384, wire_13829, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13680, wire_8793, wire_4428, wire_4384, wire_13801, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13708, wire_8791, wire_4428, wire_4384};
    // CHNAXY TOTAL: 636
    assign wire_8671 = lut_tile_6_8_chanxy_out[0];
    assign wire_8673 = lut_tile_6_8_chanxy_out[1];
    assign wire_8675 = lut_tile_6_8_chanxy_out[2];
    assign wire_8677 = lut_tile_6_8_chanxy_out[3];
    assign wire_8679 = lut_tile_6_8_chanxy_out[4];
    assign wire_8681 = lut_tile_6_8_chanxy_out[5];
    assign wire_8683 = lut_tile_6_8_chanxy_out[6];
    assign wire_8685 = lut_tile_6_8_chanxy_out[7];
    assign wire_8687 = lut_tile_6_8_chanxy_out[8];
    assign wire_8689 = lut_tile_6_8_chanxy_out[9];
    assign wire_8691 = lut_tile_6_8_chanxy_out[10];
    assign wire_8693 = lut_tile_6_8_chanxy_out[11];
    assign wire_8695 = lut_tile_6_8_chanxy_out[12];
    assign wire_8697 = lut_tile_6_8_chanxy_out[13];
    assign wire_8699 = lut_tile_6_8_chanxy_out[14];
    assign wire_8760 = lut_tile_6_8_chanxy_out[15];
    assign wire_8762 = lut_tile_6_8_chanxy_out[16];
    assign wire_8764 = lut_tile_6_8_chanxy_out[17];
    assign wire_8766 = lut_tile_6_8_chanxy_out[18];
    assign wire_8768 = lut_tile_6_8_chanxy_out[19];
    assign wire_8770 = lut_tile_6_8_chanxy_out[20];
    assign wire_8772 = lut_tile_6_8_chanxy_out[21];
    assign wire_8774 = lut_tile_6_8_chanxy_out[22];
    assign wire_8776 = lut_tile_6_8_chanxy_out[23];
    assign wire_8778 = lut_tile_6_8_chanxy_out[24];
    assign wire_8780 = lut_tile_6_8_chanxy_out[25];
    assign wire_8782 = lut_tile_6_8_chanxy_out[26];
    assign wire_8784 = lut_tile_6_8_chanxy_out[27];
    assign wire_8786 = lut_tile_6_8_chanxy_out[28];
    assign wire_8788 = lut_tile_6_8_chanxy_out[29];
    assign wire_13681 = lut_tile_6_8_chanxy_out[30];
    assign wire_13683 = lut_tile_6_8_chanxy_out[31];
    assign wire_13685 = lut_tile_6_8_chanxy_out[32];
    assign wire_13687 = lut_tile_6_8_chanxy_out[33];
    assign wire_13689 = lut_tile_6_8_chanxy_out[34];
    assign wire_13691 = lut_tile_6_8_chanxy_out[35];
    assign wire_13693 = lut_tile_6_8_chanxy_out[36];
    assign wire_13695 = lut_tile_6_8_chanxy_out[37];
    assign wire_13697 = lut_tile_6_8_chanxy_out[38];
    assign wire_13699 = lut_tile_6_8_chanxy_out[39];
    assign wire_13701 = lut_tile_6_8_chanxy_out[40];
    assign wire_13703 = lut_tile_6_8_chanxy_out[41];
    assign wire_13705 = lut_tile_6_8_chanxy_out[42];
    assign wire_13707 = lut_tile_6_8_chanxy_out[43];
    assign wire_13709 = lut_tile_6_8_chanxy_out[44];
    assign wire_13770 = lut_tile_6_8_chanxy_out[45];
    assign wire_13772 = lut_tile_6_8_chanxy_out[46];
    assign wire_13774 = lut_tile_6_8_chanxy_out[47];
    assign wire_13776 = lut_tile_6_8_chanxy_out[48];
    assign wire_13778 = lut_tile_6_8_chanxy_out[49];
    assign wire_13780 = lut_tile_6_8_chanxy_out[50];
    assign wire_13782 = lut_tile_6_8_chanxy_out[51];
    assign wire_13784 = lut_tile_6_8_chanxy_out[52];
    assign wire_13786 = lut_tile_6_8_chanxy_out[53];
    assign wire_13788 = lut_tile_6_8_chanxy_out[54];
    assign wire_13790 = lut_tile_6_8_chanxy_out[55];
    assign wire_13792 = lut_tile_6_8_chanxy_out[56];
    assign wire_13794 = lut_tile_6_8_chanxy_out[57];
    assign wire_13796 = lut_tile_6_8_chanxy_out[58];
    assign wire_13798 = lut_tile_6_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_9_chanxy_in = {wire_14068, wire_8431, wire_8369, wire_8368, wire_8359, wire_8358, wire_8349, wire_8348, wire_8312, wire_5415, wire_14066, wire_8459, wire_8429, wire_8428, wire_8419, wire_8418, wire_8409, wire_8408, wire_8314, wire_5415, wire_14064, wire_8457, wire_8399, wire_8398, wire_8389, wire_8388, wire_8379, wire_8378, wire_8316, wire_5415, wire_14062, wire_8455, wire_8367, wire_8366, wire_8357, wire_8356, wire_8347, wire_8346, wire_8318, wire_4905, wire_14060, wire_8453, wire_8427, wire_8426, wire_8417, wire_8416, wire_8407, wire_8406, wire_8320, wire_4905, wire_14058, wire_8451, wire_8397, wire_8396, wire_8387, wire_8386, wire_8377, wire_8376, wire_8322, wire_4905, wire_14056, wire_8449, wire_8365, wire_8364, wire_8355, wire_8354, wire_8345, wire_8344, wire_8324, wire_5419, wire_4905, wire_14054, wire_8447, wire_8425, wire_8424, wire_8415, wire_8414, wire_8405, wire_8404, wire_8326, wire_5419, wire_4905, wire_14052, wire_8445, wire_8395, wire_8394, wire_8385, wire_8384, wire_8375, wire_8374, wire_8328, wire_5419, wire_4905, wire_14050, wire_8443, wire_8363, wire_8362, wire_8353, wire_8352, wire_8343, wire_8342, wire_8330, wire_5419, wire_4901, wire_14048, wire_8441, wire_8423, wire_8422, wire_8413, wire_8412, wire_8403, wire_8402, wire_8332, wire_5419, wire_4901, wire_14046, wire_8439, wire_8393, wire_8392, wire_8383, wire_8382, wire_8373, wire_8372, wire_8334, wire_5419, wire_4901, wire_14044, wire_8437, wire_8361, wire_8360, wire_8351, wire_8350, wire_8341, wire_8340, wire_8336, wire_5415, wire_4901, wire_14042, wire_8435, wire_8421, wire_8420, wire_8411, wire_8410, wire_8401, wire_8400, wire_8338, wire_5415, wire_4901, wire_14040, wire_8433, wire_8391, wire_8390, wire_8381, wire_8380, wire_8371, wire_8370, wire_8310, wire_5415, wire_4901, wire_14219, wire_8849, wire_8819, wire_8818, wire_8809, wire_8808, wire_8799, wire_8798, wire_8700, wire_5415, wire_14217, wire_8821, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8728, wire_5415, wire_14215, wire_8823, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8726, wire_5415, wire_14213, wire_8825, wire_8817, wire_8816, wire_8807, wire_8806, wire_8797, wire_8796, wire_8724, wire_4905, wire_14211, wire_8827, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8722, wire_4905, wire_14209, wire_8829, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8720, wire_4905, wire_14207, wire_8831, wire_8815, wire_8814, wire_8805, wire_8804, wire_8795, wire_8794, wire_8718, wire_5419, wire_4905, wire_14205, wire_8833, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8716, wire_5419, wire_4905, wire_14203, wire_8835, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8714, wire_5419, wire_4905, wire_14201, wire_8837, wire_8813, wire_8812, wire_8803, wire_8802, wire_8793, wire_8792, wire_8712, wire_5419, wire_4901, wire_14199, wire_8839, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8710, wire_5419, wire_4901, wire_14197, wire_8841, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8708, wire_5419, wire_4901, wire_14195, wire_8843, wire_8811, wire_8810, wire_8801, wire_8800, wire_8791, wire_8790, wire_8706, wire_5415, wire_4901, wire_14193, wire_8845, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8704, wire_5415, wire_4901, wire_14191, wire_8847, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8702, wire_5415, wire_4901, wire_13827, wire_13739, wire_13738, wire_13729, wire_13728, wire_13719, wire_13718, wire_13708, wire_8698, wire_4944, wire_13825, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13680, wire_8696, wire_4944, wire_13823, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13682, wire_8694, wire_4944, wire_13821, wire_13737, wire_13736, wire_13727, wire_13726, wire_13717, wire_13716, wire_13684, wire_8692, wire_4904, wire_13819, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13686, wire_8690, wire_4904, wire_13817, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13688, wire_8688, wire_4904, wire_13815, wire_13735, wire_13734, wire_13725, wire_13724, wire_13715, wire_13714, wire_13690, wire_8686, wire_4948, wire_4904, wire_13813, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13692, wire_8684, wire_4948, wire_4904, wire_13811, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13694, wire_8682, wire_4948, wire_4904, wire_13809, wire_13733, wire_13732, wire_13723, wire_13722, wire_13713, wire_13712, wire_13696, wire_8680, wire_4948, wire_4900, wire_13807, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13698, wire_8678, wire_4948, wire_4900, wire_13805, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13700, wire_8676, wire_4948, wire_4900, wire_13803, wire_13731, wire_13730, wire_13721, wire_13720, wire_13711, wire_13710, wire_13702, wire_8674, wire_4944, wire_4900, wire_13801, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13704, wire_8672, wire_4944, wire_4900, wire_13829, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13706, wire_8670, wire_4944, wire_4900, wire_14193, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14096, wire_8849, wire_4944, wire_14195, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14094, wire_8847, wire_4944, wire_14197, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14092, wire_8845, wire_4944, wire_14199, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14090, wire_8843, wire_4904, wire_14201, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14088, wire_8841, wire_4904, wire_14203, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14086, wire_8839, wire_4904, wire_14205, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14084, wire_8837, wire_4948, wire_4904, wire_14207, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14082, wire_8835, wire_4948, wire_4904, wire_14209, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14080, wire_8833, wire_4948, wire_4904, wire_14211, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14078, wire_8831, wire_4948, wire_4900, wire_14213, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14076, wire_8829, wire_4948, wire_4900, wire_14215, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14074, wire_8827, wire_4948, wire_4900, wire_14217, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14072, wire_8825, wire_4944, wire_4900, wire_14219, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14070, wire_8823, wire_4944, wire_4900, wire_14191, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14098, wire_8821, wire_4944, wire_4900};
    // CHNAXY TOTAL: 636
    assign wire_8701 = lut_tile_6_9_chanxy_out[0];
    assign wire_8703 = lut_tile_6_9_chanxy_out[1];
    assign wire_8705 = lut_tile_6_9_chanxy_out[2];
    assign wire_8707 = lut_tile_6_9_chanxy_out[3];
    assign wire_8709 = lut_tile_6_9_chanxy_out[4];
    assign wire_8711 = lut_tile_6_9_chanxy_out[5];
    assign wire_8713 = lut_tile_6_9_chanxy_out[6];
    assign wire_8715 = lut_tile_6_9_chanxy_out[7];
    assign wire_8717 = lut_tile_6_9_chanxy_out[8];
    assign wire_8719 = lut_tile_6_9_chanxy_out[9];
    assign wire_8721 = lut_tile_6_9_chanxy_out[10];
    assign wire_8723 = lut_tile_6_9_chanxy_out[11];
    assign wire_8725 = lut_tile_6_9_chanxy_out[12];
    assign wire_8727 = lut_tile_6_9_chanxy_out[13];
    assign wire_8729 = lut_tile_6_9_chanxy_out[14];
    assign wire_8790 = lut_tile_6_9_chanxy_out[15];
    assign wire_8792 = lut_tile_6_9_chanxy_out[16];
    assign wire_8794 = lut_tile_6_9_chanxy_out[17];
    assign wire_8796 = lut_tile_6_9_chanxy_out[18];
    assign wire_8798 = lut_tile_6_9_chanxy_out[19];
    assign wire_8800 = lut_tile_6_9_chanxy_out[20];
    assign wire_8802 = lut_tile_6_9_chanxy_out[21];
    assign wire_8804 = lut_tile_6_9_chanxy_out[22];
    assign wire_8806 = lut_tile_6_9_chanxy_out[23];
    assign wire_8808 = lut_tile_6_9_chanxy_out[24];
    assign wire_8810 = lut_tile_6_9_chanxy_out[25];
    assign wire_8812 = lut_tile_6_9_chanxy_out[26];
    assign wire_8814 = lut_tile_6_9_chanxy_out[27];
    assign wire_8816 = lut_tile_6_9_chanxy_out[28];
    assign wire_8818 = lut_tile_6_9_chanxy_out[29];
    assign wire_14071 = lut_tile_6_9_chanxy_out[30];
    assign wire_14073 = lut_tile_6_9_chanxy_out[31];
    assign wire_14075 = lut_tile_6_9_chanxy_out[32];
    assign wire_14077 = lut_tile_6_9_chanxy_out[33];
    assign wire_14079 = lut_tile_6_9_chanxy_out[34];
    assign wire_14081 = lut_tile_6_9_chanxy_out[35];
    assign wire_14083 = lut_tile_6_9_chanxy_out[36];
    assign wire_14085 = lut_tile_6_9_chanxy_out[37];
    assign wire_14087 = lut_tile_6_9_chanxy_out[38];
    assign wire_14089 = lut_tile_6_9_chanxy_out[39];
    assign wire_14091 = lut_tile_6_9_chanxy_out[40];
    assign wire_14093 = lut_tile_6_9_chanxy_out[41];
    assign wire_14095 = lut_tile_6_9_chanxy_out[42];
    assign wire_14097 = lut_tile_6_9_chanxy_out[43];
    assign wire_14099 = lut_tile_6_9_chanxy_out[44];
    assign wire_14160 = lut_tile_6_9_chanxy_out[45];
    assign wire_14162 = lut_tile_6_9_chanxy_out[46];
    assign wire_14164 = lut_tile_6_9_chanxy_out[47];
    assign wire_14166 = lut_tile_6_9_chanxy_out[48];
    assign wire_14168 = lut_tile_6_9_chanxy_out[49];
    assign wire_14170 = lut_tile_6_9_chanxy_out[50];
    assign wire_14172 = lut_tile_6_9_chanxy_out[51];
    assign wire_14174 = lut_tile_6_9_chanxy_out[52];
    assign wire_14176 = lut_tile_6_9_chanxy_out[53];
    assign wire_14178 = lut_tile_6_9_chanxy_out[54];
    assign wire_14180 = lut_tile_6_9_chanxy_out[55];
    assign wire_14182 = lut_tile_6_9_chanxy_out[56];
    assign wire_14184 = lut_tile_6_9_chanxy_out[57];
    assign wire_14186 = lut_tile_6_9_chanxy_out[58];
    assign wire_14188 = lut_tile_6_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_6_10_chanxy_in = {wire_14458, wire_8436, wire_8414, wire_8392, wire_8368, wire_5926, wire_5920, wire_5911, wire_5905, wire_14456, wire_8458, wire_8406, wire_8384, wire_8360, wire_5926, wire_5920, wire_5911, wire_5905, wire_14454, wire_8450, wire_8428, wire_8376, wire_8352, wire_5926, wire_5920, wire_5911, wire_5905, wire_14452, wire_8442, wire_8420, wire_8398, wire_8344, wire_5926, wire_5917, wire_5911, wire_5421, wire_14450, wire_8434, wire_8412, wire_8390, wire_8366, wire_5926, wire_5917, wire_5911, wire_5421, wire_14448, wire_8456, wire_8404, wire_8382, wire_8358, wire_5926, wire_5917, wire_5911, wire_5421, wire_14446, wire_8448, wire_8426, wire_8374, wire_8350, wire_5923, wire_5917, wire_5908, wire_5421, wire_14444, wire_8440, wire_8418, wire_8396, wire_8342, wire_5923, wire_5917, wire_5908, wire_5421, wire_14442, wire_8432, wire_8410, wire_8388, wire_8364, wire_5923, wire_5917, wire_5908, wire_5421, wire_14440, wire_8454, wire_8402, wire_8380, wire_8356, wire_5923, wire_5914, wire_5908, wire_5417, wire_14438, wire_8446, wire_8424, wire_8372, wire_8348, wire_5923, wire_5914, wire_5908, wire_5417, wire_14436, wire_8438, wire_8416, wire_8394, wire_8340, wire_5923, wire_5914, wire_5908, wire_5417, wire_14434, wire_8430, wire_8408, wire_8386, wire_8362, wire_5920, wire_5914, wire_5905, wire_5417, wire_14432, wire_8452, wire_8400, wire_8378, wire_8354, wire_5920, wire_5914, wire_5905, wire_5417, wire_14430, wire_8444, wire_8422, wire_8370, wire_8346, wire_5920, wire_5914, wire_5905, wire_5417, wire_14609, wire_8848, wire_8796, wire_8774, wire_8752, wire_5926, wire_5920, wire_5911, wire_5905, wire_14607, wire_8840, wire_8818, wire_8766, wire_8744, wire_5926, wire_5920, wire_5911, wire_5905, wire_14605, wire_8832, wire_8810, wire_8788, wire_8736, wire_5926, wire_5920, wire_5911, wire_5905, wire_14603, wire_8824, wire_8802, wire_8780, wire_8758, wire_5926, wire_5917, wire_5911, wire_5421, wire_14601, wire_8846, wire_8794, wire_8772, wire_8750, wire_5926, wire_5917, wire_5911, wire_5421, wire_14599, wire_8838, wire_8816, wire_8764, wire_8742, wire_5926, wire_5917, wire_5911, wire_5421, wire_14597, wire_8830, wire_8808, wire_8786, wire_8734, wire_5923, wire_5917, wire_5908, wire_5421, wire_14595, wire_8822, wire_8800, wire_8778, wire_8756, wire_5923, wire_5917, wire_5908, wire_5421, wire_14593, wire_8844, wire_8792, wire_8770, wire_8748, wire_5923, wire_5917, wire_5908, wire_5421, wire_14591, wire_8836, wire_8814, wire_8762, wire_8740, wire_5923, wire_5914, wire_5908, wire_5417, wire_14589, wire_8828, wire_8806, wire_8784, wire_8732, wire_5923, wire_5914, wire_5908, wire_5417, wire_14587, wire_8820, wire_8798, wire_8776, wire_8754, wire_5923, wire_5914, wire_5908, wire_5417, wire_14585, wire_8842, wire_8790, wire_8768, wire_8746, wire_5920, wire_5914, wire_5905, wire_5417, wire_14583, wire_8834, wire_8812, wire_8760, wire_8738, wire_5920, wire_5914, wire_5905, wire_5417, wire_14581, wire_8826, wire_8804, wire_8782, wire_8730, wire_5920, wire_5914, wire_5905, wire_5417, wire_14579, wire_14578, wire_14217, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14098, wire_8728, wire_5460, wire_14609, wire_14488, wire_14215, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14070, wire_8726, wire_5460, wire_14503, wire_14502, wire_14213, wire_14129, wire_14128, wire_14119, wire_14118, wire_14109, wire_14108, wire_14072, wire_8724, wire_5460, wire_14561, wire_14560, wire_14211, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14074, wire_8722, wire_5420, wire_14591, wire_14470, wire_14209, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14076, wire_8720, wire_5420, wire_14515, wire_14514, wire_14207, wire_14127, wire_14126, wire_14117, wire_14116, wire_14107, wire_14106, wire_14078, wire_8718, wire_5420, wire_14573, wire_14572, wire_14205, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14080, wire_8716, wire_5464, wire_5420, wire_14603, wire_14482, wire_14203, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14082, wire_8714, wire_5464, wire_5420, wire_14497, wire_14496, wire_14201, wire_14125, wire_14124, wire_14115, wire_14114, wire_14105, wire_14104, wire_14084, wire_8712, wire_5464, wire_5420, wire_14555, wire_14554, wire_5464, wire_14199, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14086, wire_8710, wire_5464, wire_5416, wire_14585, wire_14464, wire_5464, wire_14197, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14088, wire_8708, wire_5464, wire_5416, wire_14509, wire_14508, wire_5460, wire_14195, wire_14123, wire_14122, wire_14113, wire_14112, wire_14103, wire_14102, wire_14090, wire_8706, wire_5464, wire_5416, wire_14567, wire_14566, wire_5420, wire_14193, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14092, wire_8704, wire_5460, wire_5416, wire_14597, wire_14476, wire_5420, wire_14191, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14094, wire_8702, wire_5460, wire_5416, wire_14491, wire_14490, wire_5416, wire_14219, wire_14121, wire_14120, wire_14111, wire_14110, wire_14101, wire_14100, wire_14096, wire_8700, wire_5460, wire_5416, wire_14549, wire_14548, wire_14533, wire_14532, wire_14517, wire_14516, wire_14531, wire_14530, wire_14545, wire_14544, wire_14499, wire_14498, wire_14543, wire_14542, wire_14527, wire_14526, wire_14511, wire_14510, wire_14525, wire_14524, wire_5464, wire_14539, wire_14538, wire_5464, wire_14493, wire_14492, wire_5460, wire_14537, wire_14536, wire_5420, wire_14521, wire_14520, wire_5420, wire_14505, wire_14504, wire_5416, wire_14563, wire_14562, wire_14577, wire_14576, wire_14607, wire_14486, wire_14575, wire_14574, wire_14559, wire_14558, wire_14589, wire_14468, wire_14557, wire_14556, wire_14571, wire_14570, wire_14601, wire_14480, wire_14569, wire_14568, wire_5464, wire_14553, wire_14552, wire_5460, wire_14583, wire_14462, wire_5460, wire_14551, wire_14550, wire_5420, wire_14565, wire_14564, wire_5416, wire_14595, wire_14474, wire_5416, wire_14519, wire_14518, wire_14547, wire_14546, wire_14593, wire_14472, wire_14501, wire_14500, wire_14529, wire_14528, wire_14605, wire_14484, wire_14513, wire_14512, wire_14541, wire_14540, wire_14587, wire_14466, wire_14495, wire_14494, wire_5464, wire_14523, wire_14522, wire_5460, wire_14599, wire_14478, wire_5460, wire_14507, wire_14506, wire_5420, wire_14535, wire_14534, wire_5416, wire_14581, wire_14460, wire_5416};
    // CHNAXY TOTAL: 573
    assign wire_8731 = lut_tile_6_10_chanxy_out[0];
    assign wire_8733 = lut_tile_6_10_chanxy_out[1];
    assign wire_8735 = lut_tile_6_10_chanxy_out[2];
    assign wire_8737 = lut_tile_6_10_chanxy_out[3];
    assign wire_8739 = lut_tile_6_10_chanxy_out[4];
    assign wire_8741 = lut_tile_6_10_chanxy_out[5];
    assign wire_8743 = lut_tile_6_10_chanxy_out[6];
    assign wire_8745 = lut_tile_6_10_chanxy_out[7];
    assign wire_8747 = lut_tile_6_10_chanxy_out[8];
    assign wire_8749 = lut_tile_6_10_chanxy_out[9];
    assign wire_8751 = lut_tile_6_10_chanxy_out[10];
    assign wire_8753 = lut_tile_6_10_chanxy_out[11];
    assign wire_8755 = lut_tile_6_10_chanxy_out[12];
    assign wire_8757 = lut_tile_6_10_chanxy_out[13];
    assign wire_8759 = lut_tile_6_10_chanxy_out[14];
    assign wire_8761 = lut_tile_6_10_chanxy_out[15];
    assign wire_8763 = lut_tile_6_10_chanxy_out[16];
    assign wire_8765 = lut_tile_6_10_chanxy_out[17];
    assign wire_8767 = lut_tile_6_10_chanxy_out[18];
    assign wire_8769 = lut_tile_6_10_chanxy_out[19];
    assign wire_8771 = lut_tile_6_10_chanxy_out[20];
    assign wire_8773 = lut_tile_6_10_chanxy_out[21];
    assign wire_8775 = lut_tile_6_10_chanxy_out[22];
    assign wire_8777 = lut_tile_6_10_chanxy_out[23];
    assign wire_8779 = lut_tile_6_10_chanxy_out[24];
    assign wire_8781 = lut_tile_6_10_chanxy_out[25];
    assign wire_8783 = lut_tile_6_10_chanxy_out[26];
    assign wire_8785 = lut_tile_6_10_chanxy_out[27];
    assign wire_8787 = lut_tile_6_10_chanxy_out[28];
    assign wire_8789 = lut_tile_6_10_chanxy_out[29];
    assign wire_8791 = lut_tile_6_10_chanxy_out[30];
    assign wire_8793 = lut_tile_6_10_chanxy_out[31];
    assign wire_8795 = lut_tile_6_10_chanxy_out[32];
    assign wire_8797 = lut_tile_6_10_chanxy_out[33];
    assign wire_8799 = lut_tile_6_10_chanxy_out[34];
    assign wire_8801 = lut_tile_6_10_chanxy_out[35];
    assign wire_8803 = lut_tile_6_10_chanxy_out[36];
    assign wire_8805 = lut_tile_6_10_chanxy_out[37];
    assign wire_8807 = lut_tile_6_10_chanxy_out[38];
    assign wire_8809 = lut_tile_6_10_chanxy_out[39];
    assign wire_8811 = lut_tile_6_10_chanxy_out[40];
    assign wire_8813 = lut_tile_6_10_chanxy_out[41];
    assign wire_8815 = lut_tile_6_10_chanxy_out[42];
    assign wire_8817 = lut_tile_6_10_chanxy_out[43];
    assign wire_8819 = lut_tile_6_10_chanxy_out[44];
    assign wire_8820 = lut_tile_6_10_chanxy_out[45];
    assign wire_8821 = lut_tile_6_10_chanxy_out[46];
    assign wire_8822 = lut_tile_6_10_chanxy_out[47];
    assign wire_8823 = lut_tile_6_10_chanxy_out[48];
    assign wire_8824 = lut_tile_6_10_chanxy_out[49];
    assign wire_8825 = lut_tile_6_10_chanxy_out[50];
    assign wire_8826 = lut_tile_6_10_chanxy_out[51];
    assign wire_8827 = lut_tile_6_10_chanxy_out[52];
    assign wire_8828 = lut_tile_6_10_chanxy_out[53];
    assign wire_8829 = lut_tile_6_10_chanxy_out[54];
    assign wire_8830 = lut_tile_6_10_chanxy_out[55];
    assign wire_8831 = lut_tile_6_10_chanxy_out[56];
    assign wire_8832 = lut_tile_6_10_chanxy_out[57];
    assign wire_8833 = lut_tile_6_10_chanxy_out[58];
    assign wire_8834 = lut_tile_6_10_chanxy_out[59];
    assign wire_8835 = lut_tile_6_10_chanxy_out[60];
    assign wire_8836 = lut_tile_6_10_chanxy_out[61];
    assign wire_8837 = lut_tile_6_10_chanxy_out[62];
    assign wire_8838 = lut_tile_6_10_chanxy_out[63];
    assign wire_8839 = lut_tile_6_10_chanxy_out[64];
    assign wire_8840 = lut_tile_6_10_chanxy_out[65];
    assign wire_8841 = lut_tile_6_10_chanxy_out[66];
    assign wire_8842 = lut_tile_6_10_chanxy_out[67];
    assign wire_8843 = lut_tile_6_10_chanxy_out[68];
    assign wire_8844 = lut_tile_6_10_chanxy_out[69];
    assign wire_8845 = lut_tile_6_10_chanxy_out[70];
    assign wire_8846 = lut_tile_6_10_chanxy_out[71];
    assign wire_8847 = lut_tile_6_10_chanxy_out[72];
    assign wire_8848 = lut_tile_6_10_chanxy_out[73];
    assign wire_8849 = lut_tile_6_10_chanxy_out[74];
    assign wire_14461 = lut_tile_6_10_chanxy_out[75];
    assign wire_14463 = lut_tile_6_10_chanxy_out[76];
    assign wire_14465 = lut_tile_6_10_chanxy_out[77];
    assign wire_14467 = lut_tile_6_10_chanxy_out[78];
    assign wire_14469 = lut_tile_6_10_chanxy_out[79];
    assign wire_14471 = lut_tile_6_10_chanxy_out[80];
    assign wire_14473 = lut_tile_6_10_chanxy_out[81];
    assign wire_14475 = lut_tile_6_10_chanxy_out[82];
    assign wire_14477 = lut_tile_6_10_chanxy_out[83];
    assign wire_14479 = lut_tile_6_10_chanxy_out[84];
    assign wire_14481 = lut_tile_6_10_chanxy_out[85];
    assign wire_14483 = lut_tile_6_10_chanxy_out[86];
    assign wire_14485 = lut_tile_6_10_chanxy_out[87];
    assign wire_14487 = lut_tile_6_10_chanxy_out[88];
    assign wire_14489 = lut_tile_6_10_chanxy_out[89];
    assign wire_14550 = lut_tile_6_10_chanxy_out[90];
    assign wire_14552 = lut_tile_6_10_chanxy_out[91];
    assign wire_14554 = lut_tile_6_10_chanxy_out[92];
    assign wire_14556 = lut_tile_6_10_chanxy_out[93];
    assign wire_14558 = lut_tile_6_10_chanxy_out[94];
    assign wire_14560 = lut_tile_6_10_chanxy_out[95];
    assign wire_14562 = lut_tile_6_10_chanxy_out[96];
    assign wire_14564 = lut_tile_6_10_chanxy_out[97];
    assign wire_14566 = lut_tile_6_10_chanxy_out[98];
    assign wire_14568 = lut_tile_6_10_chanxy_out[99];
    assign wire_14570 = lut_tile_6_10_chanxy_out[100];
    assign wire_14572 = lut_tile_6_10_chanxy_out[101];
    assign wire_14574 = lut_tile_6_10_chanxy_out[102];
    assign wire_14576 = lut_tile_6_10_chanxy_out[103];
    assign wire_14578 = lut_tile_6_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_7_1_chanxy_in = {wire_10978, wire_8581, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_8474, wire_1329, wire_10976, wire_8609, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_8482, wire_1329, wire_10974, wire_8607, wire_8573, wire_8572, wire_8533, wire_8532, wire_8493, wire_8492, wire_8490, wire_1329, wire_10972, wire_8605, wire_8569, wire_8568, wire_8529, wire_8528, wire_8498, wire_8489, wire_8488, wire_819, wire_10970, wire_8603, wire_8567, wire_8566, wire_8527, wire_8526, wire_8506, wire_8487, wire_8486, wire_819, wire_10968, wire_8601, wire_8565, wire_8564, wire_8525, wire_8524, wire_8514, wire_8485, wire_8484, wire_819, wire_10966, wire_8599, wire_8561, wire_8560, wire_8522, wire_8521, wire_8520, wire_8481, wire_8480, wire_1333, wire_819, wire_10964, wire_8597, wire_8559, wire_8558, wire_8530, wire_8519, wire_8518, wire_8479, wire_8478, wire_1333, wire_819, wire_10962, wire_8595, wire_8557, wire_8556, wire_8538, wire_8517, wire_8516, wire_8477, wire_8476, wire_1333, wire_819, wire_10960, wire_8593, wire_8553, wire_8552, wire_8546, wire_8513, wire_8512, wire_8473, wire_8472, wire_1333, wire_815, wire_10958, wire_8591, wire_8554, wire_8551, wire_8550, wire_8511, wire_8510, wire_8471, wire_8470, wire_1333, wire_815, wire_10956, wire_8589, wire_8562, wire_8549, wire_8548, wire_8509, wire_8508, wire_8469, wire_8468, wire_1333, wire_815, wire_10954, wire_8587, wire_8570, wire_8545, wire_8544, wire_8505, wire_8504, wire_8465, wire_8464, wire_1329, wire_815, wire_10952, wire_8585, wire_8578, wire_8543, wire_8542, wire_8503, wire_8502, wire_8463, wire_8462, wire_1329, wire_815, wire_10950, wire_8583, wire_8541, wire_8540, wire_8501, wire_8500, wire_8466, wire_8461, wire_8460, wire_1329, wire_815, wire_11129, wire_8999, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8850, wire_1329, wire_11127, wire_8971, wire_8967, wire_8966, wire_8962, wire_8927, wire_8926, wire_8887, wire_8886, wire_1329, wire_11125, wire_8973, wire_8965, wire_8964, wire_8954, wire_8925, wire_8924, wire_8885, wire_8884, wire_1329, wire_11123, wire_8975, wire_8961, wire_8960, wire_8946, wire_8921, wire_8920, wire_8881, wire_8880, wire_819, wire_11121, wire_8977, wire_8959, wire_8958, wire_8938, wire_8919, wire_8918, wire_8879, wire_8878, wire_819, wire_11119, wire_8979, wire_8957, wire_8956, wire_8930, wire_8917, wire_8916, wire_8877, wire_8876, wire_819, wire_11117, wire_8981, wire_8953, wire_8952, wire_8922, wire_8913, wire_8912, wire_8873, wire_8872, wire_1333, wire_819, wire_11115, wire_8983, wire_8951, wire_8950, wire_8914, wire_8911, wire_8910, wire_8871, wire_8870, wire_1333, wire_819, wire_11113, wire_8985, wire_8949, wire_8948, wire_8909, wire_8908, wire_8906, wire_8869, wire_8868, wire_1333, wire_819, wire_11111, wire_8987, wire_8945, wire_8944, wire_8905, wire_8904, wire_8898, wire_8865, wire_8864, wire_1333, wire_815, wire_11109, wire_8989, wire_8943, wire_8942, wire_8903, wire_8902, wire_8890, wire_8863, wire_8862, wire_1333, wire_815, wire_11107, wire_8991, wire_8941, wire_8940, wire_8901, wire_8900, wire_8882, wire_8861, wire_8860, wire_1333, wire_815, wire_11105, wire_8993, wire_8937, wire_8936, wire_8897, wire_8896, wire_8874, wire_8857, wire_8856, wire_1329, wire_815, wire_11103, wire_8995, wire_8935, wire_8934, wire_8895, wire_8894, wire_8866, wire_8855, wire_8854, wire_1329, wire_815, wire_11101, wire_8997, wire_8933, wire_8932, wire_8893, wire_8892, wire_8858, wire_8853, wire_8852, wire_1329, wire_815, wire_10723, wire_10602, wire_10739, wire_10618, wire_10709, wire_10708, wire_11103, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11006, wire_8999, wire_858, wire_10693, wire_10692, wire_10679, wire_10678, wire_10649, wire_10648, wire_10663, wire_10662, wire_11105, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_11004, wire_8997, wire_858, wire_10737, wire_10616, wire_10707, wire_10706, wire_10633, wire_10632, wire_10677, wire_10676, wire_11107, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_11002, wire_8995, wire_858, wire_10647, wire_10646, wire_10735, wire_10614, wire_10721, wire_10600, wire_10691, wire_10690, wire_11109, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11000, wire_8993, wire_818, wire_10705, wire_10704, wire_10661, wire_10660, wire_10631, wire_10630, wire_10675, wire_10674, wire_11111, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_10998, wire_8991, wire_818, wire_10719, wire_10598, wire_10689, wire_10688, wire_10645, wire_10644, wire_10659, wire_10658, wire_11113, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10996, wire_8989, wire_818, wire_10629, wire_10628, wire_10717, wire_10596, wire_10733, wire_10612, wire_10703, wire_10702, wire_11115, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_10994, wire_8987, wire_862, wire_818, wire_10687, wire_10686, wire_10673, wire_10672, wire_10643, wire_10642, wire_10657, wire_10656, wire_11117, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_10992, wire_8985, wire_862, wire_818, wire_10731, wire_10610, wire_10701, wire_10700, wire_10627, wire_10626, wire_10671, wire_10670, wire_11119, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10990, wire_8983, wire_862, wire_818, wire_10641, wire_10640, wire_10729, wire_10608, wire_862, wire_10715, wire_10594, wire_862, wire_10685, wire_10684, wire_862, wire_11121, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_10988, wire_8981, wire_862, wire_814, wire_10699, wire_10698, wire_862, wire_10655, wire_10654, wire_862, wire_10625, wire_10624, wire_862, wire_10669, wire_10668, wire_858, wire_11123, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_10986, wire_8979, wire_862, wire_814, wire_10713, wire_10592, wire_858, wire_10683, wire_10682, wire_858, wire_10639, wire_10638, wire_858, wire_10653, wire_10652, wire_858, wire_11125, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_10984, wire_8977, wire_862, wire_814, wire_10623, wire_10622, wire_858, wire_10711, wire_10590, wire_818, wire_10727, wire_10606, wire_818, wire_10697, wire_10696, wire_818, wire_11127, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_10982, wire_8975, wire_858, wire_814, wire_10681, wire_10680, wire_818, wire_10667, wire_10666, wire_818, wire_10637, wire_10636, wire_818, wire_10651, wire_10650, wire_814, wire_11129, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_10980, wire_8973, wire_858, wire_814, wire_10725, wire_10604, wire_814, wire_10695, wire_10694, wire_814, wire_10621, wire_10620, wire_814, wire_10665, wire_10664, wire_814, wire_11101, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_11008, wire_8971, wire_858, wire_814, wire_10635, wire_10634, wire_814};
    // CHNAXY TOTAL: 621
    assign wire_8850 = lut_tile_7_1_chanxy_out[0];
    assign wire_8851 = lut_tile_7_1_chanxy_out[1];
    assign wire_8852 = lut_tile_7_1_chanxy_out[2];
    assign wire_8854 = lut_tile_7_1_chanxy_out[3];
    assign wire_8856 = lut_tile_7_1_chanxy_out[4];
    assign wire_8858 = lut_tile_7_1_chanxy_out[5];
    assign wire_8859 = lut_tile_7_1_chanxy_out[6];
    assign wire_8860 = lut_tile_7_1_chanxy_out[7];
    assign wire_8862 = lut_tile_7_1_chanxy_out[8];
    assign wire_8864 = lut_tile_7_1_chanxy_out[9];
    assign wire_8866 = lut_tile_7_1_chanxy_out[10];
    assign wire_8867 = lut_tile_7_1_chanxy_out[11];
    assign wire_8868 = lut_tile_7_1_chanxy_out[12];
    assign wire_8870 = lut_tile_7_1_chanxy_out[13];
    assign wire_8872 = lut_tile_7_1_chanxy_out[14];
    assign wire_8874 = lut_tile_7_1_chanxy_out[15];
    assign wire_8875 = lut_tile_7_1_chanxy_out[16];
    assign wire_8876 = lut_tile_7_1_chanxy_out[17];
    assign wire_8878 = lut_tile_7_1_chanxy_out[18];
    assign wire_8880 = lut_tile_7_1_chanxy_out[19];
    assign wire_8882 = lut_tile_7_1_chanxy_out[20];
    assign wire_8883 = lut_tile_7_1_chanxy_out[21];
    assign wire_8884 = lut_tile_7_1_chanxy_out[22];
    assign wire_8886 = lut_tile_7_1_chanxy_out[23];
    assign wire_8888 = lut_tile_7_1_chanxy_out[24];
    assign wire_8890 = lut_tile_7_1_chanxy_out[25];
    assign wire_8891 = lut_tile_7_1_chanxy_out[26];
    assign wire_8892 = lut_tile_7_1_chanxy_out[27];
    assign wire_8894 = lut_tile_7_1_chanxy_out[28];
    assign wire_8896 = lut_tile_7_1_chanxy_out[29];
    assign wire_8898 = lut_tile_7_1_chanxy_out[30];
    assign wire_8899 = lut_tile_7_1_chanxy_out[31];
    assign wire_8900 = lut_tile_7_1_chanxy_out[32];
    assign wire_8902 = lut_tile_7_1_chanxy_out[33];
    assign wire_8904 = lut_tile_7_1_chanxy_out[34];
    assign wire_8906 = lut_tile_7_1_chanxy_out[35];
    assign wire_8907 = lut_tile_7_1_chanxy_out[36];
    assign wire_8908 = lut_tile_7_1_chanxy_out[37];
    assign wire_8910 = lut_tile_7_1_chanxy_out[38];
    assign wire_8912 = lut_tile_7_1_chanxy_out[39];
    assign wire_8914 = lut_tile_7_1_chanxy_out[40];
    assign wire_8915 = lut_tile_7_1_chanxy_out[41];
    assign wire_8916 = lut_tile_7_1_chanxy_out[42];
    assign wire_8918 = lut_tile_7_1_chanxy_out[43];
    assign wire_8920 = lut_tile_7_1_chanxy_out[44];
    assign wire_8922 = lut_tile_7_1_chanxy_out[45];
    assign wire_8923 = lut_tile_7_1_chanxy_out[46];
    assign wire_8924 = lut_tile_7_1_chanxy_out[47];
    assign wire_8926 = lut_tile_7_1_chanxy_out[48];
    assign wire_8928 = lut_tile_7_1_chanxy_out[49];
    assign wire_8930 = lut_tile_7_1_chanxy_out[50];
    assign wire_8931 = lut_tile_7_1_chanxy_out[51];
    assign wire_8932 = lut_tile_7_1_chanxy_out[52];
    assign wire_8934 = lut_tile_7_1_chanxy_out[53];
    assign wire_8936 = lut_tile_7_1_chanxy_out[54];
    assign wire_8938 = lut_tile_7_1_chanxy_out[55];
    assign wire_8939 = lut_tile_7_1_chanxy_out[56];
    assign wire_8940 = lut_tile_7_1_chanxy_out[57];
    assign wire_8942 = lut_tile_7_1_chanxy_out[58];
    assign wire_8944 = lut_tile_7_1_chanxy_out[59];
    assign wire_8946 = lut_tile_7_1_chanxy_out[60];
    assign wire_8947 = lut_tile_7_1_chanxy_out[61];
    assign wire_8948 = lut_tile_7_1_chanxy_out[62];
    assign wire_8950 = lut_tile_7_1_chanxy_out[63];
    assign wire_8952 = lut_tile_7_1_chanxy_out[64];
    assign wire_8954 = lut_tile_7_1_chanxy_out[65];
    assign wire_8955 = lut_tile_7_1_chanxy_out[66];
    assign wire_8956 = lut_tile_7_1_chanxy_out[67];
    assign wire_8958 = lut_tile_7_1_chanxy_out[68];
    assign wire_8960 = lut_tile_7_1_chanxy_out[69];
    assign wire_8962 = lut_tile_7_1_chanxy_out[70];
    assign wire_8963 = lut_tile_7_1_chanxy_out[71];
    assign wire_8964 = lut_tile_7_1_chanxy_out[72];
    assign wire_8966 = lut_tile_7_1_chanxy_out[73];
    assign wire_8968 = lut_tile_7_1_chanxy_out[74];
    assign wire_10981 = lut_tile_7_1_chanxy_out[75];
    assign wire_10983 = lut_tile_7_1_chanxy_out[76];
    assign wire_10985 = lut_tile_7_1_chanxy_out[77];
    assign wire_10987 = lut_tile_7_1_chanxy_out[78];
    assign wire_10989 = lut_tile_7_1_chanxy_out[79];
    assign wire_10991 = lut_tile_7_1_chanxy_out[80];
    assign wire_10993 = lut_tile_7_1_chanxy_out[81];
    assign wire_10995 = lut_tile_7_1_chanxy_out[82];
    assign wire_10997 = lut_tile_7_1_chanxy_out[83];
    assign wire_10999 = lut_tile_7_1_chanxy_out[84];
    assign wire_11001 = lut_tile_7_1_chanxy_out[85];
    assign wire_11003 = lut_tile_7_1_chanxy_out[86];
    assign wire_11005 = lut_tile_7_1_chanxy_out[87];
    assign wire_11007 = lut_tile_7_1_chanxy_out[88];
    assign wire_11009 = lut_tile_7_1_chanxy_out[89];
    assign wire_11070 = lut_tile_7_1_chanxy_out[90];
    assign wire_11072 = lut_tile_7_1_chanxy_out[91];
    assign wire_11074 = lut_tile_7_1_chanxy_out[92];
    assign wire_11076 = lut_tile_7_1_chanxy_out[93];
    assign wire_11078 = lut_tile_7_1_chanxy_out[94];
    assign wire_11080 = lut_tile_7_1_chanxy_out[95];
    assign wire_11082 = lut_tile_7_1_chanxy_out[96];
    assign wire_11084 = lut_tile_7_1_chanxy_out[97];
    assign wire_11086 = lut_tile_7_1_chanxy_out[98];
    assign wire_11088 = lut_tile_7_1_chanxy_out[99];
    assign wire_11090 = lut_tile_7_1_chanxy_out[100];
    assign wire_11092 = lut_tile_7_1_chanxy_out[101];
    assign wire_11094 = lut_tile_7_1_chanxy_out[102];
    assign wire_11096 = lut_tile_7_1_chanxy_out[103];
    assign wire_11098 = lut_tile_7_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_7_2_chanxy_in = {wire_11368, wire_8611, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8468, wire_1845, wire_11366, wire_8639, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_8476, wire_1845, wire_11364, wire_8637, wire_8575, wire_8574, wire_8535, wire_8534, wire_8495, wire_8494, wire_8484, wire_1845, wire_11362, wire_8635, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8492, wire_1335, wire_11360, wire_8633, wire_8569, wire_8568, wire_8529, wire_8528, wire_8500, wire_8489, wire_8488, wire_1335, wire_11358, wire_8631, wire_8567, wire_8566, wire_8527, wire_8526, wire_8508, wire_8487, wire_8486, wire_1335, wire_11356, wire_8629, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8516, wire_1849, wire_1335, wire_11354, wire_8627, wire_8561, wire_8560, wire_8524, wire_8521, wire_8520, wire_8481, wire_8480, wire_1849, wire_1335, wire_11352, wire_8625, wire_8559, wire_8558, wire_8532, wire_8519, wire_8518, wire_8479, wire_8478, wire_1849, wire_1335, wire_11350, wire_8623, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8540, wire_1849, wire_1331, wire_11348, wire_8621, wire_8553, wire_8552, wire_8548, wire_8513, wire_8512, wire_8473, wire_8472, wire_1849, wire_1331, wire_11346, wire_8619, wire_8556, wire_8551, wire_8550, wire_8511, wire_8510, wire_8471, wire_8470, wire_1849, wire_1331, wire_11344, wire_8617, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8564, wire_1845, wire_1331, wire_11342, wire_8615, wire_8572, wire_8545, wire_8544, wire_8505, wire_8504, wire_8465, wire_8464, wire_1845, wire_1331, wire_11340, wire_8613, wire_8543, wire_8542, wire_8503, wire_8502, wire_8463, wire_8462, wire_8460, wire_1845, wire_1331, wire_11519, wire_9029, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8852, wire_1845, wire_11517, wire_9001, wire_8967, wire_8966, wire_8964, wire_8927, wire_8926, wire_8887, wire_8886, wire_1845, wire_11515, wire_9003, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8956, wire_1845, wire_11513, wire_9005, wire_8961, wire_8960, wire_8948, wire_8921, wire_8920, wire_8881, wire_8880, wire_1335, wire_11511, wire_9007, wire_8959, wire_8958, wire_8940, wire_8919, wire_8918, wire_8879, wire_8878, wire_1335, wire_11509, wire_9009, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8932, wire_1335, wire_11507, wire_9011, wire_8953, wire_8952, wire_8924, wire_8913, wire_8912, wire_8873, wire_8872, wire_1849, wire_1335, wire_11505, wire_9013, wire_8951, wire_8950, wire_8916, wire_8911, wire_8910, wire_8871, wire_8870, wire_1849, wire_1335, wire_11503, wire_9015, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8908, wire_1849, wire_1335, wire_11501, wire_9017, wire_8945, wire_8944, wire_8905, wire_8904, wire_8900, wire_8865, wire_8864, wire_1849, wire_1331, wire_11499, wire_9019, wire_8943, wire_8942, wire_8903, wire_8902, wire_8892, wire_8863, wire_8862, wire_1849, wire_1331, wire_11497, wire_9021, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8884, wire_1849, wire_1331, wire_11495, wire_9023, wire_8937, wire_8936, wire_8897, wire_8896, wire_8876, wire_8857, wire_8856, wire_1845, wire_1331, wire_11493, wire_9025, wire_8935, wire_8934, wire_8895, wire_8894, wire_8868, wire_8855, wire_8854, wire_1845, wire_1331, wire_11491, wire_9027, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8860, wire_1845, wire_1331, wire_11127, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11008, wire_8962, wire_1374, wire_11125, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_10980, wire_8954, wire_1374, wire_11123, wire_11039, wire_11038, wire_11029, wire_11028, wire_11019, wire_11018, wire_10982, wire_8946, wire_1374, wire_11121, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_10984, wire_8938, wire_1334, wire_11119, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_10986, wire_8930, wire_1334, wire_11117, wire_11037, wire_11036, wire_11027, wire_11026, wire_11017, wire_11016, wire_10988, wire_8922, wire_1334, wire_11115, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_10990, wire_8914, wire_1378, wire_1334, wire_11113, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_10992, wire_8906, wire_1378, wire_1334, wire_11111, wire_11035, wire_11034, wire_11025, wire_11024, wire_11015, wire_11014, wire_10994, wire_8898, wire_1378, wire_1334, wire_11109, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_10996, wire_8890, wire_1378, wire_1330, wire_11107, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_10998, wire_8882, wire_1378, wire_1330, wire_11105, wire_11033, wire_11032, wire_11023, wire_11022, wire_11013, wire_11012, wire_11000, wire_8874, wire_1378, wire_1330, wire_11103, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11002, wire_8866, wire_1374, wire_1330, wire_11101, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_11004, wire_8858, wire_1374, wire_1330, wire_11129, wire_11031, wire_11030, wire_11021, wire_11020, wire_11011, wire_11010, wire_11006, wire_8850, wire_1374, wire_1330, wire_11493, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11396, wire_9029, wire_1374, wire_11495, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11394, wire_9027, wire_1374, wire_11497, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11392, wire_9025, wire_1374, wire_11499, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11390, wire_9023, wire_1334, wire_11501, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11388, wire_9021, wire_1334, wire_11503, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11386, wire_9019, wire_1334, wire_11505, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11384, wire_9017, wire_1378, wire_1334, wire_11507, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11382, wire_9015, wire_1378, wire_1334, wire_11509, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11380, wire_9013, wire_1378, wire_1334, wire_11511, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11378, wire_9011, wire_1378, wire_1330, wire_11513, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11376, wire_9009, wire_1378, wire_1330, wire_11515, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11374, wire_9007, wire_1378, wire_1330, wire_11517, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11372, wire_9005, wire_1374, wire_1330, wire_11519, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11370, wire_9003, wire_1374, wire_1330, wire_11491, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11398, wire_9001, wire_1374, wire_1330};
    // CHNAXY TOTAL: 636
    assign wire_8853 = lut_tile_7_2_chanxy_out[0];
    assign wire_8861 = lut_tile_7_2_chanxy_out[1];
    assign wire_8869 = lut_tile_7_2_chanxy_out[2];
    assign wire_8877 = lut_tile_7_2_chanxy_out[3];
    assign wire_8885 = lut_tile_7_2_chanxy_out[4];
    assign wire_8893 = lut_tile_7_2_chanxy_out[5];
    assign wire_8901 = lut_tile_7_2_chanxy_out[6];
    assign wire_8909 = lut_tile_7_2_chanxy_out[7];
    assign wire_8917 = lut_tile_7_2_chanxy_out[8];
    assign wire_8925 = lut_tile_7_2_chanxy_out[9];
    assign wire_8933 = lut_tile_7_2_chanxy_out[10];
    assign wire_8941 = lut_tile_7_2_chanxy_out[11];
    assign wire_8949 = lut_tile_7_2_chanxy_out[12];
    assign wire_8957 = lut_tile_7_2_chanxy_out[13];
    assign wire_8965 = lut_tile_7_2_chanxy_out[14];
    assign wire_8970 = lut_tile_7_2_chanxy_out[15];
    assign wire_8972 = lut_tile_7_2_chanxy_out[16];
    assign wire_8974 = lut_tile_7_2_chanxy_out[17];
    assign wire_8976 = lut_tile_7_2_chanxy_out[18];
    assign wire_8978 = lut_tile_7_2_chanxy_out[19];
    assign wire_8980 = lut_tile_7_2_chanxy_out[20];
    assign wire_8982 = lut_tile_7_2_chanxy_out[21];
    assign wire_8984 = lut_tile_7_2_chanxy_out[22];
    assign wire_8986 = lut_tile_7_2_chanxy_out[23];
    assign wire_8988 = lut_tile_7_2_chanxy_out[24];
    assign wire_8990 = lut_tile_7_2_chanxy_out[25];
    assign wire_8992 = lut_tile_7_2_chanxy_out[26];
    assign wire_8994 = lut_tile_7_2_chanxy_out[27];
    assign wire_8996 = lut_tile_7_2_chanxy_out[28];
    assign wire_8998 = lut_tile_7_2_chanxy_out[29];
    assign wire_11371 = lut_tile_7_2_chanxy_out[30];
    assign wire_11373 = lut_tile_7_2_chanxy_out[31];
    assign wire_11375 = lut_tile_7_2_chanxy_out[32];
    assign wire_11377 = lut_tile_7_2_chanxy_out[33];
    assign wire_11379 = lut_tile_7_2_chanxy_out[34];
    assign wire_11381 = lut_tile_7_2_chanxy_out[35];
    assign wire_11383 = lut_tile_7_2_chanxy_out[36];
    assign wire_11385 = lut_tile_7_2_chanxy_out[37];
    assign wire_11387 = lut_tile_7_2_chanxy_out[38];
    assign wire_11389 = lut_tile_7_2_chanxy_out[39];
    assign wire_11391 = lut_tile_7_2_chanxy_out[40];
    assign wire_11393 = lut_tile_7_2_chanxy_out[41];
    assign wire_11395 = lut_tile_7_2_chanxy_out[42];
    assign wire_11397 = lut_tile_7_2_chanxy_out[43];
    assign wire_11399 = lut_tile_7_2_chanxy_out[44];
    assign wire_11460 = lut_tile_7_2_chanxy_out[45];
    assign wire_11462 = lut_tile_7_2_chanxy_out[46];
    assign wire_11464 = lut_tile_7_2_chanxy_out[47];
    assign wire_11466 = lut_tile_7_2_chanxy_out[48];
    assign wire_11468 = lut_tile_7_2_chanxy_out[49];
    assign wire_11470 = lut_tile_7_2_chanxy_out[50];
    assign wire_11472 = lut_tile_7_2_chanxy_out[51];
    assign wire_11474 = lut_tile_7_2_chanxy_out[52];
    assign wire_11476 = lut_tile_7_2_chanxy_out[53];
    assign wire_11478 = lut_tile_7_2_chanxy_out[54];
    assign wire_11480 = lut_tile_7_2_chanxy_out[55];
    assign wire_11482 = lut_tile_7_2_chanxy_out[56];
    assign wire_11484 = lut_tile_7_2_chanxy_out[57];
    assign wire_11486 = lut_tile_7_2_chanxy_out[58];
    assign wire_11488 = lut_tile_7_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_3_chanxy_in = {wire_11758, wire_8641, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8470, wire_2361, wire_11756, wire_8669, wire_8577, wire_8576, wire_8537, wire_8536, wire_8497, wire_8496, wire_8478, wire_2361, wire_11754, wire_8667, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8486, wire_2361, wire_11752, wire_8665, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8494, wire_1851, wire_11750, wire_8663, wire_8569, wire_8568, wire_8529, wire_8528, wire_8502, wire_8489, wire_8488, wire_1851, wire_11748, wire_8661, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8510, wire_1851, wire_11746, wire_8659, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8518, wire_2365, wire_1851, wire_11744, wire_8657, wire_8561, wire_8560, wire_8526, wire_8521, wire_8520, wire_8481, wire_8480, wire_2365, wire_1851, wire_11742, wire_8655, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8534, wire_2365, wire_1851, wire_11740, wire_8653, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8542, wire_2365, wire_1847, wire_11738, wire_8651, wire_8553, wire_8552, wire_8550, wire_8513, wire_8512, wire_8473, wire_8472, wire_2365, wire_1847, wire_11736, wire_8649, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8558, wire_2365, wire_1847, wire_11734, wire_8647, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8566, wire_2361, wire_1847, wire_11732, wire_8645, wire_8574, wire_8545, wire_8544, wire_8505, wire_8504, wire_8465, wire_8464, wire_2361, wire_1847, wire_11730, wire_8643, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8462, wire_2361, wire_1847, wire_11909, wire_9059, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8854, wire_2361, wire_11907, wire_9031, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8966, wire_2361, wire_11905, wire_9033, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8958, wire_2361, wire_11903, wire_9035, wire_8961, wire_8960, wire_8950, wire_8921, wire_8920, wire_8881, wire_8880, wire_1851, wire_11901, wire_9037, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8942, wire_1851, wire_11899, wire_9039, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8934, wire_1851, wire_11897, wire_9041, wire_8953, wire_8952, wire_8926, wire_8913, wire_8912, wire_8873, wire_8872, wire_2365, wire_1851, wire_11895, wire_9043, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8918, wire_2365, wire_1851, wire_11893, wire_9045, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8910, wire_2365, wire_1851, wire_11891, wire_9047, wire_8945, wire_8944, wire_8905, wire_8904, wire_8902, wire_8865, wire_8864, wire_2365, wire_1847, wire_11889, wire_9049, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8894, wire_2365, wire_1847, wire_11887, wire_9051, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8886, wire_2365, wire_1847, wire_11885, wire_9053, wire_8937, wire_8936, wire_8897, wire_8896, wire_8878, wire_8857, wire_8856, wire_2361, wire_1847, wire_11883, wire_9055, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8870, wire_2361, wire_1847, wire_11881, wire_9057, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8862, wire_2361, wire_1847, wire_11517, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11398, wire_8964, wire_1890, wire_11515, wire_11429, wire_11428, wire_11419, wire_11418, wire_11409, wire_11408, wire_11370, wire_8956, wire_1890, wire_11513, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11372, wire_8948, wire_1890, wire_11511, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11374, wire_8940, wire_1850, wire_11509, wire_11427, wire_11426, wire_11417, wire_11416, wire_11407, wire_11406, wire_11376, wire_8932, wire_1850, wire_11507, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11378, wire_8924, wire_1850, wire_11505, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11380, wire_8916, wire_1894, wire_1850, wire_11503, wire_11425, wire_11424, wire_11415, wire_11414, wire_11405, wire_11404, wire_11382, wire_8908, wire_1894, wire_1850, wire_11501, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11384, wire_8900, wire_1894, wire_1850, wire_11499, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11386, wire_8892, wire_1894, wire_1846, wire_11497, wire_11423, wire_11422, wire_11413, wire_11412, wire_11403, wire_11402, wire_11388, wire_8884, wire_1894, wire_1846, wire_11495, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11390, wire_8876, wire_1894, wire_1846, wire_11493, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11392, wire_8868, wire_1890, wire_1846, wire_11491, wire_11421, wire_11420, wire_11411, wire_11410, wire_11401, wire_11400, wire_11394, wire_8860, wire_1890, wire_1846, wire_11519, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11396, wire_8852, wire_1890, wire_1846, wire_11883, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11786, wire_9059, wire_1890, wire_11885, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11784, wire_9057, wire_1890, wire_11887, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11782, wire_9055, wire_1890, wire_11889, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11780, wire_9053, wire_1850, wire_11891, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11778, wire_9051, wire_1850, wire_11893, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11776, wire_9049, wire_1850, wire_11895, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11774, wire_9047, wire_1894, wire_1850, wire_11897, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11772, wire_9045, wire_1894, wire_1850, wire_11899, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11770, wire_9043, wire_1894, wire_1850, wire_11901, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11768, wire_9041, wire_1894, wire_1846, wire_11903, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11766, wire_9039, wire_1894, wire_1846, wire_11905, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11764, wire_9037, wire_1894, wire_1846, wire_11907, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11762, wire_9035, wire_1890, wire_1846, wire_11909, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11760, wire_9033, wire_1890, wire_1846, wire_11881, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11788, wire_9031, wire_1890, wire_1846};
    // CHNAXY TOTAL: 636
    assign wire_8855 = lut_tile_7_3_chanxy_out[0];
    assign wire_8863 = lut_tile_7_3_chanxy_out[1];
    assign wire_8871 = lut_tile_7_3_chanxy_out[2];
    assign wire_8879 = lut_tile_7_3_chanxy_out[3];
    assign wire_8887 = lut_tile_7_3_chanxy_out[4];
    assign wire_8895 = lut_tile_7_3_chanxy_out[5];
    assign wire_8903 = lut_tile_7_3_chanxy_out[6];
    assign wire_8911 = lut_tile_7_3_chanxy_out[7];
    assign wire_8919 = lut_tile_7_3_chanxy_out[8];
    assign wire_8927 = lut_tile_7_3_chanxy_out[9];
    assign wire_8935 = lut_tile_7_3_chanxy_out[10];
    assign wire_8943 = lut_tile_7_3_chanxy_out[11];
    assign wire_8951 = lut_tile_7_3_chanxy_out[12];
    assign wire_8959 = lut_tile_7_3_chanxy_out[13];
    assign wire_8967 = lut_tile_7_3_chanxy_out[14];
    assign wire_9000 = lut_tile_7_3_chanxy_out[15];
    assign wire_9002 = lut_tile_7_3_chanxy_out[16];
    assign wire_9004 = lut_tile_7_3_chanxy_out[17];
    assign wire_9006 = lut_tile_7_3_chanxy_out[18];
    assign wire_9008 = lut_tile_7_3_chanxy_out[19];
    assign wire_9010 = lut_tile_7_3_chanxy_out[20];
    assign wire_9012 = lut_tile_7_3_chanxy_out[21];
    assign wire_9014 = lut_tile_7_3_chanxy_out[22];
    assign wire_9016 = lut_tile_7_3_chanxy_out[23];
    assign wire_9018 = lut_tile_7_3_chanxy_out[24];
    assign wire_9020 = lut_tile_7_3_chanxy_out[25];
    assign wire_9022 = lut_tile_7_3_chanxy_out[26];
    assign wire_9024 = lut_tile_7_3_chanxy_out[27];
    assign wire_9026 = lut_tile_7_3_chanxy_out[28];
    assign wire_9028 = lut_tile_7_3_chanxy_out[29];
    assign wire_11761 = lut_tile_7_3_chanxy_out[30];
    assign wire_11763 = lut_tile_7_3_chanxy_out[31];
    assign wire_11765 = lut_tile_7_3_chanxy_out[32];
    assign wire_11767 = lut_tile_7_3_chanxy_out[33];
    assign wire_11769 = lut_tile_7_3_chanxy_out[34];
    assign wire_11771 = lut_tile_7_3_chanxy_out[35];
    assign wire_11773 = lut_tile_7_3_chanxy_out[36];
    assign wire_11775 = lut_tile_7_3_chanxy_out[37];
    assign wire_11777 = lut_tile_7_3_chanxy_out[38];
    assign wire_11779 = lut_tile_7_3_chanxy_out[39];
    assign wire_11781 = lut_tile_7_3_chanxy_out[40];
    assign wire_11783 = lut_tile_7_3_chanxy_out[41];
    assign wire_11785 = lut_tile_7_3_chanxy_out[42];
    assign wire_11787 = lut_tile_7_3_chanxy_out[43];
    assign wire_11789 = lut_tile_7_3_chanxy_out[44];
    assign wire_11850 = lut_tile_7_3_chanxy_out[45];
    assign wire_11852 = lut_tile_7_3_chanxy_out[46];
    assign wire_11854 = lut_tile_7_3_chanxy_out[47];
    assign wire_11856 = lut_tile_7_3_chanxy_out[48];
    assign wire_11858 = lut_tile_7_3_chanxy_out[49];
    assign wire_11860 = lut_tile_7_3_chanxy_out[50];
    assign wire_11862 = lut_tile_7_3_chanxy_out[51];
    assign wire_11864 = lut_tile_7_3_chanxy_out[52];
    assign wire_11866 = lut_tile_7_3_chanxy_out[53];
    assign wire_11868 = lut_tile_7_3_chanxy_out[54];
    assign wire_11870 = lut_tile_7_3_chanxy_out[55];
    assign wire_11872 = lut_tile_7_3_chanxy_out[56];
    assign wire_11874 = lut_tile_7_3_chanxy_out[57];
    assign wire_11876 = lut_tile_7_3_chanxy_out[58];
    assign wire_11878 = lut_tile_7_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_4_chanxy_in = {wire_12148, wire_8671, wire_8609, wire_8608, wire_8599, wire_8598, wire_8589, wire_8588, wire_8472, wire_2877, wire_12146, wire_8699, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8480, wire_2877, wire_12144, wire_8697, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8488, wire_2877, wire_12142, wire_8695, wire_8607, wire_8606, wire_8597, wire_8596, wire_8587, wire_8586, wire_8496, wire_2367, wire_12140, wire_8693, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8504, wire_2367, wire_12138, wire_8691, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8512, wire_2367, wire_12136, wire_8689, wire_8605, wire_8604, wire_8595, wire_8594, wire_8585, wire_8584, wire_8520, wire_2881, wire_2367, wire_12134, wire_8687, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8528, wire_2881, wire_2367, wire_12132, wire_8685, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8536, wire_2881, wire_2367, wire_12130, wire_8683, wire_8603, wire_8602, wire_8593, wire_8592, wire_8583, wire_8582, wire_8544, wire_2881, wire_2363, wire_12128, wire_8681, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8552, wire_2881, wire_2363, wire_12126, wire_8679, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8560, wire_2881, wire_2363, wire_12124, wire_8677, wire_8601, wire_8600, wire_8591, wire_8590, wire_8581, wire_8580, wire_8568, wire_2877, wire_2363, wire_12122, wire_8675, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8576, wire_2877, wire_2363, wire_12120, wire_8673, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8464, wire_2877, wire_2363, wire_12299, wire_9089, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8856, wire_2877, wire_12297, wire_9061, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8968, wire_2877, wire_12295, wire_9063, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8960, wire_2877, wire_12293, wire_9065, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8952, wire_2367, wire_12291, wire_9067, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8944, wire_2367, wire_12289, wire_9069, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8936, wire_2367, wire_12287, wire_9071, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8928, wire_2881, wire_2367, wire_12285, wire_9073, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8920, wire_2881, wire_2367, wire_12283, wire_9075, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8912, wire_2881, wire_2367, wire_12281, wire_9077, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8904, wire_2881, wire_2363, wire_12279, wire_9079, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8896, wire_2881, wire_2363, wire_12277, wire_9081, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8888, wire_2881, wire_2363, wire_12275, wire_9083, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8880, wire_2877, wire_2363, wire_12273, wire_9085, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8872, wire_2877, wire_2363, wire_12271, wire_9087, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8864, wire_2877, wire_2363, wire_11907, wire_11819, wire_11818, wire_11809, wire_11808, wire_11799, wire_11798, wire_11788, wire_8966, wire_2406, wire_11905, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11760, wire_8958, wire_2406, wire_11903, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11762, wire_8950, wire_2406, wire_11901, wire_11817, wire_11816, wire_11807, wire_11806, wire_11797, wire_11796, wire_11764, wire_8942, wire_2366, wire_11899, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11766, wire_8934, wire_2366, wire_11897, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11768, wire_8926, wire_2366, wire_11895, wire_11815, wire_11814, wire_11805, wire_11804, wire_11795, wire_11794, wire_11770, wire_8918, wire_2410, wire_2366, wire_11893, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11772, wire_8910, wire_2410, wire_2366, wire_11891, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11774, wire_8902, wire_2410, wire_2366, wire_11889, wire_11813, wire_11812, wire_11803, wire_11802, wire_11793, wire_11792, wire_11776, wire_8894, wire_2410, wire_2362, wire_11887, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11778, wire_8886, wire_2410, wire_2362, wire_11885, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11780, wire_8878, wire_2410, wire_2362, wire_11883, wire_11811, wire_11810, wire_11801, wire_11800, wire_11791, wire_11790, wire_11782, wire_8870, wire_2406, wire_2362, wire_11881, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11784, wire_8862, wire_2406, wire_2362, wire_11909, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11786, wire_8854, wire_2406, wire_2362, wire_12273, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12176, wire_9089, wire_2406, wire_12275, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12174, wire_9087, wire_2406, wire_12277, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12172, wire_9085, wire_2406, wire_12279, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12170, wire_9083, wire_2366, wire_12281, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12168, wire_9081, wire_2366, wire_12283, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12166, wire_9079, wire_2366, wire_12285, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12164, wire_9077, wire_2410, wire_2366, wire_12287, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12162, wire_9075, wire_2410, wire_2366, wire_12289, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12160, wire_9073, wire_2410, wire_2366, wire_12291, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12158, wire_9071, wire_2410, wire_2362, wire_12293, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12156, wire_9069, wire_2410, wire_2362, wire_12295, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12154, wire_9067, wire_2410, wire_2362, wire_12297, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12152, wire_9065, wire_2406, wire_2362, wire_12299, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12150, wire_9063, wire_2406, wire_2362, wire_12271, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12178, wire_9061, wire_2406, wire_2362};
    // CHNAXY TOTAL: 636
    assign wire_8857 = lut_tile_7_4_chanxy_out[0];
    assign wire_8865 = lut_tile_7_4_chanxy_out[1];
    assign wire_8873 = lut_tile_7_4_chanxy_out[2];
    assign wire_8881 = lut_tile_7_4_chanxy_out[3];
    assign wire_8889 = lut_tile_7_4_chanxy_out[4];
    assign wire_8897 = lut_tile_7_4_chanxy_out[5];
    assign wire_8905 = lut_tile_7_4_chanxy_out[6];
    assign wire_8913 = lut_tile_7_4_chanxy_out[7];
    assign wire_8921 = lut_tile_7_4_chanxy_out[8];
    assign wire_8929 = lut_tile_7_4_chanxy_out[9];
    assign wire_8937 = lut_tile_7_4_chanxy_out[10];
    assign wire_8945 = lut_tile_7_4_chanxy_out[11];
    assign wire_8953 = lut_tile_7_4_chanxy_out[12];
    assign wire_8961 = lut_tile_7_4_chanxy_out[13];
    assign wire_8969 = lut_tile_7_4_chanxy_out[14];
    assign wire_9030 = lut_tile_7_4_chanxy_out[15];
    assign wire_9032 = lut_tile_7_4_chanxy_out[16];
    assign wire_9034 = lut_tile_7_4_chanxy_out[17];
    assign wire_9036 = lut_tile_7_4_chanxy_out[18];
    assign wire_9038 = lut_tile_7_4_chanxy_out[19];
    assign wire_9040 = lut_tile_7_4_chanxy_out[20];
    assign wire_9042 = lut_tile_7_4_chanxy_out[21];
    assign wire_9044 = lut_tile_7_4_chanxy_out[22];
    assign wire_9046 = lut_tile_7_4_chanxy_out[23];
    assign wire_9048 = lut_tile_7_4_chanxy_out[24];
    assign wire_9050 = lut_tile_7_4_chanxy_out[25];
    assign wire_9052 = lut_tile_7_4_chanxy_out[26];
    assign wire_9054 = lut_tile_7_4_chanxy_out[27];
    assign wire_9056 = lut_tile_7_4_chanxy_out[28];
    assign wire_9058 = lut_tile_7_4_chanxy_out[29];
    assign wire_12151 = lut_tile_7_4_chanxy_out[30];
    assign wire_12153 = lut_tile_7_4_chanxy_out[31];
    assign wire_12155 = lut_tile_7_4_chanxy_out[32];
    assign wire_12157 = lut_tile_7_4_chanxy_out[33];
    assign wire_12159 = lut_tile_7_4_chanxy_out[34];
    assign wire_12161 = lut_tile_7_4_chanxy_out[35];
    assign wire_12163 = lut_tile_7_4_chanxy_out[36];
    assign wire_12165 = lut_tile_7_4_chanxy_out[37];
    assign wire_12167 = lut_tile_7_4_chanxy_out[38];
    assign wire_12169 = lut_tile_7_4_chanxy_out[39];
    assign wire_12171 = lut_tile_7_4_chanxy_out[40];
    assign wire_12173 = lut_tile_7_4_chanxy_out[41];
    assign wire_12175 = lut_tile_7_4_chanxy_out[42];
    assign wire_12177 = lut_tile_7_4_chanxy_out[43];
    assign wire_12179 = lut_tile_7_4_chanxy_out[44];
    assign wire_12240 = lut_tile_7_4_chanxy_out[45];
    assign wire_12242 = lut_tile_7_4_chanxy_out[46];
    assign wire_12244 = lut_tile_7_4_chanxy_out[47];
    assign wire_12246 = lut_tile_7_4_chanxy_out[48];
    assign wire_12248 = lut_tile_7_4_chanxy_out[49];
    assign wire_12250 = lut_tile_7_4_chanxy_out[50];
    assign wire_12252 = lut_tile_7_4_chanxy_out[51];
    assign wire_12254 = lut_tile_7_4_chanxy_out[52];
    assign wire_12256 = lut_tile_7_4_chanxy_out[53];
    assign wire_12258 = lut_tile_7_4_chanxy_out[54];
    assign wire_12260 = lut_tile_7_4_chanxy_out[55];
    assign wire_12262 = lut_tile_7_4_chanxy_out[56];
    assign wire_12264 = lut_tile_7_4_chanxy_out[57];
    assign wire_12266 = lut_tile_7_4_chanxy_out[58];
    assign wire_12268 = lut_tile_7_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_5_chanxy_in = {wire_12538, wire_8701, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8582, wire_3393, wire_12536, wire_8729, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8584, wire_3393, wire_12534, wire_8727, wire_8639, wire_8638, wire_8629, wire_8628, wire_8619, wire_8618, wire_8586, wire_3393, wire_12532, wire_8725, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8588, wire_2883, wire_12530, wire_8723, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8590, wire_2883, wire_12528, wire_8721, wire_8637, wire_8636, wire_8627, wire_8626, wire_8617, wire_8616, wire_8592, wire_2883, wire_12526, wire_8719, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8594, wire_3397, wire_2883, wire_12524, wire_8717, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8596, wire_3397, wire_2883, wire_12522, wire_8715, wire_8635, wire_8634, wire_8625, wire_8624, wire_8615, wire_8614, wire_8598, wire_3397, wire_2883, wire_12520, wire_8713, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8600, wire_3397, wire_2879, wire_12518, wire_8711, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8602, wire_3397, wire_2879, wire_12516, wire_8709, wire_8633, wire_8632, wire_8623, wire_8622, wire_8613, wire_8612, wire_8604, wire_3397, wire_2879, wire_12514, wire_8707, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8606, wire_3393, wire_2879, wire_12512, wire_8705, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8608, wire_3393, wire_2879, wire_12510, wire_8703, wire_8631, wire_8630, wire_8621, wire_8620, wire_8611, wire_8610, wire_8580, wire_3393, wire_2879, wire_12689, wire_9119, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_8970, wire_3393, wire_12687, wire_9091, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8998, wire_3393, wire_12685, wire_9093, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8996, wire_3393, wire_12683, wire_9095, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_8994, wire_2883, wire_12681, wire_9097, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8992, wire_2883, wire_12679, wire_9099, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8990, wire_2883, wire_12677, wire_9101, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_8988, wire_3397, wire_2883, wire_12675, wire_9103, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8986, wire_3397, wire_2883, wire_12673, wire_9105, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8984, wire_3397, wire_2883, wire_12671, wire_9107, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_8982, wire_3397, wire_2879, wire_12669, wire_9109, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8980, wire_3397, wire_2879, wire_12667, wire_9111, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8978, wire_3397, wire_2879, wire_12665, wire_9113, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_8976, wire_3393, wire_2879, wire_12663, wire_9115, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8974, wire_3393, wire_2879, wire_12661, wire_9117, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8972, wire_3393, wire_2879, wire_12297, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12178, wire_8968, wire_2922, wire_12295, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12150, wire_8960, wire_2922, wire_12293, wire_12209, wire_12208, wire_12199, wire_12198, wire_12189, wire_12188, wire_12152, wire_8952, wire_2922, wire_12291, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12154, wire_8944, wire_2882, wire_12289, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12156, wire_8936, wire_2882, wire_12287, wire_12207, wire_12206, wire_12197, wire_12196, wire_12187, wire_12186, wire_12158, wire_8928, wire_2882, wire_12285, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12160, wire_8920, wire_2926, wire_2882, wire_12283, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12162, wire_8912, wire_2926, wire_2882, wire_12281, wire_12205, wire_12204, wire_12195, wire_12194, wire_12185, wire_12184, wire_12164, wire_8904, wire_2926, wire_2882, wire_12279, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12166, wire_8896, wire_2926, wire_2878, wire_12277, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12168, wire_8888, wire_2926, wire_2878, wire_12275, wire_12203, wire_12202, wire_12193, wire_12192, wire_12183, wire_12182, wire_12170, wire_8880, wire_2926, wire_2878, wire_12273, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12172, wire_8872, wire_2922, wire_2878, wire_12271, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12174, wire_8864, wire_2922, wire_2878, wire_12299, wire_12201, wire_12200, wire_12191, wire_12190, wire_12181, wire_12180, wire_12176, wire_8856, wire_2922, wire_2878, wire_12663, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12566, wire_9119, wire_2922, wire_12665, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12564, wire_9117, wire_2922, wire_12667, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12562, wire_9115, wire_2922, wire_12669, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12560, wire_9113, wire_2882, wire_12671, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12558, wire_9111, wire_2882, wire_12673, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12556, wire_9109, wire_2882, wire_12675, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12554, wire_9107, wire_2926, wire_2882, wire_12677, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12552, wire_9105, wire_2926, wire_2882, wire_12679, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12550, wire_9103, wire_2926, wire_2882, wire_12681, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12548, wire_9101, wire_2926, wire_2878, wire_12683, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12546, wire_9099, wire_2926, wire_2878, wire_12685, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12544, wire_9097, wire_2926, wire_2878, wire_12687, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12542, wire_9095, wire_2922, wire_2878, wire_12689, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12540, wire_9093, wire_2922, wire_2878, wire_12661, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12568, wire_9091, wire_2922, wire_2878};
    // CHNAXY TOTAL: 636
    assign wire_8971 = lut_tile_7_5_chanxy_out[0];
    assign wire_8973 = lut_tile_7_5_chanxy_out[1];
    assign wire_8975 = lut_tile_7_5_chanxy_out[2];
    assign wire_8977 = lut_tile_7_5_chanxy_out[3];
    assign wire_8979 = lut_tile_7_5_chanxy_out[4];
    assign wire_8981 = lut_tile_7_5_chanxy_out[5];
    assign wire_8983 = lut_tile_7_5_chanxy_out[6];
    assign wire_8985 = lut_tile_7_5_chanxy_out[7];
    assign wire_8987 = lut_tile_7_5_chanxy_out[8];
    assign wire_8989 = lut_tile_7_5_chanxy_out[9];
    assign wire_8991 = lut_tile_7_5_chanxy_out[10];
    assign wire_8993 = lut_tile_7_5_chanxy_out[11];
    assign wire_8995 = lut_tile_7_5_chanxy_out[12];
    assign wire_8997 = lut_tile_7_5_chanxy_out[13];
    assign wire_8999 = lut_tile_7_5_chanxy_out[14];
    assign wire_9060 = lut_tile_7_5_chanxy_out[15];
    assign wire_9062 = lut_tile_7_5_chanxy_out[16];
    assign wire_9064 = lut_tile_7_5_chanxy_out[17];
    assign wire_9066 = lut_tile_7_5_chanxy_out[18];
    assign wire_9068 = lut_tile_7_5_chanxy_out[19];
    assign wire_9070 = lut_tile_7_5_chanxy_out[20];
    assign wire_9072 = lut_tile_7_5_chanxy_out[21];
    assign wire_9074 = lut_tile_7_5_chanxy_out[22];
    assign wire_9076 = lut_tile_7_5_chanxy_out[23];
    assign wire_9078 = lut_tile_7_5_chanxy_out[24];
    assign wire_9080 = lut_tile_7_5_chanxy_out[25];
    assign wire_9082 = lut_tile_7_5_chanxy_out[26];
    assign wire_9084 = lut_tile_7_5_chanxy_out[27];
    assign wire_9086 = lut_tile_7_5_chanxy_out[28];
    assign wire_9088 = lut_tile_7_5_chanxy_out[29];
    assign wire_12541 = lut_tile_7_5_chanxy_out[30];
    assign wire_12543 = lut_tile_7_5_chanxy_out[31];
    assign wire_12545 = lut_tile_7_5_chanxy_out[32];
    assign wire_12547 = lut_tile_7_5_chanxy_out[33];
    assign wire_12549 = lut_tile_7_5_chanxy_out[34];
    assign wire_12551 = lut_tile_7_5_chanxy_out[35];
    assign wire_12553 = lut_tile_7_5_chanxy_out[36];
    assign wire_12555 = lut_tile_7_5_chanxy_out[37];
    assign wire_12557 = lut_tile_7_5_chanxy_out[38];
    assign wire_12559 = lut_tile_7_5_chanxy_out[39];
    assign wire_12561 = lut_tile_7_5_chanxy_out[40];
    assign wire_12563 = lut_tile_7_5_chanxy_out[41];
    assign wire_12565 = lut_tile_7_5_chanxy_out[42];
    assign wire_12567 = lut_tile_7_5_chanxy_out[43];
    assign wire_12569 = lut_tile_7_5_chanxy_out[44];
    assign wire_12630 = lut_tile_7_5_chanxy_out[45];
    assign wire_12632 = lut_tile_7_5_chanxy_out[46];
    assign wire_12634 = lut_tile_7_5_chanxy_out[47];
    assign wire_12636 = lut_tile_7_5_chanxy_out[48];
    assign wire_12638 = lut_tile_7_5_chanxy_out[49];
    assign wire_12640 = lut_tile_7_5_chanxy_out[50];
    assign wire_12642 = lut_tile_7_5_chanxy_out[51];
    assign wire_12644 = lut_tile_7_5_chanxy_out[52];
    assign wire_12646 = lut_tile_7_5_chanxy_out[53];
    assign wire_12648 = lut_tile_7_5_chanxy_out[54];
    assign wire_12650 = lut_tile_7_5_chanxy_out[55];
    assign wire_12652 = lut_tile_7_5_chanxy_out[56];
    assign wire_12654 = lut_tile_7_5_chanxy_out[57];
    assign wire_12656 = lut_tile_7_5_chanxy_out[58];
    assign wire_12658 = lut_tile_7_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_6_chanxy_in = {wire_12928, wire_8731, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8612, wire_3909, wire_12926, wire_8759, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8614, wire_3909, wire_12924, wire_8757, wire_8669, wire_8668, wire_8659, wire_8658, wire_8649, wire_8648, wire_8616, wire_3909, wire_12922, wire_8755, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8618, wire_3399, wire_12920, wire_8753, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8620, wire_3399, wire_12918, wire_8751, wire_8667, wire_8666, wire_8657, wire_8656, wire_8647, wire_8646, wire_8622, wire_3399, wire_12916, wire_8749, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8624, wire_3913, wire_3399, wire_12914, wire_8747, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8626, wire_3913, wire_3399, wire_12912, wire_8745, wire_8665, wire_8664, wire_8655, wire_8654, wire_8645, wire_8644, wire_8628, wire_3913, wire_3399, wire_12910, wire_8743, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8630, wire_3913, wire_3395, wire_12908, wire_8741, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8632, wire_3913, wire_3395, wire_12906, wire_8739, wire_8663, wire_8662, wire_8653, wire_8652, wire_8643, wire_8642, wire_8634, wire_3913, wire_3395, wire_12904, wire_8737, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8636, wire_3909, wire_3395, wire_12902, wire_8735, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8638, wire_3909, wire_3395, wire_12900, wire_8733, wire_8661, wire_8660, wire_8651, wire_8650, wire_8641, wire_8640, wire_8610, wire_3909, wire_3395, wire_13079, wire_9149, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9000, wire_3909, wire_13077, wire_9121, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_9028, wire_3909, wire_13075, wire_9123, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9026, wire_3909, wire_13073, wire_9125, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9024, wire_3399, wire_13071, wire_9127, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_9022, wire_3399, wire_13069, wire_9129, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9020, wire_3399, wire_13067, wire_9131, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9018, wire_3913, wire_3399, wire_13065, wire_9133, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_9016, wire_3913, wire_3399, wire_13063, wire_9135, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9014, wire_3913, wire_3399, wire_13061, wire_9137, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9012, wire_3913, wire_3395, wire_13059, wire_9139, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_9010, wire_3913, wire_3395, wire_13057, wire_9141, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9008, wire_3913, wire_3395, wire_13055, wire_9143, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9006, wire_3909, wire_3395, wire_13053, wire_9145, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_9004, wire_3909, wire_3395, wire_13051, wire_9147, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9002, wire_3909, wire_3395, wire_12687, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12568, wire_8998, wire_3438, wire_12685, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12540, wire_8996, wire_3438, wire_12683, wire_12599, wire_12598, wire_12589, wire_12588, wire_12579, wire_12578, wire_12542, wire_8994, wire_3438, wire_12681, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12544, wire_8992, wire_3398, wire_12679, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12546, wire_8990, wire_3398, wire_12677, wire_12597, wire_12596, wire_12587, wire_12586, wire_12577, wire_12576, wire_12548, wire_8988, wire_3398, wire_12675, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12550, wire_8986, wire_3442, wire_3398, wire_12673, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12552, wire_8984, wire_3442, wire_3398, wire_12671, wire_12595, wire_12594, wire_12585, wire_12584, wire_12575, wire_12574, wire_12554, wire_8982, wire_3442, wire_3398, wire_12669, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12556, wire_8980, wire_3442, wire_3394, wire_12667, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12558, wire_8978, wire_3442, wire_3394, wire_12665, wire_12593, wire_12592, wire_12583, wire_12582, wire_12573, wire_12572, wire_12560, wire_8976, wire_3442, wire_3394, wire_12663, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12562, wire_8974, wire_3438, wire_3394, wire_12661, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12564, wire_8972, wire_3438, wire_3394, wire_12689, wire_12591, wire_12590, wire_12581, wire_12580, wire_12571, wire_12570, wire_12566, wire_8970, wire_3438, wire_3394, wire_13053, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12956, wire_9149, wire_3438, wire_13055, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12954, wire_9147, wire_3438, wire_13057, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12952, wire_9145, wire_3438, wire_13059, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12950, wire_9143, wire_3398, wire_13061, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12948, wire_9141, wire_3398, wire_13063, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12946, wire_9139, wire_3398, wire_13065, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12944, wire_9137, wire_3442, wire_3398, wire_13067, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12942, wire_9135, wire_3442, wire_3398, wire_13069, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12940, wire_9133, wire_3442, wire_3398, wire_13071, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12938, wire_9131, wire_3442, wire_3394, wire_13073, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12936, wire_9129, wire_3442, wire_3394, wire_13075, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12934, wire_9127, wire_3442, wire_3394, wire_13077, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12932, wire_9125, wire_3438, wire_3394, wire_13079, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12930, wire_9123, wire_3438, wire_3394, wire_13051, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12958, wire_9121, wire_3438, wire_3394};
    // CHNAXY TOTAL: 636
    assign wire_9001 = lut_tile_7_6_chanxy_out[0];
    assign wire_9003 = lut_tile_7_6_chanxy_out[1];
    assign wire_9005 = lut_tile_7_6_chanxy_out[2];
    assign wire_9007 = lut_tile_7_6_chanxy_out[3];
    assign wire_9009 = lut_tile_7_6_chanxy_out[4];
    assign wire_9011 = lut_tile_7_6_chanxy_out[5];
    assign wire_9013 = lut_tile_7_6_chanxy_out[6];
    assign wire_9015 = lut_tile_7_6_chanxy_out[7];
    assign wire_9017 = lut_tile_7_6_chanxy_out[8];
    assign wire_9019 = lut_tile_7_6_chanxy_out[9];
    assign wire_9021 = lut_tile_7_6_chanxy_out[10];
    assign wire_9023 = lut_tile_7_6_chanxy_out[11];
    assign wire_9025 = lut_tile_7_6_chanxy_out[12];
    assign wire_9027 = lut_tile_7_6_chanxy_out[13];
    assign wire_9029 = lut_tile_7_6_chanxy_out[14];
    assign wire_9090 = lut_tile_7_6_chanxy_out[15];
    assign wire_9092 = lut_tile_7_6_chanxy_out[16];
    assign wire_9094 = lut_tile_7_6_chanxy_out[17];
    assign wire_9096 = lut_tile_7_6_chanxy_out[18];
    assign wire_9098 = lut_tile_7_6_chanxy_out[19];
    assign wire_9100 = lut_tile_7_6_chanxy_out[20];
    assign wire_9102 = lut_tile_7_6_chanxy_out[21];
    assign wire_9104 = lut_tile_7_6_chanxy_out[22];
    assign wire_9106 = lut_tile_7_6_chanxy_out[23];
    assign wire_9108 = lut_tile_7_6_chanxy_out[24];
    assign wire_9110 = lut_tile_7_6_chanxy_out[25];
    assign wire_9112 = lut_tile_7_6_chanxy_out[26];
    assign wire_9114 = lut_tile_7_6_chanxy_out[27];
    assign wire_9116 = lut_tile_7_6_chanxy_out[28];
    assign wire_9118 = lut_tile_7_6_chanxy_out[29];
    assign wire_12931 = lut_tile_7_6_chanxy_out[30];
    assign wire_12933 = lut_tile_7_6_chanxy_out[31];
    assign wire_12935 = lut_tile_7_6_chanxy_out[32];
    assign wire_12937 = lut_tile_7_6_chanxy_out[33];
    assign wire_12939 = lut_tile_7_6_chanxy_out[34];
    assign wire_12941 = lut_tile_7_6_chanxy_out[35];
    assign wire_12943 = lut_tile_7_6_chanxy_out[36];
    assign wire_12945 = lut_tile_7_6_chanxy_out[37];
    assign wire_12947 = lut_tile_7_6_chanxy_out[38];
    assign wire_12949 = lut_tile_7_6_chanxy_out[39];
    assign wire_12951 = lut_tile_7_6_chanxy_out[40];
    assign wire_12953 = lut_tile_7_6_chanxy_out[41];
    assign wire_12955 = lut_tile_7_6_chanxy_out[42];
    assign wire_12957 = lut_tile_7_6_chanxy_out[43];
    assign wire_12959 = lut_tile_7_6_chanxy_out[44];
    assign wire_13020 = lut_tile_7_6_chanxy_out[45];
    assign wire_13022 = lut_tile_7_6_chanxy_out[46];
    assign wire_13024 = lut_tile_7_6_chanxy_out[47];
    assign wire_13026 = lut_tile_7_6_chanxy_out[48];
    assign wire_13028 = lut_tile_7_6_chanxy_out[49];
    assign wire_13030 = lut_tile_7_6_chanxy_out[50];
    assign wire_13032 = lut_tile_7_6_chanxy_out[51];
    assign wire_13034 = lut_tile_7_6_chanxy_out[52];
    assign wire_13036 = lut_tile_7_6_chanxy_out[53];
    assign wire_13038 = lut_tile_7_6_chanxy_out[54];
    assign wire_13040 = lut_tile_7_6_chanxy_out[55];
    assign wire_13042 = lut_tile_7_6_chanxy_out[56];
    assign wire_13044 = lut_tile_7_6_chanxy_out[57];
    assign wire_13046 = lut_tile_7_6_chanxy_out[58];
    assign wire_13048 = lut_tile_7_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_7_chanxy_in = {wire_13318, wire_8761, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8642, wire_4425, wire_13316, wire_8789, wire_8699, wire_8698, wire_8689, wire_8688, wire_8679, wire_8678, wire_8644, wire_4425, wire_13314, wire_8787, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8646, wire_4425, wire_13312, wire_8785, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8648, wire_3915, wire_13310, wire_8783, wire_8697, wire_8696, wire_8687, wire_8686, wire_8677, wire_8676, wire_8650, wire_3915, wire_13308, wire_8781, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8652, wire_3915, wire_13306, wire_8779, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8654, wire_4429, wire_3915, wire_13304, wire_8777, wire_8695, wire_8694, wire_8685, wire_8684, wire_8675, wire_8674, wire_8656, wire_4429, wire_3915, wire_13302, wire_8775, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8658, wire_4429, wire_3915, wire_13300, wire_8773, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8660, wire_4429, wire_3911, wire_13298, wire_8771, wire_8693, wire_8692, wire_8683, wire_8682, wire_8673, wire_8672, wire_8662, wire_4429, wire_3911, wire_13296, wire_8769, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8664, wire_4429, wire_3911, wire_13294, wire_8767, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8666, wire_4425, wire_3911, wire_13292, wire_8765, wire_8691, wire_8690, wire_8681, wire_8680, wire_8671, wire_8670, wire_8668, wire_4425, wire_3911, wire_13290, wire_8763, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8640, wire_4425, wire_3911, wire_13469, wire_9179, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9030, wire_4425, wire_13467, wire_9151, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9058, wire_4425, wire_13465, wire_9153, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9056, wire_4425, wire_13463, wire_9155, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9054, wire_3915, wire_13461, wire_9157, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9052, wire_3915, wire_13459, wire_9159, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9050, wire_3915, wire_13457, wire_9161, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9048, wire_4429, wire_3915, wire_13455, wire_9163, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9046, wire_4429, wire_3915, wire_13453, wire_9165, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9044, wire_4429, wire_3915, wire_13451, wire_9167, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9042, wire_4429, wire_3911, wire_13449, wire_9169, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9040, wire_4429, wire_3911, wire_13447, wire_9171, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9038, wire_4429, wire_3911, wire_13445, wire_9173, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9036, wire_4425, wire_3911, wire_13443, wire_9175, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9034, wire_4425, wire_3911, wire_13441, wire_9177, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9032, wire_4425, wire_3911, wire_13077, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12958, wire_9028, wire_3954, wire_13075, wire_12989, wire_12988, wire_12979, wire_12978, wire_12969, wire_12968, wire_12930, wire_9026, wire_3954, wire_13073, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12932, wire_9024, wire_3954, wire_13071, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12934, wire_9022, wire_3914, wire_13069, wire_12987, wire_12986, wire_12977, wire_12976, wire_12967, wire_12966, wire_12936, wire_9020, wire_3914, wire_13067, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12938, wire_9018, wire_3914, wire_13065, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12940, wire_9016, wire_3958, wire_3914, wire_13063, wire_12985, wire_12984, wire_12975, wire_12974, wire_12965, wire_12964, wire_12942, wire_9014, wire_3958, wire_3914, wire_13061, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12944, wire_9012, wire_3958, wire_3914, wire_13059, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12946, wire_9010, wire_3958, wire_3910, wire_13057, wire_12983, wire_12982, wire_12973, wire_12972, wire_12963, wire_12962, wire_12948, wire_9008, wire_3958, wire_3910, wire_13055, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12950, wire_9006, wire_3958, wire_3910, wire_13053, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12952, wire_9004, wire_3954, wire_3910, wire_13051, wire_12981, wire_12980, wire_12971, wire_12970, wire_12961, wire_12960, wire_12954, wire_9002, wire_3954, wire_3910, wire_13079, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12956, wire_9000, wire_3954, wire_3910, wire_13443, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13346, wire_9179, wire_3954, wire_13445, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13344, wire_9177, wire_3954, wire_13447, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13342, wire_9175, wire_3954, wire_13449, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13340, wire_9173, wire_3914, wire_13451, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13338, wire_9171, wire_3914, wire_13453, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13336, wire_9169, wire_3914, wire_13455, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13334, wire_9167, wire_3958, wire_3914, wire_13457, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13332, wire_9165, wire_3958, wire_3914, wire_13459, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13330, wire_9163, wire_3958, wire_3914, wire_13461, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13328, wire_9161, wire_3958, wire_3910, wire_13463, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13326, wire_9159, wire_3958, wire_3910, wire_13465, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13324, wire_9157, wire_3958, wire_3910, wire_13467, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13322, wire_9155, wire_3954, wire_3910, wire_13469, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13320, wire_9153, wire_3954, wire_3910, wire_13441, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13348, wire_9151, wire_3954, wire_3910};
    // CHNAXY TOTAL: 636
    assign wire_9031 = lut_tile_7_7_chanxy_out[0];
    assign wire_9033 = lut_tile_7_7_chanxy_out[1];
    assign wire_9035 = lut_tile_7_7_chanxy_out[2];
    assign wire_9037 = lut_tile_7_7_chanxy_out[3];
    assign wire_9039 = lut_tile_7_7_chanxy_out[4];
    assign wire_9041 = lut_tile_7_7_chanxy_out[5];
    assign wire_9043 = lut_tile_7_7_chanxy_out[6];
    assign wire_9045 = lut_tile_7_7_chanxy_out[7];
    assign wire_9047 = lut_tile_7_7_chanxy_out[8];
    assign wire_9049 = lut_tile_7_7_chanxy_out[9];
    assign wire_9051 = lut_tile_7_7_chanxy_out[10];
    assign wire_9053 = lut_tile_7_7_chanxy_out[11];
    assign wire_9055 = lut_tile_7_7_chanxy_out[12];
    assign wire_9057 = lut_tile_7_7_chanxy_out[13];
    assign wire_9059 = lut_tile_7_7_chanxy_out[14];
    assign wire_9120 = lut_tile_7_7_chanxy_out[15];
    assign wire_9122 = lut_tile_7_7_chanxy_out[16];
    assign wire_9124 = lut_tile_7_7_chanxy_out[17];
    assign wire_9126 = lut_tile_7_7_chanxy_out[18];
    assign wire_9128 = lut_tile_7_7_chanxy_out[19];
    assign wire_9130 = lut_tile_7_7_chanxy_out[20];
    assign wire_9132 = lut_tile_7_7_chanxy_out[21];
    assign wire_9134 = lut_tile_7_7_chanxy_out[22];
    assign wire_9136 = lut_tile_7_7_chanxy_out[23];
    assign wire_9138 = lut_tile_7_7_chanxy_out[24];
    assign wire_9140 = lut_tile_7_7_chanxy_out[25];
    assign wire_9142 = lut_tile_7_7_chanxy_out[26];
    assign wire_9144 = lut_tile_7_7_chanxy_out[27];
    assign wire_9146 = lut_tile_7_7_chanxy_out[28];
    assign wire_9148 = lut_tile_7_7_chanxy_out[29];
    assign wire_13321 = lut_tile_7_7_chanxy_out[30];
    assign wire_13323 = lut_tile_7_7_chanxy_out[31];
    assign wire_13325 = lut_tile_7_7_chanxy_out[32];
    assign wire_13327 = lut_tile_7_7_chanxy_out[33];
    assign wire_13329 = lut_tile_7_7_chanxy_out[34];
    assign wire_13331 = lut_tile_7_7_chanxy_out[35];
    assign wire_13333 = lut_tile_7_7_chanxy_out[36];
    assign wire_13335 = lut_tile_7_7_chanxy_out[37];
    assign wire_13337 = lut_tile_7_7_chanxy_out[38];
    assign wire_13339 = lut_tile_7_7_chanxy_out[39];
    assign wire_13341 = lut_tile_7_7_chanxy_out[40];
    assign wire_13343 = lut_tile_7_7_chanxy_out[41];
    assign wire_13345 = lut_tile_7_7_chanxy_out[42];
    assign wire_13347 = lut_tile_7_7_chanxy_out[43];
    assign wire_13349 = lut_tile_7_7_chanxy_out[44];
    assign wire_13410 = lut_tile_7_7_chanxy_out[45];
    assign wire_13412 = lut_tile_7_7_chanxy_out[46];
    assign wire_13414 = lut_tile_7_7_chanxy_out[47];
    assign wire_13416 = lut_tile_7_7_chanxy_out[48];
    assign wire_13418 = lut_tile_7_7_chanxy_out[49];
    assign wire_13420 = lut_tile_7_7_chanxy_out[50];
    assign wire_13422 = lut_tile_7_7_chanxy_out[51];
    assign wire_13424 = lut_tile_7_7_chanxy_out[52];
    assign wire_13426 = lut_tile_7_7_chanxy_out[53];
    assign wire_13428 = lut_tile_7_7_chanxy_out[54];
    assign wire_13430 = lut_tile_7_7_chanxy_out[55];
    assign wire_13432 = lut_tile_7_7_chanxy_out[56];
    assign wire_13434 = lut_tile_7_7_chanxy_out[57];
    assign wire_13436 = lut_tile_7_7_chanxy_out[58];
    assign wire_13438 = lut_tile_7_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_8_chanxy_in = {wire_13708, wire_8791, wire_8729, wire_8728, wire_8719, wire_8718, wire_8709, wire_8708, wire_8672, wire_4941, wire_13706, wire_8819, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8674, wire_4941, wire_13704, wire_8817, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8676, wire_4941, wire_13702, wire_8815, wire_8727, wire_8726, wire_8717, wire_8716, wire_8707, wire_8706, wire_8678, wire_4431, wire_13700, wire_8813, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8680, wire_4431, wire_13698, wire_8811, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8682, wire_4431, wire_13696, wire_8809, wire_8725, wire_8724, wire_8715, wire_8714, wire_8705, wire_8704, wire_8684, wire_4945, wire_4431, wire_13694, wire_8807, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8686, wire_4945, wire_4431, wire_13692, wire_8805, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8688, wire_4945, wire_4431, wire_13690, wire_8803, wire_8723, wire_8722, wire_8713, wire_8712, wire_8703, wire_8702, wire_8690, wire_4945, wire_4427, wire_13688, wire_8801, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8692, wire_4945, wire_4427, wire_13686, wire_8799, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8694, wire_4945, wire_4427, wire_13684, wire_8797, wire_8721, wire_8720, wire_8711, wire_8710, wire_8701, wire_8700, wire_8696, wire_4941, wire_4427, wire_13682, wire_8795, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8698, wire_4941, wire_4427, wire_13680, wire_8793, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8670, wire_4941, wire_4427, wire_13859, wire_9209, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9060, wire_4941, wire_13857, wire_9181, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9088, wire_4941, wire_13855, wire_9183, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9086, wire_4941, wire_13853, wire_9185, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9084, wire_4431, wire_13851, wire_9187, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9082, wire_4431, wire_13849, wire_9189, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9080, wire_4431, wire_13847, wire_9191, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9078, wire_4945, wire_4431, wire_13845, wire_9193, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9076, wire_4945, wire_4431, wire_13843, wire_9195, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9074, wire_4945, wire_4431, wire_13841, wire_9197, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9072, wire_4945, wire_4427, wire_13839, wire_9199, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9070, wire_4945, wire_4427, wire_13837, wire_9201, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9068, wire_4945, wire_4427, wire_13835, wire_9203, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9066, wire_4941, wire_4427, wire_13833, wire_9205, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9064, wire_4941, wire_4427, wire_13831, wire_9207, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9062, wire_4941, wire_4427, wire_13467, wire_13379, wire_13378, wire_13369, wire_13368, wire_13359, wire_13358, wire_13348, wire_9058, wire_4470, wire_13465, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13320, wire_9056, wire_4470, wire_13463, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13322, wire_9054, wire_4470, wire_13461, wire_13377, wire_13376, wire_13367, wire_13366, wire_13357, wire_13356, wire_13324, wire_9052, wire_4430, wire_13459, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13326, wire_9050, wire_4430, wire_13457, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13328, wire_9048, wire_4430, wire_13455, wire_13375, wire_13374, wire_13365, wire_13364, wire_13355, wire_13354, wire_13330, wire_9046, wire_4474, wire_4430, wire_13453, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13332, wire_9044, wire_4474, wire_4430, wire_13451, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13334, wire_9042, wire_4474, wire_4430, wire_13449, wire_13373, wire_13372, wire_13363, wire_13362, wire_13353, wire_13352, wire_13336, wire_9040, wire_4474, wire_4426, wire_13447, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13338, wire_9038, wire_4474, wire_4426, wire_13445, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13340, wire_9036, wire_4474, wire_4426, wire_13443, wire_13371, wire_13370, wire_13361, wire_13360, wire_13351, wire_13350, wire_13342, wire_9034, wire_4470, wire_4426, wire_13441, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13344, wire_9032, wire_4470, wire_4426, wire_13469, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13346, wire_9030, wire_4470, wire_4426, wire_13833, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13736, wire_9209, wire_4470, wire_13835, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13734, wire_9207, wire_4470, wire_13837, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13732, wire_9205, wire_4470, wire_13839, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13730, wire_9203, wire_4430, wire_13841, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13728, wire_9201, wire_4430, wire_13843, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13726, wire_9199, wire_4430, wire_13845, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13724, wire_9197, wire_4474, wire_4430, wire_13847, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13722, wire_9195, wire_4474, wire_4430, wire_13849, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13720, wire_9193, wire_4474, wire_4430, wire_13851, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13718, wire_9191, wire_4474, wire_4426, wire_13853, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13716, wire_9189, wire_4474, wire_4426, wire_13855, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13714, wire_9187, wire_4474, wire_4426, wire_13857, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13712, wire_9185, wire_4470, wire_4426, wire_13859, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13710, wire_9183, wire_4470, wire_4426, wire_13831, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13738, wire_9181, wire_4470, wire_4426};
    // CHNAXY TOTAL: 636
    assign wire_9061 = lut_tile_7_8_chanxy_out[0];
    assign wire_9063 = lut_tile_7_8_chanxy_out[1];
    assign wire_9065 = lut_tile_7_8_chanxy_out[2];
    assign wire_9067 = lut_tile_7_8_chanxy_out[3];
    assign wire_9069 = lut_tile_7_8_chanxy_out[4];
    assign wire_9071 = lut_tile_7_8_chanxy_out[5];
    assign wire_9073 = lut_tile_7_8_chanxy_out[6];
    assign wire_9075 = lut_tile_7_8_chanxy_out[7];
    assign wire_9077 = lut_tile_7_8_chanxy_out[8];
    assign wire_9079 = lut_tile_7_8_chanxy_out[9];
    assign wire_9081 = lut_tile_7_8_chanxy_out[10];
    assign wire_9083 = lut_tile_7_8_chanxy_out[11];
    assign wire_9085 = lut_tile_7_8_chanxy_out[12];
    assign wire_9087 = lut_tile_7_8_chanxy_out[13];
    assign wire_9089 = lut_tile_7_8_chanxy_out[14];
    assign wire_9150 = lut_tile_7_8_chanxy_out[15];
    assign wire_9152 = lut_tile_7_8_chanxy_out[16];
    assign wire_9154 = lut_tile_7_8_chanxy_out[17];
    assign wire_9156 = lut_tile_7_8_chanxy_out[18];
    assign wire_9158 = lut_tile_7_8_chanxy_out[19];
    assign wire_9160 = lut_tile_7_8_chanxy_out[20];
    assign wire_9162 = lut_tile_7_8_chanxy_out[21];
    assign wire_9164 = lut_tile_7_8_chanxy_out[22];
    assign wire_9166 = lut_tile_7_8_chanxy_out[23];
    assign wire_9168 = lut_tile_7_8_chanxy_out[24];
    assign wire_9170 = lut_tile_7_8_chanxy_out[25];
    assign wire_9172 = lut_tile_7_8_chanxy_out[26];
    assign wire_9174 = lut_tile_7_8_chanxy_out[27];
    assign wire_9176 = lut_tile_7_8_chanxy_out[28];
    assign wire_9178 = lut_tile_7_8_chanxy_out[29];
    assign wire_13711 = lut_tile_7_8_chanxy_out[30];
    assign wire_13713 = lut_tile_7_8_chanxy_out[31];
    assign wire_13715 = lut_tile_7_8_chanxy_out[32];
    assign wire_13717 = lut_tile_7_8_chanxy_out[33];
    assign wire_13719 = lut_tile_7_8_chanxy_out[34];
    assign wire_13721 = lut_tile_7_8_chanxy_out[35];
    assign wire_13723 = lut_tile_7_8_chanxy_out[36];
    assign wire_13725 = lut_tile_7_8_chanxy_out[37];
    assign wire_13727 = lut_tile_7_8_chanxy_out[38];
    assign wire_13729 = lut_tile_7_8_chanxy_out[39];
    assign wire_13731 = lut_tile_7_8_chanxy_out[40];
    assign wire_13733 = lut_tile_7_8_chanxy_out[41];
    assign wire_13735 = lut_tile_7_8_chanxy_out[42];
    assign wire_13737 = lut_tile_7_8_chanxy_out[43];
    assign wire_13739 = lut_tile_7_8_chanxy_out[44];
    assign wire_13800 = lut_tile_7_8_chanxy_out[45];
    assign wire_13802 = lut_tile_7_8_chanxy_out[46];
    assign wire_13804 = lut_tile_7_8_chanxy_out[47];
    assign wire_13806 = lut_tile_7_8_chanxy_out[48];
    assign wire_13808 = lut_tile_7_8_chanxy_out[49];
    assign wire_13810 = lut_tile_7_8_chanxy_out[50];
    assign wire_13812 = lut_tile_7_8_chanxy_out[51];
    assign wire_13814 = lut_tile_7_8_chanxy_out[52];
    assign wire_13816 = lut_tile_7_8_chanxy_out[53];
    assign wire_13818 = lut_tile_7_8_chanxy_out[54];
    assign wire_13820 = lut_tile_7_8_chanxy_out[55];
    assign wire_13822 = lut_tile_7_8_chanxy_out[56];
    assign wire_13824 = lut_tile_7_8_chanxy_out[57];
    assign wire_13826 = lut_tile_7_8_chanxy_out[58];
    assign wire_13828 = lut_tile_7_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_9_chanxy_in = {wire_14098, wire_8821, wire_8819, wire_8818, wire_8809, wire_8808, wire_8799, wire_8798, wire_8702, wire_5457, wire_14096, wire_8849, wire_8789, wire_8788, wire_8779, wire_8778, wire_8769, wire_8768, wire_8704, wire_5457, wire_14094, wire_8847, wire_8759, wire_8758, wire_8749, wire_8748, wire_8739, wire_8738, wire_8706, wire_5457, wire_14092, wire_8845, wire_8817, wire_8816, wire_8807, wire_8806, wire_8797, wire_8796, wire_8708, wire_4947, wire_14090, wire_8843, wire_8787, wire_8786, wire_8777, wire_8776, wire_8767, wire_8766, wire_8710, wire_4947, wire_14088, wire_8841, wire_8757, wire_8756, wire_8747, wire_8746, wire_8737, wire_8736, wire_8712, wire_4947, wire_14086, wire_8839, wire_8815, wire_8814, wire_8805, wire_8804, wire_8795, wire_8794, wire_8714, wire_5461, wire_4947, wire_14084, wire_8837, wire_8785, wire_8784, wire_8775, wire_8774, wire_8765, wire_8764, wire_8716, wire_5461, wire_4947, wire_14082, wire_8835, wire_8755, wire_8754, wire_8745, wire_8744, wire_8735, wire_8734, wire_8718, wire_5461, wire_4947, wire_14080, wire_8833, wire_8813, wire_8812, wire_8803, wire_8802, wire_8793, wire_8792, wire_8720, wire_5461, wire_4943, wire_14078, wire_8831, wire_8783, wire_8782, wire_8773, wire_8772, wire_8763, wire_8762, wire_8722, wire_5461, wire_4943, wire_14076, wire_8829, wire_8753, wire_8752, wire_8743, wire_8742, wire_8733, wire_8732, wire_8724, wire_5461, wire_4943, wire_14074, wire_8827, wire_8811, wire_8810, wire_8801, wire_8800, wire_8791, wire_8790, wire_8726, wire_5457, wire_4943, wire_14072, wire_8825, wire_8781, wire_8780, wire_8771, wire_8770, wire_8761, wire_8760, wire_8728, wire_5457, wire_4943, wire_14070, wire_8823, wire_8751, wire_8750, wire_8741, wire_8740, wire_8731, wire_8730, wire_8700, wire_5457, wire_4943, wire_14249, wire_9239, wire_9209, wire_9208, wire_9199, wire_9198, wire_9189, wire_9188, wire_9090, wire_5457, wire_14247, wire_9211, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9118, wire_5457, wire_14245, wire_9213, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9116, wire_5457, wire_14243, wire_9215, wire_9207, wire_9206, wire_9197, wire_9196, wire_9187, wire_9186, wire_9114, wire_4947, wire_14241, wire_9217, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9112, wire_4947, wire_14239, wire_9219, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9110, wire_4947, wire_14237, wire_9221, wire_9205, wire_9204, wire_9195, wire_9194, wire_9185, wire_9184, wire_9108, wire_5461, wire_4947, wire_14235, wire_9223, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9106, wire_5461, wire_4947, wire_14233, wire_9225, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9104, wire_5461, wire_4947, wire_14231, wire_9227, wire_9203, wire_9202, wire_9193, wire_9192, wire_9183, wire_9182, wire_9102, wire_5461, wire_4943, wire_14229, wire_9229, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9100, wire_5461, wire_4943, wire_14227, wire_9231, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9098, wire_5461, wire_4943, wire_14225, wire_9233, wire_9201, wire_9200, wire_9191, wire_9190, wire_9181, wire_9180, wire_9096, wire_5457, wire_4943, wire_14223, wire_9235, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9094, wire_5457, wire_4943, wire_14221, wire_9237, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9092, wire_5457, wire_4943, wire_13857, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13738, wire_9088, wire_4986, wire_13855, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13710, wire_9086, wire_4986, wire_13853, wire_13769, wire_13768, wire_13759, wire_13758, wire_13749, wire_13748, wire_13712, wire_9084, wire_4986, wire_13851, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13714, wire_9082, wire_4946, wire_13849, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13716, wire_9080, wire_4946, wire_13847, wire_13767, wire_13766, wire_13757, wire_13756, wire_13747, wire_13746, wire_13718, wire_9078, wire_4946, wire_13845, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13720, wire_9076, wire_4990, wire_4946, wire_13843, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13722, wire_9074, wire_4990, wire_4946, wire_13841, wire_13765, wire_13764, wire_13755, wire_13754, wire_13745, wire_13744, wire_13724, wire_9072, wire_4990, wire_4946, wire_13839, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13726, wire_9070, wire_4990, wire_4942, wire_13837, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13728, wire_9068, wire_4990, wire_4942, wire_13835, wire_13763, wire_13762, wire_13753, wire_13752, wire_13743, wire_13742, wire_13730, wire_9066, wire_4990, wire_4942, wire_13833, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13732, wire_9064, wire_4986, wire_4942, wire_13831, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13734, wire_9062, wire_4986, wire_4942, wire_13859, wire_13761, wire_13760, wire_13751, wire_13750, wire_13741, wire_13740, wire_13736, wire_9060, wire_4986, wire_4942, wire_14223, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14126, wire_9239, wire_4986, wire_14225, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14124, wire_9237, wire_4986, wire_14227, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14122, wire_9235, wire_4986, wire_14229, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14120, wire_9233, wire_4946, wire_14231, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14118, wire_9231, wire_4946, wire_14233, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14116, wire_9229, wire_4946, wire_14235, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14114, wire_9227, wire_4990, wire_4946, wire_14237, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14112, wire_9225, wire_4990, wire_4946, wire_14239, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14110, wire_9223, wire_4990, wire_4946, wire_14241, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14108, wire_9221, wire_4990, wire_4942, wire_14243, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14106, wire_9219, wire_4990, wire_4942, wire_14245, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14104, wire_9217, wire_4990, wire_4942, wire_14247, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14102, wire_9215, wire_4986, wire_4942, wire_14249, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14100, wire_9213, wire_4986, wire_4942, wire_14221, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14128, wire_9211, wire_4986, wire_4942};
    // CHNAXY TOTAL: 636
    assign wire_9091 = lut_tile_7_9_chanxy_out[0];
    assign wire_9093 = lut_tile_7_9_chanxy_out[1];
    assign wire_9095 = lut_tile_7_9_chanxy_out[2];
    assign wire_9097 = lut_tile_7_9_chanxy_out[3];
    assign wire_9099 = lut_tile_7_9_chanxy_out[4];
    assign wire_9101 = lut_tile_7_9_chanxy_out[5];
    assign wire_9103 = lut_tile_7_9_chanxy_out[6];
    assign wire_9105 = lut_tile_7_9_chanxy_out[7];
    assign wire_9107 = lut_tile_7_9_chanxy_out[8];
    assign wire_9109 = lut_tile_7_9_chanxy_out[9];
    assign wire_9111 = lut_tile_7_9_chanxy_out[10];
    assign wire_9113 = lut_tile_7_9_chanxy_out[11];
    assign wire_9115 = lut_tile_7_9_chanxy_out[12];
    assign wire_9117 = lut_tile_7_9_chanxy_out[13];
    assign wire_9119 = lut_tile_7_9_chanxy_out[14];
    assign wire_9180 = lut_tile_7_9_chanxy_out[15];
    assign wire_9182 = lut_tile_7_9_chanxy_out[16];
    assign wire_9184 = lut_tile_7_9_chanxy_out[17];
    assign wire_9186 = lut_tile_7_9_chanxy_out[18];
    assign wire_9188 = lut_tile_7_9_chanxy_out[19];
    assign wire_9190 = lut_tile_7_9_chanxy_out[20];
    assign wire_9192 = lut_tile_7_9_chanxy_out[21];
    assign wire_9194 = lut_tile_7_9_chanxy_out[22];
    assign wire_9196 = lut_tile_7_9_chanxy_out[23];
    assign wire_9198 = lut_tile_7_9_chanxy_out[24];
    assign wire_9200 = lut_tile_7_9_chanxy_out[25];
    assign wire_9202 = lut_tile_7_9_chanxy_out[26];
    assign wire_9204 = lut_tile_7_9_chanxy_out[27];
    assign wire_9206 = lut_tile_7_9_chanxy_out[28];
    assign wire_9208 = lut_tile_7_9_chanxy_out[29];
    assign wire_14101 = lut_tile_7_9_chanxy_out[30];
    assign wire_14103 = lut_tile_7_9_chanxy_out[31];
    assign wire_14105 = lut_tile_7_9_chanxy_out[32];
    assign wire_14107 = lut_tile_7_9_chanxy_out[33];
    assign wire_14109 = lut_tile_7_9_chanxy_out[34];
    assign wire_14111 = lut_tile_7_9_chanxy_out[35];
    assign wire_14113 = lut_tile_7_9_chanxy_out[36];
    assign wire_14115 = lut_tile_7_9_chanxy_out[37];
    assign wire_14117 = lut_tile_7_9_chanxy_out[38];
    assign wire_14119 = lut_tile_7_9_chanxy_out[39];
    assign wire_14121 = lut_tile_7_9_chanxy_out[40];
    assign wire_14123 = lut_tile_7_9_chanxy_out[41];
    assign wire_14125 = lut_tile_7_9_chanxy_out[42];
    assign wire_14127 = lut_tile_7_9_chanxy_out[43];
    assign wire_14129 = lut_tile_7_9_chanxy_out[44];
    assign wire_14190 = lut_tile_7_9_chanxy_out[45];
    assign wire_14192 = lut_tile_7_9_chanxy_out[46];
    assign wire_14194 = lut_tile_7_9_chanxy_out[47];
    assign wire_14196 = lut_tile_7_9_chanxy_out[48];
    assign wire_14198 = lut_tile_7_9_chanxy_out[49];
    assign wire_14200 = lut_tile_7_9_chanxy_out[50];
    assign wire_14202 = lut_tile_7_9_chanxy_out[51];
    assign wire_14204 = lut_tile_7_9_chanxy_out[52];
    assign wire_14206 = lut_tile_7_9_chanxy_out[53];
    assign wire_14208 = lut_tile_7_9_chanxy_out[54];
    assign wire_14210 = lut_tile_7_9_chanxy_out[55];
    assign wire_14212 = lut_tile_7_9_chanxy_out[56];
    assign wire_14214 = lut_tile_7_9_chanxy_out[57];
    assign wire_14216 = lut_tile_7_9_chanxy_out[58];
    assign wire_14218 = lut_tile_7_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_7_10_chanxy_in = {wire_14488, wire_8848, wire_8796, wire_8774, wire_8752, wire_5974, wire_5968, wire_5959, wire_5953, wire_14486, wire_8840, wire_8818, wire_8766, wire_8744, wire_5974, wire_5968, wire_5959, wire_5953, wire_14484, wire_8832, wire_8810, wire_8788, wire_8736, wire_5974, wire_5968, wire_5959, wire_5953, wire_14482, wire_8824, wire_8802, wire_8780, wire_8758, wire_5974, wire_5965, wire_5959, wire_5463, wire_14480, wire_8846, wire_8794, wire_8772, wire_8750, wire_5974, wire_5965, wire_5959, wire_5463, wire_14478, wire_8838, wire_8816, wire_8764, wire_8742, wire_5974, wire_5965, wire_5959, wire_5463, wire_14476, wire_8830, wire_8808, wire_8786, wire_8734, wire_5971, wire_5965, wire_5956, wire_5463, wire_14474, wire_8822, wire_8800, wire_8778, wire_8756, wire_5971, wire_5965, wire_5956, wire_5463, wire_14472, wire_8844, wire_8792, wire_8770, wire_8748, wire_5971, wire_5965, wire_5956, wire_5463, wire_14470, wire_8836, wire_8814, wire_8762, wire_8740, wire_5971, wire_5962, wire_5956, wire_5459, wire_14468, wire_8828, wire_8806, wire_8784, wire_8732, wire_5971, wire_5962, wire_5956, wire_5459, wire_14466, wire_8820, wire_8798, wire_8776, wire_8754, wire_5971, wire_5962, wire_5956, wire_5459, wire_14464, wire_8842, wire_8790, wire_8768, wire_8746, wire_5968, wire_5962, wire_5953, wire_5459, wire_14462, wire_8834, wire_8812, wire_8760, wire_8738, wire_5968, wire_5962, wire_5953, wire_5459, wire_14460, wire_8826, wire_8804, wire_8782, wire_8730, wire_5968, wire_5962, wire_5953, wire_5459, wire_14639, wire_9232, wire_9208, wire_9156, wire_9134, wire_5974, wire_5968, wire_5959, wire_5953, wire_14637, wire_9224, wire_9200, wire_9178, wire_9126, wire_5974, wire_5968, wire_5959, wire_5953, wire_14635, wire_9216, wire_9192, wire_9170, wire_9148, wire_5974, wire_5968, wire_5959, wire_5953, wire_14633, wire_9238, wire_9184, wire_9162, wire_9140, wire_5974, wire_5965, wire_5959, wire_5463, wire_14631, wire_9230, wire_9206, wire_9154, wire_9132, wire_5974, wire_5965, wire_5959, wire_5463, wire_14629, wire_9222, wire_9198, wire_9176, wire_9124, wire_5974, wire_5965, wire_5959, wire_5463, wire_14627, wire_9214, wire_9190, wire_9168, wire_9146, wire_5971, wire_5965, wire_5956, wire_5463, wire_14625, wire_9236, wire_9182, wire_9160, wire_9138, wire_5971, wire_5965, wire_5956, wire_5463, wire_14623, wire_9228, wire_9204, wire_9152, wire_9130, wire_5971, wire_5965, wire_5956, wire_5463, wire_14621, wire_9220, wire_9196, wire_9174, wire_9122, wire_5971, wire_5962, wire_5956, wire_5459, wire_14619, wire_9212, wire_9188, wire_9166, wire_9144, wire_5971, wire_5962, wire_5956, wire_5459, wire_14617, wire_9234, wire_9180, wire_9158, wire_9136, wire_5971, wire_5962, wire_5956, wire_5459, wire_14615, wire_9226, wire_9202, wire_9150, wire_9128, wire_5968, wire_5962, wire_5953, wire_5459, wire_14613, wire_9218, wire_9194, wire_9172, wire_9120, wire_5968, wire_5962, wire_5953, wire_5459, wire_14611, wire_9210, wire_9186, wire_9164, wire_9142, wire_5968, wire_5962, wire_5953, wire_5459, wire_14639, wire_14518, wire_14247, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14128, wire_9118, wire_5502, wire_14547, wire_14546, wire_14245, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14100, wire_9116, wire_5502, wire_14593, wire_14592, wire_14243, wire_14159, wire_14158, wire_14149, wire_14148, wire_14139, wire_14138, wire_14102, wire_9114, wire_5502, wire_14621, wire_14500, wire_14241, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14104, wire_9112, wire_5462, wire_14529, wire_14528, wire_14239, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14106, wire_9110, wire_5462, wire_14605, wire_14604, wire_14237, wire_14157, wire_14156, wire_14147, wire_14146, wire_14137, wire_14136, wire_14108, wire_9108, wire_5462, wire_14633, wire_14512, wire_14235, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14110, wire_9106, wire_5506, wire_5462, wire_14541, wire_14540, wire_14233, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14112, wire_9104, wire_5506, wire_5462, wire_14587, wire_14586, wire_14231, wire_14155, wire_14154, wire_14145, wire_14144, wire_14135, wire_14134, wire_14114, wire_9102, wire_5506, wire_5462, wire_14615, wire_14494, wire_5506, wire_14229, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14116, wire_9100, wire_5506, wire_5458, wire_14523, wire_14522, wire_5502, wire_14227, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14118, wire_9098, wire_5506, wire_5458, wire_14599, wire_14598, wire_5502, wire_14225, wire_14153, wire_14152, wire_14143, wire_14142, wire_14133, wire_14132, wire_14120, wire_9096, wire_5506, wire_5458, wire_14627, wire_14506, wire_5462, wire_14223, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14122, wire_9094, wire_5502, wire_5458, wire_14535, wire_14534, wire_5458, wire_14221, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14124, wire_9092, wire_5502, wire_5458, wire_14581, wire_14580, wire_5458, wire_14249, wire_14151, wire_14150, wire_14141, wire_14140, wire_14131, wire_14130, wire_14126, wire_9090, wire_5502, wire_5458, wire_14579, wire_14578, wire_14609, wire_14608, wire_14623, wire_14502, wire_14561, wire_14560, wire_14591, wire_14590, wire_14635, wire_14514, wire_14573, wire_14572, wire_14603, wire_14602, wire_14617, wire_14496, wire_14555, wire_14554, wire_5506, wire_14585, wire_14584, wire_5506, wire_14629, wire_14508, wire_5502, wire_14567, wire_14566, wire_5462, wire_14597, wire_14596, wire_5462, wire_14611, wire_14490, wire_5458, wire_14549, wire_14548, wire_14533, wire_14532, wire_14637, wire_14516, wire_14531, wire_14530, wire_14545, wire_14544, wire_14619, wire_14498, wire_14543, wire_14542, wire_14527, wire_14526, wire_14631, wire_14510, wire_14525, wire_14524, wire_5506, wire_14539, wire_14538, wire_5506, wire_14613, wire_14492, wire_5502, wire_14537, wire_14536, wire_5462, wire_14521, wire_14520, wire_5462, wire_14625, wire_14504, wire_5458, wire_14563, wire_14562, wire_14577, wire_14576, wire_14607, wire_14606, wire_14575, wire_14574, wire_14559, wire_14558, wire_14589, wire_14588, wire_14557, wire_14556, wire_14571, wire_14570, wire_14601, wire_14600, wire_14569, wire_14568, wire_5506, wire_14553, wire_14552, wire_5502, wire_14583, wire_14582, wire_5502, wire_14551, wire_14550, wire_5462, wire_14565, wire_14564, wire_5458, wire_14595, wire_14594, wire_5458};
    // CHNAXY TOTAL: 573
    assign wire_9121 = lut_tile_7_10_chanxy_out[0];
    assign wire_9123 = lut_tile_7_10_chanxy_out[1];
    assign wire_9125 = lut_tile_7_10_chanxy_out[2];
    assign wire_9127 = lut_tile_7_10_chanxy_out[3];
    assign wire_9129 = lut_tile_7_10_chanxy_out[4];
    assign wire_9131 = lut_tile_7_10_chanxy_out[5];
    assign wire_9133 = lut_tile_7_10_chanxy_out[6];
    assign wire_9135 = lut_tile_7_10_chanxy_out[7];
    assign wire_9137 = lut_tile_7_10_chanxy_out[8];
    assign wire_9139 = lut_tile_7_10_chanxy_out[9];
    assign wire_9141 = lut_tile_7_10_chanxy_out[10];
    assign wire_9143 = lut_tile_7_10_chanxy_out[11];
    assign wire_9145 = lut_tile_7_10_chanxy_out[12];
    assign wire_9147 = lut_tile_7_10_chanxy_out[13];
    assign wire_9149 = lut_tile_7_10_chanxy_out[14];
    assign wire_9151 = lut_tile_7_10_chanxy_out[15];
    assign wire_9153 = lut_tile_7_10_chanxy_out[16];
    assign wire_9155 = lut_tile_7_10_chanxy_out[17];
    assign wire_9157 = lut_tile_7_10_chanxy_out[18];
    assign wire_9159 = lut_tile_7_10_chanxy_out[19];
    assign wire_9161 = lut_tile_7_10_chanxy_out[20];
    assign wire_9163 = lut_tile_7_10_chanxy_out[21];
    assign wire_9165 = lut_tile_7_10_chanxy_out[22];
    assign wire_9167 = lut_tile_7_10_chanxy_out[23];
    assign wire_9169 = lut_tile_7_10_chanxy_out[24];
    assign wire_9171 = lut_tile_7_10_chanxy_out[25];
    assign wire_9173 = lut_tile_7_10_chanxy_out[26];
    assign wire_9175 = lut_tile_7_10_chanxy_out[27];
    assign wire_9177 = lut_tile_7_10_chanxy_out[28];
    assign wire_9179 = lut_tile_7_10_chanxy_out[29];
    assign wire_9181 = lut_tile_7_10_chanxy_out[30];
    assign wire_9183 = lut_tile_7_10_chanxy_out[31];
    assign wire_9185 = lut_tile_7_10_chanxy_out[32];
    assign wire_9187 = lut_tile_7_10_chanxy_out[33];
    assign wire_9189 = lut_tile_7_10_chanxy_out[34];
    assign wire_9191 = lut_tile_7_10_chanxy_out[35];
    assign wire_9193 = lut_tile_7_10_chanxy_out[36];
    assign wire_9195 = lut_tile_7_10_chanxy_out[37];
    assign wire_9197 = lut_tile_7_10_chanxy_out[38];
    assign wire_9199 = lut_tile_7_10_chanxy_out[39];
    assign wire_9201 = lut_tile_7_10_chanxy_out[40];
    assign wire_9203 = lut_tile_7_10_chanxy_out[41];
    assign wire_9205 = lut_tile_7_10_chanxy_out[42];
    assign wire_9207 = lut_tile_7_10_chanxy_out[43];
    assign wire_9209 = lut_tile_7_10_chanxy_out[44];
    assign wire_9210 = lut_tile_7_10_chanxy_out[45];
    assign wire_9211 = lut_tile_7_10_chanxy_out[46];
    assign wire_9212 = lut_tile_7_10_chanxy_out[47];
    assign wire_9213 = lut_tile_7_10_chanxy_out[48];
    assign wire_9214 = lut_tile_7_10_chanxy_out[49];
    assign wire_9215 = lut_tile_7_10_chanxy_out[50];
    assign wire_9216 = lut_tile_7_10_chanxy_out[51];
    assign wire_9217 = lut_tile_7_10_chanxy_out[52];
    assign wire_9218 = lut_tile_7_10_chanxy_out[53];
    assign wire_9219 = lut_tile_7_10_chanxy_out[54];
    assign wire_9220 = lut_tile_7_10_chanxy_out[55];
    assign wire_9221 = lut_tile_7_10_chanxy_out[56];
    assign wire_9222 = lut_tile_7_10_chanxy_out[57];
    assign wire_9223 = lut_tile_7_10_chanxy_out[58];
    assign wire_9224 = lut_tile_7_10_chanxy_out[59];
    assign wire_9225 = lut_tile_7_10_chanxy_out[60];
    assign wire_9226 = lut_tile_7_10_chanxy_out[61];
    assign wire_9227 = lut_tile_7_10_chanxy_out[62];
    assign wire_9228 = lut_tile_7_10_chanxy_out[63];
    assign wire_9229 = lut_tile_7_10_chanxy_out[64];
    assign wire_9230 = lut_tile_7_10_chanxy_out[65];
    assign wire_9231 = lut_tile_7_10_chanxy_out[66];
    assign wire_9232 = lut_tile_7_10_chanxy_out[67];
    assign wire_9233 = lut_tile_7_10_chanxy_out[68];
    assign wire_9234 = lut_tile_7_10_chanxy_out[69];
    assign wire_9235 = lut_tile_7_10_chanxy_out[70];
    assign wire_9236 = lut_tile_7_10_chanxy_out[71];
    assign wire_9237 = lut_tile_7_10_chanxy_out[72];
    assign wire_9238 = lut_tile_7_10_chanxy_out[73];
    assign wire_9239 = lut_tile_7_10_chanxy_out[74];
    assign wire_14491 = lut_tile_7_10_chanxy_out[75];
    assign wire_14493 = lut_tile_7_10_chanxy_out[76];
    assign wire_14495 = lut_tile_7_10_chanxy_out[77];
    assign wire_14497 = lut_tile_7_10_chanxy_out[78];
    assign wire_14499 = lut_tile_7_10_chanxy_out[79];
    assign wire_14501 = lut_tile_7_10_chanxy_out[80];
    assign wire_14503 = lut_tile_7_10_chanxy_out[81];
    assign wire_14505 = lut_tile_7_10_chanxy_out[82];
    assign wire_14507 = lut_tile_7_10_chanxy_out[83];
    assign wire_14509 = lut_tile_7_10_chanxy_out[84];
    assign wire_14511 = lut_tile_7_10_chanxy_out[85];
    assign wire_14513 = lut_tile_7_10_chanxy_out[86];
    assign wire_14515 = lut_tile_7_10_chanxy_out[87];
    assign wire_14517 = lut_tile_7_10_chanxy_out[88];
    assign wire_14519 = lut_tile_7_10_chanxy_out[89];
    assign wire_14580 = lut_tile_7_10_chanxy_out[90];
    assign wire_14582 = lut_tile_7_10_chanxy_out[91];
    assign wire_14584 = lut_tile_7_10_chanxy_out[92];
    assign wire_14586 = lut_tile_7_10_chanxy_out[93];
    assign wire_14588 = lut_tile_7_10_chanxy_out[94];
    assign wire_14590 = lut_tile_7_10_chanxy_out[95];
    assign wire_14592 = lut_tile_7_10_chanxy_out[96];
    assign wire_14594 = lut_tile_7_10_chanxy_out[97];
    assign wire_14596 = lut_tile_7_10_chanxy_out[98];
    assign wire_14598 = lut_tile_7_10_chanxy_out[99];
    assign wire_14600 = lut_tile_7_10_chanxy_out[100];
    assign wire_14602 = lut_tile_7_10_chanxy_out[101];
    assign wire_14604 = lut_tile_7_10_chanxy_out[102];
    assign wire_14606 = lut_tile_7_10_chanxy_out[103];
    assign wire_14608 = lut_tile_7_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_8_1_chanxy_in = {wire_11008, wire_8971, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8858, wire_1371, wire_11006, wire_8999, wire_8967, wire_8966, wire_8927, wire_8926, wire_8887, wire_8886, wire_8866, wire_1371, wire_11004, wire_8997, wire_8965, wire_8964, wire_8925, wire_8924, wire_8885, wire_8884, wire_8874, wire_1371, wire_11002, wire_8995, wire_8961, wire_8960, wire_8921, wire_8920, wire_8882, wire_8881, wire_8880, wire_861, wire_11000, wire_8993, wire_8959, wire_8958, wire_8919, wire_8918, wire_8890, wire_8879, wire_8878, wire_861, wire_10998, wire_8991, wire_8957, wire_8956, wire_8917, wire_8916, wire_8898, wire_8877, wire_8876, wire_861, wire_10996, wire_8989, wire_8953, wire_8952, wire_8913, wire_8912, wire_8906, wire_8873, wire_8872, wire_1375, wire_861, wire_10994, wire_8987, wire_8951, wire_8950, wire_8914, wire_8911, wire_8910, wire_8871, wire_8870, wire_1375, wire_861, wire_10992, wire_8985, wire_8949, wire_8948, wire_8922, wire_8909, wire_8908, wire_8869, wire_8868, wire_1375, wire_861, wire_10990, wire_8983, wire_8945, wire_8944, wire_8930, wire_8905, wire_8904, wire_8865, wire_8864, wire_1375, wire_857, wire_10988, wire_8981, wire_8943, wire_8942, wire_8938, wire_8903, wire_8902, wire_8863, wire_8862, wire_1375, wire_857, wire_10986, wire_8979, wire_8946, wire_8941, wire_8940, wire_8901, wire_8900, wire_8861, wire_8860, wire_1375, wire_857, wire_10984, wire_8977, wire_8954, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856, wire_1371, wire_857, wire_10982, wire_8975, wire_8962, wire_8935, wire_8934, wire_8895, wire_8894, wire_8855, wire_8854, wire_1371, wire_857, wire_10980, wire_8973, wire_8933, wire_8932, wire_8893, wire_8892, wire_8853, wire_8852, wire_8850, wire_1371, wire_857, wire_11159, wire_9389, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_9242, wire_1371, wire_11157, wire_9361, wire_9357, wire_9356, wire_9354, wire_9317, wire_9316, wire_9277, wire_9276, wire_1371, wire_11155, wire_9363, wire_9353, wire_9352, wire_9346, wire_9313, wire_9312, wire_9273, wire_9272, wire_1371, wire_11153, wire_9365, wire_9351, wire_9350, wire_9338, wire_9311, wire_9310, wire_9271, wire_9270, wire_861, wire_11151, wire_9367, wire_9349, wire_9348, wire_9330, wire_9309, wire_9308, wire_9269, wire_9268, wire_861, wire_11149, wire_9369, wire_9345, wire_9344, wire_9322, wire_9305, wire_9304, wire_9265, wire_9264, wire_861, wire_11147, wire_9371, wire_9343, wire_9342, wire_9314, wire_9303, wire_9302, wire_9263, wire_9262, wire_1375, wire_861, wire_11145, wire_9373, wire_9341, wire_9340, wire_9306, wire_9301, wire_9300, wire_9261, wire_9260, wire_1375, wire_861, wire_11143, wire_9375, wire_9337, wire_9336, wire_9298, wire_9297, wire_9296, wire_9257, wire_9256, wire_1375, wire_861, wire_11141, wire_9377, wire_9335, wire_9334, wire_9295, wire_9294, wire_9290, wire_9255, wire_9254, wire_1375, wire_857, wire_11139, wire_9379, wire_9333, wire_9332, wire_9293, wire_9292, wire_9282, wire_9253, wire_9252, wire_1375, wire_857, wire_11137, wire_9381, wire_9329, wire_9328, wire_9289, wire_9288, wire_9274, wire_9249, wire_9248, wire_1375, wire_857, wire_11135, wire_9383, wire_9327, wire_9326, wire_9287, wire_9286, wire_9266, wire_9247, wire_9246, wire_1371, wire_857, wire_11133, wire_9385, wire_9325, wire_9324, wire_9285, wire_9284, wire_9258, wire_9245, wire_9244, wire_1371, wire_857, wire_11131, wire_9387, wire_9321, wire_9320, wire_9281, wire_9280, wire_9250, wire_9241, wire_9240, wire_1371, wire_857, wire_10723, wire_10722, wire_10739, wire_10738, wire_11133, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11036, wire_9389, wire_900, wire_10709, wire_10708, wire_10693, wire_10692, wire_10679, wire_10678, wire_10769, wire_10648, wire_11135, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_11034, wire_9387, wire_900, wire_10663, wire_10662, wire_10737, wire_10736, wire_10707, wire_10706, wire_10753, wire_10632, wire_11137, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11032, wire_9385, wire_900, wire_10677, wire_10676, wire_10767, wire_10646, wire_10735, wire_10734, wire_10721, wire_10720, wire_11139, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11030, wire_9383, wire_860, wire_10691, wire_10690, wire_10705, wire_10704, wire_10661, wire_10660, wire_10751, wire_10630, wire_11141, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_11028, wire_9381, wire_860, wire_10675, wire_10674, wire_10719, wire_10718, wire_10689, wire_10688, wire_10765, wire_10644, wire_11143, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11026, wire_9379, wire_860, wire_10659, wire_10658, wire_10749, wire_10628, wire_10717, wire_10716, wire_10733, wire_10732, wire_11145, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11024, wire_9377, wire_904, wire_860, wire_10703, wire_10702, wire_10687, wire_10686, wire_10673, wire_10672, wire_10763, wire_10642, wire_11147, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_11022, wire_9375, wire_904, wire_860, wire_10657, wire_10656, wire_10731, wire_10730, wire_10701, wire_10700, wire_10747, wire_10626, wire_11149, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11020, wire_9373, wire_904, wire_860, wire_10671, wire_10670, wire_10761, wire_10640, wire_10729, wire_10728, wire_904, wire_10715, wire_10714, wire_904, wire_11151, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11018, wire_9371, wire_904, wire_856, wire_10685, wire_10684, wire_904, wire_10699, wire_10698, wire_904, wire_10655, wire_10654, wire_904, wire_10745, wire_10624, wire_904, wire_11153, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_11016, wire_9369, wire_904, wire_856, wire_10669, wire_10668, wire_900, wire_10713, wire_10712, wire_900, wire_10683, wire_10682, wire_900, wire_10759, wire_10638, wire_900, wire_11155, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11014, wire_9367, wire_904, wire_856, wire_10653, wire_10652, wire_900, wire_10743, wire_10622, wire_900, wire_10711, wire_10710, wire_860, wire_10727, wire_10726, wire_860, wire_11157, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11012, wire_9365, wire_900, wire_856, wire_10697, wire_10696, wire_860, wire_10681, wire_10680, wire_860, wire_10667, wire_10666, wire_860, wire_10757, wire_10636, wire_860, wire_11159, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_11010, wire_9363, wire_900, wire_856, wire_10651, wire_10650, wire_856, wire_10725, wire_10724, wire_856, wire_10695, wire_10694, wire_856, wire_10741, wire_10620, wire_856, wire_11131, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11038, wire_9361, wire_900, wire_856, wire_10665, wire_10664, wire_856, wire_10755, wire_10634, wire_856};
    // CHNAXY TOTAL: 621
    assign wire_9240 = lut_tile_8_1_chanxy_out[0];
    assign wire_9242 = lut_tile_8_1_chanxy_out[1];
    assign wire_9243 = lut_tile_8_1_chanxy_out[2];
    assign wire_9244 = lut_tile_8_1_chanxy_out[3];
    assign wire_9246 = lut_tile_8_1_chanxy_out[4];
    assign wire_9248 = lut_tile_8_1_chanxy_out[5];
    assign wire_9250 = lut_tile_8_1_chanxy_out[6];
    assign wire_9251 = lut_tile_8_1_chanxy_out[7];
    assign wire_9252 = lut_tile_8_1_chanxy_out[8];
    assign wire_9254 = lut_tile_8_1_chanxy_out[9];
    assign wire_9256 = lut_tile_8_1_chanxy_out[10];
    assign wire_9258 = lut_tile_8_1_chanxy_out[11];
    assign wire_9259 = lut_tile_8_1_chanxy_out[12];
    assign wire_9260 = lut_tile_8_1_chanxy_out[13];
    assign wire_9262 = lut_tile_8_1_chanxy_out[14];
    assign wire_9264 = lut_tile_8_1_chanxy_out[15];
    assign wire_9266 = lut_tile_8_1_chanxy_out[16];
    assign wire_9267 = lut_tile_8_1_chanxy_out[17];
    assign wire_9268 = lut_tile_8_1_chanxy_out[18];
    assign wire_9270 = lut_tile_8_1_chanxy_out[19];
    assign wire_9272 = lut_tile_8_1_chanxy_out[20];
    assign wire_9274 = lut_tile_8_1_chanxy_out[21];
    assign wire_9275 = lut_tile_8_1_chanxy_out[22];
    assign wire_9276 = lut_tile_8_1_chanxy_out[23];
    assign wire_9278 = lut_tile_8_1_chanxy_out[24];
    assign wire_9280 = lut_tile_8_1_chanxy_out[25];
    assign wire_9282 = lut_tile_8_1_chanxy_out[26];
    assign wire_9283 = lut_tile_8_1_chanxy_out[27];
    assign wire_9284 = lut_tile_8_1_chanxy_out[28];
    assign wire_9286 = lut_tile_8_1_chanxy_out[29];
    assign wire_9288 = lut_tile_8_1_chanxy_out[30];
    assign wire_9290 = lut_tile_8_1_chanxy_out[31];
    assign wire_9291 = lut_tile_8_1_chanxy_out[32];
    assign wire_9292 = lut_tile_8_1_chanxy_out[33];
    assign wire_9294 = lut_tile_8_1_chanxy_out[34];
    assign wire_9296 = lut_tile_8_1_chanxy_out[35];
    assign wire_9298 = lut_tile_8_1_chanxy_out[36];
    assign wire_9299 = lut_tile_8_1_chanxy_out[37];
    assign wire_9300 = lut_tile_8_1_chanxy_out[38];
    assign wire_9302 = lut_tile_8_1_chanxy_out[39];
    assign wire_9304 = lut_tile_8_1_chanxy_out[40];
    assign wire_9306 = lut_tile_8_1_chanxy_out[41];
    assign wire_9307 = lut_tile_8_1_chanxy_out[42];
    assign wire_9308 = lut_tile_8_1_chanxy_out[43];
    assign wire_9310 = lut_tile_8_1_chanxy_out[44];
    assign wire_9312 = lut_tile_8_1_chanxy_out[45];
    assign wire_9314 = lut_tile_8_1_chanxy_out[46];
    assign wire_9315 = lut_tile_8_1_chanxy_out[47];
    assign wire_9316 = lut_tile_8_1_chanxy_out[48];
    assign wire_9318 = lut_tile_8_1_chanxy_out[49];
    assign wire_9320 = lut_tile_8_1_chanxy_out[50];
    assign wire_9322 = lut_tile_8_1_chanxy_out[51];
    assign wire_9323 = lut_tile_8_1_chanxy_out[52];
    assign wire_9324 = lut_tile_8_1_chanxy_out[53];
    assign wire_9326 = lut_tile_8_1_chanxy_out[54];
    assign wire_9328 = lut_tile_8_1_chanxy_out[55];
    assign wire_9330 = lut_tile_8_1_chanxy_out[56];
    assign wire_9331 = lut_tile_8_1_chanxy_out[57];
    assign wire_9332 = lut_tile_8_1_chanxy_out[58];
    assign wire_9334 = lut_tile_8_1_chanxy_out[59];
    assign wire_9336 = lut_tile_8_1_chanxy_out[60];
    assign wire_9338 = lut_tile_8_1_chanxy_out[61];
    assign wire_9339 = lut_tile_8_1_chanxy_out[62];
    assign wire_9340 = lut_tile_8_1_chanxy_out[63];
    assign wire_9342 = lut_tile_8_1_chanxy_out[64];
    assign wire_9344 = lut_tile_8_1_chanxy_out[65];
    assign wire_9346 = lut_tile_8_1_chanxy_out[66];
    assign wire_9347 = lut_tile_8_1_chanxy_out[67];
    assign wire_9348 = lut_tile_8_1_chanxy_out[68];
    assign wire_9350 = lut_tile_8_1_chanxy_out[69];
    assign wire_9352 = lut_tile_8_1_chanxy_out[70];
    assign wire_9354 = lut_tile_8_1_chanxy_out[71];
    assign wire_9355 = lut_tile_8_1_chanxy_out[72];
    assign wire_9356 = lut_tile_8_1_chanxy_out[73];
    assign wire_9358 = lut_tile_8_1_chanxy_out[74];
    assign wire_11011 = lut_tile_8_1_chanxy_out[75];
    assign wire_11013 = lut_tile_8_1_chanxy_out[76];
    assign wire_11015 = lut_tile_8_1_chanxy_out[77];
    assign wire_11017 = lut_tile_8_1_chanxy_out[78];
    assign wire_11019 = lut_tile_8_1_chanxy_out[79];
    assign wire_11021 = lut_tile_8_1_chanxy_out[80];
    assign wire_11023 = lut_tile_8_1_chanxy_out[81];
    assign wire_11025 = lut_tile_8_1_chanxy_out[82];
    assign wire_11027 = lut_tile_8_1_chanxy_out[83];
    assign wire_11029 = lut_tile_8_1_chanxy_out[84];
    assign wire_11031 = lut_tile_8_1_chanxy_out[85];
    assign wire_11033 = lut_tile_8_1_chanxy_out[86];
    assign wire_11035 = lut_tile_8_1_chanxy_out[87];
    assign wire_11037 = lut_tile_8_1_chanxy_out[88];
    assign wire_11039 = lut_tile_8_1_chanxy_out[89];
    assign wire_11100 = lut_tile_8_1_chanxy_out[90];
    assign wire_11102 = lut_tile_8_1_chanxy_out[91];
    assign wire_11104 = lut_tile_8_1_chanxy_out[92];
    assign wire_11106 = lut_tile_8_1_chanxy_out[93];
    assign wire_11108 = lut_tile_8_1_chanxy_out[94];
    assign wire_11110 = lut_tile_8_1_chanxy_out[95];
    assign wire_11112 = lut_tile_8_1_chanxy_out[96];
    assign wire_11114 = lut_tile_8_1_chanxy_out[97];
    assign wire_11116 = lut_tile_8_1_chanxy_out[98];
    assign wire_11118 = lut_tile_8_1_chanxy_out[99];
    assign wire_11120 = lut_tile_8_1_chanxy_out[100];
    assign wire_11122 = lut_tile_8_1_chanxy_out[101];
    assign wire_11124 = lut_tile_8_1_chanxy_out[102];
    assign wire_11126 = lut_tile_8_1_chanxy_out[103];
    assign wire_11128 = lut_tile_8_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_8_2_chanxy_in = {wire_11398, wire_9001, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8860, wire_1887, wire_11396, wire_9029, wire_8967, wire_8966, wire_8927, wire_8926, wire_8887, wire_8886, wire_8868, wire_1887, wire_11394, wire_9027, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8876, wire_1887, wire_11392, wire_9025, wire_8961, wire_8960, wire_8921, wire_8920, wire_8884, wire_8881, wire_8880, wire_1377, wire_11390, wire_9023, wire_8959, wire_8958, wire_8919, wire_8918, wire_8892, wire_8879, wire_8878, wire_1377, wire_11388, wire_9021, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8900, wire_1377, wire_11386, wire_9019, wire_8953, wire_8952, wire_8913, wire_8912, wire_8908, wire_8873, wire_8872, wire_1891, wire_1377, wire_11384, wire_9017, wire_8951, wire_8950, wire_8916, wire_8911, wire_8910, wire_8871, wire_8870, wire_1891, wire_1377, wire_11382, wire_9015, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8924, wire_1891, wire_1377, wire_11380, wire_9013, wire_8945, wire_8944, wire_8932, wire_8905, wire_8904, wire_8865, wire_8864, wire_1891, wire_1373, wire_11378, wire_9011, wire_8943, wire_8942, wire_8940, wire_8903, wire_8902, wire_8863, wire_8862, wire_1891, wire_1373, wire_11376, wire_9009, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8948, wire_1891, wire_1373, wire_11374, wire_9007, wire_8956, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856, wire_1887, wire_1373, wire_11372, wire_9005, wire_8964, wire_8935, wire_8934, wire_8895, wire_8894, wire_8855, wire_8854, wire_1887, wire_1373, wire_11370, wire_9003, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8852, wire_1887, wire_1373, wire_11549, wire_9419, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_9244, wire_1887, wire_11547, wire_9391, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9356, wire_1887, wire_11545, wire_9393, wire_9353, wire_9352, wire_9348, wire_9313, wire_9312, wire_9273, wire_9272, wire_1887, wire_11543, wire_9395, wire_9351, wire_9350, wire_9340, wire_9311, wire_9310, wire_9271, wire_9270, wire_1377, wire_11541, wire_9397, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9332, wire_1377, wire_11539, wire_9399, wire_9345, wire_9344, wire_9324, wire_9305, wire_9304, wire_9265, wire_9264, wire_1377, wire_11537, wire_9401, wire_9343, wire_9342, wire_9316, wire_9303, wire_9302, wire_9263, wire_9262, wire_1891, wire_1377, wire_11535, wire_9403, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9308, wire_1891, wire_1377, wire_11533, wire_9405, wire_9337, wire_9336, wire_9300, wire_9297, wire_9296, wire_9257, wire_9256, wire_1891, wire_1377, wire_11531, wire_9407, wire_9335, wire_9334, wire_9295, wire_9294, wire_9292, wire_9255, wire_9254, wire_1891, wire_1373, wire_11529, wire_9409, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9284, wire_1891, wire_1373, wire_11527, wire_9411, wire_9329, wire_9328, wire_9289, wire_9288, wire_9276, wire_9249, wire_9248, wire_1891, wire_1373, wire_11525, wire_9413, wire_9327, wire_9326, wire_9287, wire_9286, wire_9268, wire_9247, wire_9246, wire_1887, wire_1373, wire_11523, wire_9415, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9260, wire_1887, wire_1373, wire_11521, wire_9417, wire_9321, wire_9320, wire_9281, wire_9280, wire_9252, wire_9241, wire_9240, wire_1887, wire_1373, wire_11157, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11038, wire_9354, wire_1416, wire_11155, wire_11069, wire_11068, wire_11059, wire_11058, wire_11049, wire_11048, wire_11010, wire_9346, wire_1416, wire_11153, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11012, wire_9338, wire_1416, wire_11151, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11014, wire_9330, wire_1376, wire_11149, wire_11067, wire_11066, wire_11057, wire_11056, wire_11047, wire_11046, wire_11016, wire_9322, wire_1376, wire_11147, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11018, wire_9314, wire_1376, wire_11145, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11020, wire_9306, wire_1420, wire_1376, wire_11143, wire_11065, wire_11064, wire_11055, wire_11054, wire_11045, wire_11044, wire_11022, wire_9298, wire_1420, wire_1376, wire_11141, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11024, wire_9290, wire_1420, wire_1376, wire_11139, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11026, wire_9282, wire_1420, wire_1372, wire_11137, wire_11063, wire_11062, wire_11053, wire_11052, wire_11043, wire_11042, wire_11028, wire_9274, wire_1420, wire_1372, wire_11135, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11030, wire_9266, wire_1420, wire_1372, wire_11133, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11032, wire_9258, wire_1416, wire_1372, wire_11131, wire_11061, wire_11060, wire_11051, wire_11050, wire_11041, wire_11040, wire_11034, wire_9250, wire_1416, wire_1372, wire_11159, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11036, wire_9242, wire_1416, wire_1372, wire_11523, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11426, wire_9419, wire_1416, wire_11525, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11424, wire_9417, wire_1416, wire_11527, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11422, wire_9415, wire_1416, wire_11529, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11420, wire_9413, wire_1376, wire_11531, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11418, wire_9411, wire_1376, wire_11533, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11416, wire_9409, wire_1376, wire_11535, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11414, wire_9407, wire_1420, wire_1376, wire_11537, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11412, wire_9405, wire_1420, wire_1376, wire_11539, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11410, wire_9403, wire_1420, wire_1376, wire_11541, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11408, wire_9401, wire_1420, wire_1372, wire_11543, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11406, wire_9399, wire_1420, wire_1372, wire_11545, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11404, wire_9397, wire_1420, wire_1372, wire_11547, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11402, wire_9395, wire_1416, wire_1372, wire_11549, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11400, wire_9393, wire_1416, wire_1372, wire_11521, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11428, wire_9391, wire_1416, wire_1372};
    // CHNAXY TOTAL: 636
    assign wire_9245 = lut_tile_8_2_chanxy_out[0];
    assign wire_9253 = lut_tile_8_2_chanxy_out[1];
    assign wire_9261 = lut_tile_8_2_chanxy_out[2];
    assign wire_9269 = lut_tile_8_2_chanxy_out[3];
    assign wire_9277 = lut_tile_8_2_chanxy_out[4];
    assign wire_9285 = lut_tile_8_2_chanxy_out[5];
    assign wire_9293 = lut_tile_8_2_chanxy_out[6];
    assign wire_9301 = lut_tile_8_2_chanxy_out[7];
    assign wire_9309 = lut_tile_8_2_chanxy_out[8];
    assign wire_9317 = lut_tile_8_2_chanxy_out[9];
    assign wire_9325 = lut_tile_8_2_chanxy_out[10];
    assign wire_9333 = lut_tile_8_2_chanxy_out[11];
    assign wire_9341 = lut_tile_8_2_chanxy_out[12];
    assign wire_9349 = lut_tile_8_2_chanxy_out[13];
    assign wire_9357 = lut_tile_8_2_chanxy_out[14];
    assign wire_9360 = lut_tile_8_2_chanxy_out[15];
    assign wire_9362 = lut_tile_8_2_chanxy_out[16];
    assign wire_9364 = lut_tile_8_2_chanxy_out[17];
    assign wire_9366 = lut_tile_8_2_chanxy_out[18];
    assign wire_9368 = lut_tile_8_2_chanxy_out[19];
    assign wire_9370 = lut_tile_8_2_chanxy_out[20];
    assign wire_9372 = lut_tile_8_2_chanxy_out[21];
    assign wire_9374 = lut_tile_8_2_chanxy_out[22];
    assign wire_9376 = lut_tile_8_2_chanxy_out[23];
    assign wire_9378 = lut_tile_8_2_chanxy_out[24];
    assign wire_9380 = lut_tile_8_2_chanxy_out[25];
    assign wire_9382 = lut_tile_8_2_chanxy_out[26];
    assign wire_9384 = lut_tile_8_2_chanxy_out[27];
    assign wire_9386 = lut_tile_8_2_chanxy_out[28];
    assign wire_9388 = lut_tile_8_2_chanxy_out[29];
    assign wire_11401 = lut_tile_8_2_chanxy_out[30];
    assign wire_11403 = lut_tile_8_2_chanxy_out[31];
    assign wire_11405 = lut_tile_8_2_chanxy_out[32];
    assign wire_11407 = lut_tile_8_2_chanxy_out[33];
    assign wire_11409 = lut_tile_8_2_chanxy_out[34];
    assign wire_11411 = lut_tile_8_2_chanxy_out[35];
    assign wire_11413 = lut_tile_8_2_chanxy_out[36];
    assign wire_11415 = lut_tile_8_2_chanxy_out[37];
    assign wire_11417 = lut_tile_8_2_chanxy_out[38];
    assign wire_11419 = lut_tile_8_2_chanxy_out[39];
    assign wire_11421 = lut_tile_8_2_chanxy_out[40];
    assign wire_11423 = lut_tile_8_2_chanxy_out[41];
    assign wire_11425 = lut_tile_8_2_chanxy_out[42];
    assign wire_11427 = lut_tile_8_2_chanxy_out[43];
    assign wire_11429 = lut_tile_8_2_chanxy_out[44];
    assign wire_11490 = lut_tile_8_2_chanxy_out[45];
    assign wire_11492 = lut_tile_8_2_chanxy_out[46];
    assign wire_11494 = lut_tile_8_2_chanxy_out[47];
    assign wire_11496 = lut_tile_8_2_chanxy_out[48];
    assign wire_11498 = lut_tile_8_2_chanxy_out[49];
    assign wire_11500 = lut_tile_8_2_chanxy_out[50];
    assign wire_11502 = lut_tile_8_2_chanxy_out[51];
    assign wire_11504 = lut_tile_8_2_chanxy_out[52];
    assign wire_11506 = lut_tile_8_2_chanxy_out[53];
    assign wire_11508 = lut_tile_8_2_chanxy_out[54];
    assign wire_11510 = lut_tile_8_2_chanxy_out[55];
    assign wire_11512 = lut_tile_8_2_chanxy_out[56];
    assign wire_11514 = lut_tile_8_2_chanxy_out[57];
    assign wire_11516 = lut_tile_8_2_chanxy_out[58];
    assign wire_11518 = lut_tile_8_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_3_chanxy_in = {wire_11788, wire_9031, wire_8969, wire_8968, wire_8929, wire_8928, wire_8889, wire_8888, wire_8862, wire_2403, wire_11786, wire_9059, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8870, wire_2403, wire_11784, wire_9057, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8878, wire_2403, wire_11782, wire_9055, wire_8961, wire_8960, wire_8921, wire_8920, wire_8886, wire_8881, wire_8880, wire_1893, wire_11780, wire_9053, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8894, wire_1893, wire_11778, wire_9051, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8902, wire_1893, wire_11776, wire_9049, wire_8953, wire_8952, wire_8913, wire_8912, wire_8910, wire_8873, wire_8872, wire_2407, wire_1893, wire_11774, wire_9047, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8918, wire_2407, wire_1893, wire_11772, wire_9045, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8926, wire_2407, wire_1893, wire_11770, wire_9043, wire_8945, wire_8944, wire_8934, wire_8905, wire_8904, wire_8865, wire_8864, wire_2407, wire_1889, wire_11768, wire_9041, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8942, wire_2407, wire_1889, wire_11766, wire_9039, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8950, wire_2407, wire_1889, wire_11764, wire_9037, wire_8958, wire_8937, wire_8936, wire_8897, wire_8896, wire_8857, wire_8856, wire_2403, wire_1889, wire_11762, wire_9035, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8966, wire_2403, wire_1889, wire_11760, wire_9033, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8854, wire_2403, wire_1889, wire_11939, wire_9449, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9246, wire_2403, wire_11937, wire_9421, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9358, wire_2403, wire_11935, wire_9423, wire_9353, wire_9352, wire_9350, wire_9313, wire_9312, wire_9273, wire_9272, wire_2403, wire_11933, wire_9425, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9342, wire_1893, wire_11931, wire_9427, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9334, wire_1893, wire_11929, wire_9429, wire_9345, wire_9344, wire_9326, wire_9305, wire_9304, wire_9265, wire_9264, wire_1893, wire_11927, wire_9431, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9318, wire_2407, wire_1893, wire_11925, wire_9433, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9310, wire_2407, wire_1893, wire_11923, wire_9435, wire_9337, wire_9336, wire_9302, wire_9297, wire_9296, wire_9257, wire_9256, wire_2407, wire_1893, wire_11921, wire_9437, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9294, wire_2407, wire_1889, wire_11919, wire_9439, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9286, wire_2407, wire_1889, wire_11917, wire_9441, wire_9329, wire_9328, wire_9289, wire_9288, wire_9278, wire_9249, wire_9248, wire_2407, wire_1889, wire_11915, wire_9443, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9270, wire_2403, wire_1889, wire_11913, wire_9445, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9262, wire_2403, wire_1889, wire_11911, wire_9447, wire_9321, wire_9320, wire_9281, wire_9280, wire_9254, wire_9241, wire_9240, wire_2403, wire_1889, wire_11547, wire_11459, wire_11458, wire_11449, wire_11448, wire_11439, wire_11438, wire_11428, wire_9356, wire_1932, wire_11545, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11400, wire_9348, wire_1932, wire_11543, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11402, wire_9340, wire_1932, wire_11541, wire_11457, wire_11456, wire_11447, wire_11446, wire_11437, wire_11436, wire_11404, wire_9332, wire_1892, wire_11539, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11406, wire_9324, wire_1892, wire_11537, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11408, wire_9316, wire_1892, wire_11535, wire_11455, wire_11454, wire_11445, wire_11444, wire_11435, wire_11434, wire_11410, wire_9308, wire_1936, wire_1892, wire_11533, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11412, wire_9300, wire_1936, wire_1892, wire_11531, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11414, wire_9292, wire_1936, wire_1892, wire_11529, wire_11453, wire_11452, wire_11443, wire_11442, wire_11433, wire_11432, wire_11416, wire_9284, wire_1936, wire_1888, wire_11527, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11418, wire_9276, wire_1936, wire_1888, wire_11525, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11420, wire_9268, wire_1936, wire_1888, wire_11523, wire_11451, wire_11450, wire_11441, wire_11440, wire_11431, wire_11430, wire_11422, wire_9260, wire_1932, wire_1888, wire_11521, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11424, wire_9252, wire_1932, wire_1888, wire_11549, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11426, wire_9244, wire_1932, wire_1888, wire_11913, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11816, wire_9449, wire_1932, wire_11915, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11814, wire_9447, wire_1932, wire_11917, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11812, wire_9445, wire_1932, wire_11919, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11810, wire_9443, wire_1892, wire_11921, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11808, wire_9441, wire_1892, wire_11923, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11806, wire_9439, wire_1892, wire_11925, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11804, wire_9437, wire_1936, wire_1892, wire_11927, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11802, wire_9435, wire_1936, wire_1892, wire_11929, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11800, wire_9433, wire_1936, wire_1892, wire_11931, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11798, wire_9431, wire_1936, wire_1888, wire_11933, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11796, wire_9429, wire_1936, wire_1888, wire_11935, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11794, wire_9427, wire_1936, wire_1888, wire_11937, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11792, wire_9425, wire_1932, wire_1888, wire_11939, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11790, wire_9423, wire_1932, wire_1888, wire_11911, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11818, wire_9421, wire_1932, wire_1888};
    // CHNAXY TOTAL: 636
    assign wire_9247 = lut_tile_8_3_chanxy_out[0];
    assign wire_9255 = lut_tile_8_3_chanxy_out[1];
    assign wire_9263 = lut_tile_8_3_chanxy_out[2];
    assign wire_9271 = lut_tile_8_3_chanxy_out[3];
    assign wire_9279 = lut_tile_8_3_chanxy_out[4];
    assign wire_9287 = lut_tile_8_3_chanxy_out[5];
    assign wire_9295 = lut_tile_8_3_chanxy_out[6];
    assign wire_9303 = lut_tile_8_3_chanxy_out[7];
    assign wire_9311 = lut_tile_8_3_chanxy_out[8];
    assign wire_9319 = lut_tile_8_3_chanxy_out[9];
    assign wire_9327 = lut_tile_8_3_chanxy_out[10];
    assign wire_9335 = lut_tile_8_3_chanxy_out[11];
    assign wire_9343 = lut_tile_8_3_chanxy_out[12];
    assign wire_9351 = lut_tile_8_3_chanxy_out[13];
    assign wire_9359 = lut_tile_8_3_chanxy_out[14];
    assign wire_9390 = lut_tile_8_3_chanxy_out[15];
    assign wire_9392 = lut_tile_8_3_chanxy_out[16];
    assign wire_9394 = lut_tile_8_3_chanxy_out[17];
    assign wire_9396 = lut_tile_8_3_chanxy_out[18];
    assign wire_9398 = lut_tile_8_3_chanxy_out[19];
    assign wire_9400 = lut_tile_8_3_chanxy_out[20];
    assign wire_9402 = lut_tile_8_3_chanxy_out[21];
    assign wire_9404 = lut_tile_8_3_chanxy_out[22];
    assign wire_9406 = lut_tile_8_3_chanxy_out[23];
    assign wire_9408 = lut_tile_8_3_chanxy_out[24];
    assign wire_9410 = lut_tile_8_3_chanxy_out[25];
    assign wire_9412 = lut_tile_8_3_chanxy_out[26];
    assign wire_9414 = lut_tile_8_3_chanxy_out[27];
    assign wire_9416 = lut_tile_8_3_chanxy_out[28];
    assign wire_9418 = lut_tile_8_3_chanxy_out[29];
    assign wire_11791 = lut_tile_8_3_chanxy_out[30];
    assign wire_11793 = lut_tile_8_3_chanxy_out[31];
    assign wire_11795 = lut_tile_8_3_chanxy_out[32];
    assign wire_11797 = lut_tile_8_3_chanxy_out[33];
    assign wire_11799 = lut_tile_8_3_chanxy_out[34];
    assign wire_11801 = lut_tile_8_3_chanxy_out[35];
    assign wire_11803 = lut_tile_8_3_chanxy_out[36];
    assign wire_11805 = lut_tile_8_3_chanxy_out[37];
    assign wire_11807 = lut_tile_8_3_chanxy_out[38];
    assign wire_11809 = lut_tile_8_3_chanxy_out[39];
    assign wire_11811 = lut_tile_8_3_chanxy_out[40];
    assign wire_11813 = lut_tile_8_3_chanxy_out[41];
    assign wire_11815 = lut_tile_8_3_chanxy_out[42];
    assign wire_11817 = lut_tile_8_3_chanxy_out[43];
    assign wire_11819 = lut_tile_8_3_chanxy_out[44];
    assign wire_11880 = lut_tile_8_3_chanxy_out[45];
    assign wire_11882 = lut_tile_8_3_chanxy_out[46];
    assign wire_11884 = lut_tile_8_3_chanxy_out[47];
    assign wire_11886 = lut_tile_8_3_chanxy_out[48];
    assign wire_11888 = lut_tile_8_3_chanxy_out[49];
    assign wire_11890 = lut_tile_8_3_chanxy_out[50];
    assign wire_11892 = lut_tile_8_3_chanxy_out[51];
    assign wire_11894 = lut_tile_8_3_chanxy_out[52];
    assign wire_11896 = lut_tile_8_3_chanxy_out[53];
    assign wire_11898 = lut_tile_8_3_chanxy_out[54];
    assign wire_11900 = lut_tile_8_3_chanxy_out[55];
    assign wire_11902 = lut_tile_8_3_chanxy_out[56];
    assign wire_11904 = lut_tile_8_3_chanxy_out[57];
    assign wire_11906 = lut_tile_8_3_chanxy_out[58];
    assign wire_11908 = lut_tile_8_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_4_chanxy_in = {wire_12178, wire_9061, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8864, wire_2919, wire_12176, wire_9089, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8872, wire_2919, wire_12174, wire_9087, wire_8999, wire_8998, wire_8989, wire_8988, wire_8979, wire_8978, wire_8880, wire_2919, wire_12172, wire_9085, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8888, wire_2409, wire_12170, wire_9083, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8896, wire_2409, wire_12168, wire_9081, wire_8997, wire_8996, wire_8987, wire_8986, wire_8977, wire_8976, wire_8904, wire_2409, wire_12166, wire_9079, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8912, wire_2923, wire_2409, wire_12164, wire_9077, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8920, wire_2923, wire_2409, wire_12162, wire_9075, wire_8995, wire_8994, wire_8985, wire_8984, wire_8975, wire_8974, wire_8928, wire_2923, wire_2409, wire_12160, wire_9073, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8936, wire_2923, wire_2405, wire_12158, wire_9071, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8944, wire_2923, wire_2405, wire_12156, wire_9069, wire_8993, wire_8992, wire_8983, wire_8982, wire_8973, wire_8972, wire_8952, wire_2923, wire_2405, wire_12154, wire_9067, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8960, wire_2919, wire_2405, wire_12152, wire_9065, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8968, wire_2919, wire_2405, wire_12150, wire_9063, wire_8991, wire_8990, wire_8981, wire_8980, wire_8971, wire_8970, wire_8856, wire_2919, wire_2405, wire_12329, wire_9479, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9240, wire_2919, wire_12327, wire_9451, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9352, wire_2919, wire_12325, wire_9453, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9344, wire_2919, wire_12323, wire_9455, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9336, wire_2409, wire_12321, wire_9457, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9328, wire_2409, wire_12319, wire_9459, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9320, wire_2409, wire_12317, wire_9461, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9312, wire_2923, wire_2409, wire_12315, wire_9463, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9304, wire_2923, wire_2409, wire_12313, wire_9465, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9296, wire_2923, wire_2409, wire_12311, wire_9467, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9288, wire_2923, wire_2405, wire_12309, wire_9469, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9280, wire_2923, wire_2405, wire_12307, wire_9471, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9272, wire_2923, wire_2405, wire_12305, wire_9473, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9264, wire_2919, wire_2405, wire_12303, wire_9475, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9256, wire_2919, wire_2405, wire_12301, wire_9477, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9248, wire_2919, wire_2405, wire_11937, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11818, wire_9358, wire_2448, wire_11935, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11790, wire_9350, wire_2448, wire_11933, wire_11849, wire_11848, wire_11839, wire_11838, wire_11829, wire_11828, wire_11792, wire_9342, wire_2448, wire_11931, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11794, wire_9334, wire_2408, wire_11929, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11796, wire_9326, wire_2408, wire_11927, wire_11847, wire_11846, wire_11837, wire_11836, wire_11827, wire_11826, wire_11798, wire_9318, wire_2408, wire_11925, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11800, wire_9310, wire_2452, wire_2408, wire_11923, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11802, wire_9302, wire_2452, wire_2408, wire_11921, wire_11845, wire_11844, wire_11835, wire_11834, wire_11825, wire_11824, wire_11804, wire_9294, wire_2452, wire_2408, wire_11919, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11806, wire_9286, wire_2452, wire_2404, wire_11917, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11808, wire_9278, wire_2452, wire_2404, wire_11915, wire_11843, wire_11842, wire_11833, wire_11832, wire_11823, wire_11822, wire_11810, wire_9270, wire_2452, wire_2404, wire_11913, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11812, wire_9262, wire_2448, wire_2404, wire_11911, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11814, wire_9254, wire_2448, wire_2404, wire_11939, wire_11841, wire_11840, wire_11831, wire_11830, wire_11821, wire_11820, wire_11816, wire_9246, wire_2448, wire_2404, wire_12303, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12206, wire_9479, wire_2448, wire_12305, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12204, wire_9477, wire_2448, wire_12307, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12202, wire_9475, wire_2448, wire_12309, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12200, wire_9473, wire_2408, wire_12311, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12198, wire_9471, wire_2408, wire_12313, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12196, wire_9469, wire_2408, wire_12315, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12194, wire_9467, wire_2452, wire_2408, wire_12317, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12192, wire_9465, wire_2452, wire_2408, wire_12319, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12190, wire_9463, wire_2452, wire_2408, wire_12321, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12188, wire_9461, wire_2452, wire_2404, wire_12323, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12186, wire_9459, wire_2452, wire_2404, wire_12325, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12184, wire_9457, wire_2452, wire_2404, wire_12327, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12182, wire_9455, wire_2448, wire_2404, wire_12329, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12180, wire_9453, wire_2448, wire_2404, wire_12301, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12208, wire_9451, wire_2448, wire_2404};
    // CHNAXY TOTAL: 636
    assign wire_9241 = lut_tile_8_4_chanxy_out[0];
    assign wire_9249 = lut_tile_8_4_chanxy_out[1];
    assign wire_9257 = lut_tile_8_4_chanxy_out[2];
    assign wire_9265 = lut_tile_8_4_chanxy_out[3];
    assign wire_9273 = lut_tile_8_4_chanxy_out[4];
    assign wire_9281 = lut_tile_8_4_chanxy_out[5];
    assign wire_9289 = lut_tile_8_4_chanxy_out[6];
    assign wire_9297 = lut_tile_8_4_chanxy_out[7];
    assign wire_9305 = lut_tile_8_4_chanxy_out[8];
    assign wire_9313 = lut_tile_8_4_chanxy_out[9];
    assign wire_9321 = lut_tile_8_4_chanxy_out[10];
    assign wire_9329 = lut_tile_8_4_chanxy_out[11];
    assign wire_9337 = lut_tile_8_4_chanxy_out[12];
    assign wire_9345 = lut_tile_8_4_chanxy_out[13];
    assign wire_9353 = lut_tile_8_4_chanxy_out[14];
    assign wire_9420 = lut_tile_8_4_chanxy_out[15];
    assign wire_9422 = lut_tile_8_4_chanxy_out[16];
    assign wire_9424 = lut_tile_8_4_chanxy_out[17];
    assign wire_9426 = lut_tile_8_4_chanxy_out[18];
    assign wire_9428 = lut_tile_8_4_chanxy_out[19];
    assign wire_9430 = lut_tile_8_4_chanxy_out[20];
    assign wire_9432 = lut_tile_8_4_chanxy_out[21];
    assign wire_9434 = lut_tile_8_4_chanxy_out[22];
    assign wire_9436 = lut_tile_8_4_chanxy_out[23];
    assign wire_9438 = lut_tile_8_4_chanxy_out[24];
    assign wire_9440 = lut_tile_8_4_chanxy_out[25];
    assign wire_9442 = lut_tile_8_4_chanxy_out[26];
    assign wire_9444 = lut_tile_8_4_chanxy_out[27];
    assign wire_9446 = lut_tile_8_4_chanxy_out[28];
    assign wire_9448 = lut_tile_8_4_chanxy_out[29];
    assign wire_12181 = lut_tile_8_4_chanxy_out[30];
    assign wire_12183 = lut_tile_8_4_chanxy_out[31];
    assign wire_12185 = lut_tile_8_4_chanxy_out[32];
    assign wire_12187 = lut_tile_8_4_chanxy_out[33];
    assign wire_12189 = lut_tile_8_4_chanxy_out[34];
    assign wire_12191 = lut_tile_8_4_chanxy_out[35];
    assign wire_12193 = lut_tile_8_4_chanxy_out[36];
    assign wire_12195 = lut_tile_8_4_chanxy_out[37];
    assign wire_12197 = lut_tile_8_4_chanxy_out[38];
    assign wire_12199 = lut_tile_8_4_chanxy_out[39];
    assign wire_12201 = lut_tile_8_4_chanxy_out[40];
    assign wire_12203 = lut_tile_8_4_chanxy_out[41];
    assign wire_12205 = lut_tile_8_4_chanxy_out[42];
    assign wire_12207 = lut_tile_8_4_chanxy_out[43];
    assign wire_12209 = lut_tile_8_4_chanxy_out[44];
    assign wire_12270 = lut_tile_8_4_chanxy_out[45];
    assign wire_12272 = lut_tile_8_4_chanxy_out[46];
    assign wire_12274 = lut_tile_8_4_chanxy_out[47];
    assign wire_12276 = lut_tile_8_4_chanxy_out[48];
    assign wire_12278 = lut_tile_8_4_chanxy_out[49];
    assign wire_12280 = lut_tile_8_4_chanxy_out[50];
    assign wire_12282 = lut_tile_8_4_chanxy_out[51];
    assign wire_12284 = lut_tile_8_4_chanxy_out[52];
    assign wire_12286 = lut_tile_8_4_chanxy_out[53];
    assign wire_12288 = lut_tile_8_4_chanxy_out[54];
    assign wire_12290 = lut_tile_8_4_chanxy_out[55];
    assign wire_12292 = lut_tile_8_4_chanxy_out[56];
    assign wire_12294 = lut_tile_8_4_chanxy_out[57];
    assign wire_12296 = lut_tile_8_4_chanxy_out[58];
    assign wire_12298 = lut_tile_8_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_5_chanxy_in = {wire_12568, wire_9091, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_8972, wire_3435, wire_12566, wire_9119, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_8974, wire_3435, wire_12564, wire_9117, wire_9029, wire_9028, wire_9019, wire_9018, wire_9009, wire_9008, wire_8976, wire_3435, wire_12562, wire_9115, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_8978, wire_2925, wire_12560, wire_9113, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_8980, wire_2925, wire_12558, wire_9111, wire_9027, wire_9026, wire_9017, wire_9016, wire_9007, wire_9006, wire_8982, wire_2925, wire_12556, wire_9109, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_8984, wire_3439, wire_2925, wire_12554, wire_9107, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_8986, wire_3439, wire_2925, wire_12552, wire_9105, wire_9025, wire_9024, wire_9015, wire_9014, wire_9005, wire_9004, wire_8988, wire_3439, wire_2925, wire_12550, wire_9103, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_8990, wire_3439, wire_2921, wire_12548, wire_9101, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_8992, wire_3439, wire_2921, wire_12546, wire_9099, wire_9023, wire_9022, wire_9013, wire_9012, wire_9003, wire_9002, wire_8994, wire_3439, wire_2921, wire_12544, wire_9097, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_8996, wire_3435, wire_2921, wire_12542, wire_9095, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_8998, wire_3435, wire_2921, wire_12540, wire_9093, wire_9021, wire_9020, wire_9011, wire_9010, wire_9001, wire_9000, wire_8970, wire_3435, wire_2921, wire_12719, wire_9509, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9360, wire_3435, wire_12717, wire_9481, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9388, wire_3435, wire_12715, wire_9483, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9386, wire_3435, wire_12713, wire_9485, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9384, wire_2925, wire_12711, wire_9487, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9382, wire_2925, wire_12709, wire_9489, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9380, wire_2925, wire_12707, wire_9491, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9378, wire_3439, wire_2925, wire_12705, wire_9493, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9376, wire_3439, wire_2925, wire_12703, wire_9495, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9374, wire_3439, wire_2925, wire_12701, wire_9497, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9372, wire_3439, wire_2921, wire_12699, wire_9499, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9370, wire_3439, wire_2921, wire_12697, wire_9501, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9368, wire_3439, wire_2921, wire_12695, wire_9503, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9366, wire_3435, wire_2921, wire_12693, wire_9505, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9364, wire_3435, wire_2921, wire_12691, wire_9507, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9362, wire_3435, wire_2921, wire_12327, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12208, wire_9352, wire_2964, wire_12325, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12180, wire_9344, wire_2964, wire_12323, wire_12239, wire_12238, wire_12229, wire_12228, wire_12219, wire_12218, wire_12182, wire_9336, wire_2964, wire_12321, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12184, wire_9328, wire_2924, wire_12319, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12186, wire_9320, wire_2924, wire_12317, wire_12237, wire_12236, wire_12227, wire_12226, wire_12217, wire_12216, wire_12188, wire_9312, wire_2924, wire_12315, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12190, wire_9304, wire_2968, wire_2924, wire_12313, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12192, wire_9296, wire_2968, wire_2924, wire_12311, wire_12235, wire_12234, wire_12225, wire_12224, wire_12215, wire_12214, wire_12194, wire_9288, wire_2968, wire_2924, wire_12309, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12196, wire_9280, wire_2968, wire_2920, wire_12307, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12198, wire_9272, wire_2968, wire_2920, wire_12305, wire_12233, wire_12232, wire_12223, wire_12222, wire_12213, wire_12212, wire_12200, wire_9264, wire_2968, wire_2920, wire_12303, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12202, wire_9256, wire_2964, wire_2920, wire_12301, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12204, wire_9248, wire_2964, wire_2920, wire_12329, wire_12231, wire_12230, wire_12221, wire_12220, wire_12211, wire_12210, wire_12206, wire_9240, wire_2964, wire_2920, wire_12693, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12596, wire_9509, wire_2964, wire_12695, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12594, wire_9507, wire_2964, wire_12697, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12592, wire_9505, wire_2964, wire_12699, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12590, wire_9503, wire_2924, wire_12701, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12588, wire_9501, wire_2924, wire_12703, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12586, wire_9499, wire_2924, wire_12705, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12584, wire_9497, wire_2968, wire_2924, wire_12707, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12582, wire_9495, wire_2968, wire_2924, wire_12709, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12580, wire_9493, wire_2968, wire_2924, wire_12711, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12578, wire_9491, wire_2968, wire_2920, wire_12713, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12576, wire_9489, wire_2968, wire_2920, wire_12715, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12574, wire_9487, wire_2968, wire_2920, wire_12717, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12572, wire_9485, wire_2964, wire_2920, wire_12719, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12570, wire_9483, wire_2964, wire_2920, wire_12691, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12598, wire_9481, wire_2964, wire_2920};
    // CHNAXY TOTAL: 636
    assign wire_9361 = lut_tile_8_5_chanxy_out[0];
    assign wire_9363 = lut_tile_8_5_chanxy_out[1];
    assign wire_9365 = lut_tile_8_5_chanxy_out[2];
    assign wire_9367 = lut_tile_8_5_chanxy_out[3];
    assign wire_9369 = lut_tile_8_5_chanxy_out[4];
    assign wire_9371 = lut_tile_8_5_chanxy_out[5];
    assign wire_9373 = lut_tile_8_5_chanxy_out[6];
    assign wire_9375 = lut_tile_8_5_chanxy_out[7];
    assign wire_9377 = lut_tile_8_5_chanxy_out[8];
    assign wire_9379 = lut_tile_8_5_chanxy_out[9];
    assign wire_9381 = lut_tile_8_5_chanxy_out[10];
    assign wire_9383 = lut_tile_8_5_chanxy_out[11];
    assign wire_9385 = lut_tile_8_5_chanxy_out[12];
    assign wire_9387 = lut_tile_8_5_chanxy_out[13];
    assign wire_9389 = lut_tile_8_5_chanxy_out[14];
    assign wire_9450 = lut_tile_8_5_chanxy_out[15];
    assign wire_9452 = lut_tile_8_5_chanxy_out[16];
    assign wire_9454 = lut_tile_8_5_chanxy_out[17];
    assign wire_9456 = lut_tile_8_5_chanxy_out[18];
    assign wire_9458 = lut_tile_8_5_chanxy_out[19];
    assign wire_9460 = lut_tile_8_5_chanxy_out[20];
    assign wire_9462 = lut_tile_8_5_chanxy_out[21];
    assign wire_9464 = lut_tile_8_5_chanxy_out[22];
    assign wire_9466 = lut_tile_8_5_chanxy_out[23];
    assign wire_9468 = lut_tile_8_5_chanxy_out[24];
    assign wire_9470 = lut_tile_8_5_chanxy_out[25];
    assign wire_9472 = lut_tile_8_5_chanxy_out[26];
    assign wire_9474 = lut_tile_8_5_chanxy_out[27];
    assign wire_9476 = lut_tile_8_5_chanxy_out[28];
    assign wire_9478 = lut_tile_8_5_chanxy_out[29];
    assign wire_12571 = lut_tile_8_5_chanxy_out[30];
    assign wire_12573 = lut_tile_8_5_chanxy_out[31];
    assign wire_12575 = lut_tile_8_5_chanxy_out[32];
    assign wire_12577 = lut_tile_8_5_chanxy_out[33];
    assign wire_12579 = lut_tile_8_5_chanxy_out[34];
    assign wire_12581 = lut_tile_8_5_chanxy_out[35];
    assign wire_12583 = lut_tile_8_5_chanxy_out[36];
    assign wire_12585 = lut_tile_8_5_chanxy_out[37];
    assign wire_12587 = lut_tile_8_5_chanxy_out[38];
    assign wire_12589 = lut_tile_8_5_chanxy_out[39];
    assign wire_12591 = lut_tile_8_5_chanxy_out[40];
    assign wire_12593 = lut_tile_8_5_chanxy_out[41];
    assign wire_12595 = lut_tile_8_5_chanxy_out[42];
    assign wire_12597 = lut_tile_8_5_chanxy_out[43];
    assign wire_12599 = lut_tile_8_5_chanxy_out[44];
    assign wire_12660 = lut_tile_8_5_chanxy_out[45];
    assign wire_12662 = lut_tile_8_5_chanxy_out[46];
    assign wire_12664 = lut_tile_8_5_chanxy_out[47];
    assign wire_12666 = lut_tile_8_5_chanxy_out[48];
    assign wire_12668 = lut_tile_8_5_chanxy_out[49];
    assign wire_12670 = lut_tile_8_5_chanxy_out[50];
    assign wire_12672 = lut_tile_8_5_chanxy_out[51];
    assign wire_12674 = lut_tile_8_5_chanxy_out[52];
    assign wire_12676 = lut_tile_8_5_chanxy_out[53];
    assign wire_12678 = lut_tile_8_5_chanxy_out[54];
    assign wire_12680 = lut_tile_8_5_chanxy_out[55];
    assign wire_12682 = lut_tile_8_5_chanxy_out[56];
    assign wire_12684 = lut_tile_8_5_chanxy_out[57];
    assign wire_12686 = lut_tile_8_5_chanxy_out[58];
    assign wire_12688 = lut_tile_8_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_6_chanxy_in = {wire_12958, wire_9121, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9002, wire_3951, wire_12956, wire_9149, wire_9059, wire_9058, wire_9049, wire_9048, wire_9039, wire_9038, wire_9004, wire_3951, wire_12954, wire_9147, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9006, wire_3951, wire_12952, wire_9145, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9008, wire_3441, wire_12950, wire_9143, wire_9057, wire_9056, wire_9047, wire_9046, wire_9037, wire_9036, wire_9010, wire_3441, wire_12948, wire_9141, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9012, wire_3441, wire_12946, wire_9139, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9014, wire_3955, wire_3441, wire_12944, wire_9137, wire_9055, wire_9054, wire_9045, wire_9044, wire_9035, wire_9034, wire_9016, wire_3955, wire_3441, wire_12942, wire_9135, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9018, wire_3955, wire_3441, wire_12940, wire_9133, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9020, wire_3955, wire_3437, wire_12938, wire_9131, wire_9053, wire_9052, wire_9043, wire_9042, wire_9033, wire_9032, wire_9022, wire_3955, wire_3437, wire_12936, wire_9129, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9024, wire_3955, wire_3437, wire_12934, wire_9127, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9026, wire_3951, wire_3437, wire_12932, wire_9125, wire_9051, wire_9050, wire_9041, wire_9040, wire_9031, wire_9030, wire_9028, wire_3951, wire_3437, wire_12930, wire_9123, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9000, wire_3951, wire_3437, wire_13109, wire_9539, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9390, wire_3951, wire_13107, wire_9511, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9418, wire_3951, wire_13105, wire_9513, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9416, wire_3951, wire_13103, wire_9515, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9414, wire_3441, wire_13101, wire_9517, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9412, wire_3441, wire_13099, wire_9519, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9410, wire_3441, wire_13097, wire_9521, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9408, wire_3955, wire_3441, wire_13095, wire_9523, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9406, wire_3955, wire_3441, wire_13093, wire_9525, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9404, wire_3955, wire_3441, wire_13091, wire_9527, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9402, wire_3955, wire_3437, wire_13089, wire_9529, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9400, wire_3955, wire_3437, wire_13087, wire_9531, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9398, wire_3955, wire_3437, wire_13085, wire_9533, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9396, wire_3951, wire_3437, wire_13083, wire_9535, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9394, wire_3951, wire_3437, wire_13081, wire_9537, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9392, wire_3951, wire_3437, wire_12717, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12598, wire_9388, wire_3480, wire_12715, wire_12629, wire_12628, wire_12619, wire_12618, wire_12609, wire_12608, wire_12570, wire_9386, wire_3480, wire_12713, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12572, wire_9384, wire_3480, wire_12711, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12574, wire_9382, wire_3440, wire_12709, wire_12627, wire_12626, wire_12617, wire_12616, wire_12607, wire_12606, wire_12576, wire_9380, wire_3440, wire_12707, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12578, wire_9378, wire_3440, wire_12705, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12580, wire_9376, wire_3484, wire_3440, wire_12703, wire_12625, wire_12624, wire_12615, wire_12614, wire_12605, wire_12604, wire_12582, wire_9374, wire_3484, wire_3440, wire_12701, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12584, wire_9372, wire_3484, wire_3440, wire_12699, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12586, wire_9370, wire_3484, wire_3436, wire_12697, wire_12623, wire_12622, wire_12613, wire_12612, wire_12603, wire_12602, wire_12588, wire_9368, wire_3484, wire_3436, wire_12695, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12590, wire_9366, wire_3484, wire_3436, wire_12693, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12592, wire_9364, wire_3480, wire_3436, wire_12691, wire_12621, wire_12620, wire_12611, wire_12610, wire_12601, wire_12600, wire_12594, wire_9362, wire_3480, wire_3436, wire_12719, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12596, wire_9360, wire_3480, wire_3436, wire_13083, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12986, wire_9539, wire_3480, wire_13085, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_12984, wire_9537, wire_3480, wire_13087, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12982, wire_9535, wire_3480, wire_13089, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12980, wire_9533, wire_3440, wire_13091, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_12978, wire_9531, wire_3440, wire_13093, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12976, wire_9529, wire_3440, wire_13095, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12974, wire_9527, wire_3484, wire_3440, wire_13097, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_12972, wire_9525, wire_3484, wire_3440, wire_13099, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12970, wire_9523, wire_3484, wire_3440, wire_13101, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12968, wire_9521, wire_3484, wire_3436, wire_13103, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_12966, wire_9519, wire_3484, wire_3436, wire_13105, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12964, wire_9517, wire_3484, wire_3436, wire_13107, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12962, wire_9515, wire_3480, wire_3436, wire_13109, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_12960, wire_9513, wire_3480, wire_3436, wire_13081, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12988, wire_9511, wire_3480, wire_3436};
    // CHNAXY TOTAL: 636
    assign wire_9391 = lut_tile_8_6_chanxy_out[0];
    assign wire_9393 = lut_tile_8_6_chanxy_out[1];
    assign wire_9395 = lut_tile_8_6_chanxy_out[2];
    assign wire_9397 = lut_tile_8_6_chanxy_out[3];
    assign wire_9399 = lut_tile_8_6_chanxy_out[4];
    assign wire_9401 = lut_tile_8_6_chanxy_out[5];
    assign wire_9403 = lut_tile_8_6_chanxy_out[6];
    assign wire_9405 = lut_tile_8_6_chanxy_out[7];
    assign wire_9407 = lut_tile_8_6_chanxy_out[8];
    assign wire_9409 = lut_tile_8_6_chanxy_out[9];
    assign wire_9411 = lut_tile_8_6_chanxy_out[10];
    assign wire_9413 = lut_tile_8_6_chanxy_out[11];
    assign wire_9415 = lut_tile_8_6_chanxy_out[12];
    assign wire_9417 = lut_tile_8_6_chanxy_out[13];
    assign wire_9419 = lut_tile_8_6_chanxy_out[14];
    assign wire_9480 = lut_tile_8_6_chanxy_out[15];
    assign wire_9482 = lut_tile_8_6_chanxy_out[16];
    assign wire_9484 = lut_tile_8_6_chanxy_out[17];
    assign wire_9486 = lut_tile_8_6_chanxy_out[18];
    assign wire_9488 = lut_tile_8_6_chanxy_out[19];
    assign wire_9490 = lut_tile_8_6_chanxy_out[20];
    assign wire_9492 = lut_tile_8_6_chanxy_out[21];
    assign wire_9494 = lut_tile_8_6_chanxy_out[22];
    assign wire_9496 = lut_tile_8_6_chanxy_out[23];
    assign wire_9498 = lut_tile_8_6_chanxy_out[24];
    assign wire_9500 = lut_tile_8_6_chanxy_out[25];
    assign wire_9502 = lut_tile_8_6_chanxy_out[26];
    assign wire_9504 = lut_tile_8_6_chanxy_out[27];
    assign wire_9506 = lut_tile_8_6_chanxy_out[28];
    assign wire_9508 = lut_tile_8_6_chanxy_out[29];
    assign wire_12961 = lut_tile_8_6_chanxy_out[30];
    assign wire_12963 = lut_tile_8_6_chanxy_out[31];
    assign wire_12965 = lut_tile_8_6_chanxy_out[32];
    assign wire_12967 = lut_tile_8_6_chanxy_out[33];
    assign wire_12969 = lut_tile_8_6_chanxy_out[34];
    assign wire_12971 = lut_tile_8_6_chanxy_out[35];
    assign wire_12973 = lut_tile_8_6_chanxy_out[36];
    assign wire_12975 = lut_tile_8_6_chanxy_out[37];
    assign wire_12977 = lut_tile_8_6_chanxy_out[38];
    assign wire_12979 = lut_tile_8_6_chanxy_out[39];
    assign wire_12981 = lut_tile_8_6_chanxy_out[40];
    assign wire_12983 = lut_tile_8_6_chanxy_out[41];
    assign wire_12985 = lut_tile_8_6_chanxy_out[42];
    assign wire_12987 = lut_tile_8_6_chanxy_out[43];
    assign wire_12989 = lut_tile_8_6_chanxy_out[44];
    assign wire_13050 = lut_tile_8_6_chanxy_out[45];
    assign wire_13052 = lut_tile_8_6_chanxy_out[46];
    assign wire_13054 = lut_tile_8_6_chanxy_out[47];
    assign wire_13056 = lut_tile_8_6_chanxy_out[48];
    assign wire_13058 = lut_tile_8_6_chanxy_out[49];
    assign wire_13060 = lut_tile_8_6_chanxy_out[50];
    assign wire_13062 = lut_tile_8_6_chanxy_out[51];
    assign wire_13064 = lut_tile_8_6_chanxy_out[52];
    assign wire_13066 = lut_tile_8_6_chanxy_out[53];
    assign wire_13068 = lut_tile_8_6_chanxy_out[54];
    assign wire_13070 = lut_tile_8_6_chanxy_out[55];
    assign wire_13072 = lut_tile_8_6_chanxy_out[56];
    assign wire_13074 = lut_tile_8_6_chanxy_out[57];
    assign wire_13076 = lut_tile_8_6_chanxy_out[58];
    assign wire_13078 = lut_tile_8_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_7_chanxy_in = {wire_13348, wire_9151, wire_9089, wire_9088, wire_9079, wire_9078, wire_9069, wire_9068, wire_9032, wire_4467, wire_13346, wire_9179, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9034, wire_4467, wire_13344, wire_9177, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9036, wire_4467, wire_13342, wire_9175, wire_9087, wire_9086, wire_9077, wire_9076, wire_9067, wire_9066, wire_9038, wire_3957, wire_13340, wire_9173, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9040, wire_3957, wire_13338, wire_9171, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9042, wire_3957, wire_13336, wire_9169, wire_9085, wire_9084, wire_9075, wire_9074, wire_9065, wire_9064, wire_9044, wire_4471, wire_3957, wire_13334, wire_9167, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9046, wire_4471, wire_3957, wire_13332, wire_9165, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9048, wire_4471, wire_3957, wire_13330, wire_9163, wire_9083, wire_9082, wire_9073, wire_9072, wire_9063, wire_9062, wire_9050, wire_4471, wire_3953, wire_13328, wire_9161, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9052, wire_4471, wire_3953, wire_13326, wire_9159, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9054, wire_4471, wire_3953, wire_13324, wire_9157, wire_9081, wire_9080, wire_9071, wire_9070, wire_9061, wire_9060, wire_9056, wire_4467, wire_3953, wire_13322, wire_9155, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9058, wire_4467, wire_3953, wire_13320, wire_9153, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9030, wire_4467, wire_3953, wire_13499, wire_9569, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9420, wire_4467, wire_13497, wire_9541, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9448, wire_4467, wire_13495, wire_9543, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9446, wire_4467, wire_13493, wire_9545, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9444, wire_3957, wire_13491, wire_9547, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9442, wire_3957, wire_13489, wire_9549, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9440, wire_3957, wire_13487, wire_9551, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9438, wire_4471, wire_3957, wire_13485, wire_9553, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9436, wire_4471, wire_3957, wire_13483, wire_9555, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9434, wire_4471, wire_3957, wire_13481, wire_9557, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9432, wire_4471, wire_3953, wire_13479, wire_9559, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9430, wire_4471, wire_3953, wire_13477, wire_9561, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9428, wire_4471, wire_3953, wire_13475, wire_9563, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9426, wire_4467, wire_3953, wire_13473, wire_9565, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9424, wire_4467, wire_3953, wire_13471, wire_9567, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9422, wire_4467, wire_3953, wire_13107, wire_13019, wire_13018, wire_13009, wire_13008, wire_12999, wire_12998, wire_12988, wire_9418, wire_3996, wire_13105, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_12960, wire_9416, wire_3996, wire_13103, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12962, wire_9414, wire_3996, wire_13101, wire_13017, wire_13016, wire_13007, wire_13006, wire_12997, wire_12996, wire_12964, wire_9412, wire_3956, wire_13099, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_12966, wire_9410, wire_3956, wire_13097, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12968, wire_9408, wire_3956, wire_13095, wire_13015, wire_13014, wire_13005, wire_13004, wire_12995, wire_12994, wire_12970, wire_9406, wire_4000, wire_3956, wire_13093, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_12972, wire_9404, wire_4000, wire_3956, wire_13091, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_12974, wire_9402, wire_4000, wire_3956, wire_13089, wire_13013, wire_13012, wire_13003, wire_13002, wire_12993, wire_12992, wire_12976, wire_9400, wire_4000, wire_3952, wire_13087, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_12978, wire_9398, wire_4000, wire_3952, wire_13085, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12980, wire_9396, wire_4000, wire_3952, wire_13083, wire_13011, wire_13010, wire_13001, wire_13000, wire_12991, wire_12990, wire_12982, wire_9394, wire_3996, wire_3952, wire_13081, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_12984, wire_9392, wire_3996, wire_3952, wire_13109, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_12986, wire_9390, wire_3996, wire_3952, wire_13473, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13376, wire_9569, wire_3996, wire_13475, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13374, wire_9567, wire_3996, wire_13477, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13372, wire_9565, wire_3996, wire_13479, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13370, wire_9563, wire_3956, wire_13481, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13368, wire_9561, wire_3956, wire_13483, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13366, wire_9559, wire_3956, wire_13485, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13364, wire_9557, wire_4000, wire_3956, wire_13487, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13362, wire_9555, wire_4000, wire_3956, wire_13489, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13360, wire_9553, wire_4000, wire_3956, wire_13491, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13358, wire_9551, wire_4000, wire_3952, wire_13493, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13356, wire_9549, wire_4000, wire_3952, wire_13495, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13354, wire_9547, wire_4000, wire_3952, wire_13497, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13352, wire_9545, wire_3996, wire_3952, wire_13499, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13350, wire_9543, wire_3996, wire_3952, wire_13471, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13378, wire_9541, wire_3996, wire_3952};
    // CHNAXY TOTAL: 636
    assign wire_9421 = lut_tile_8_7_chanxy_out[0];
    assign wire_9423 = lut_tile_8_7_chanxy_out[1];
    assign wire_9425 = lut_tile_8_7_chanxy_out[2];
    assign wire_9427 = lut_tile_8_7_chanxy_out[3];
    assign wire_9429 = lut_tile_8_7_chanxy_out[4];
    assign wire_9431 = lut_tile_8_7_chanxy_out[5];
    assign wire_9433 = lut_tile_8_7_chanxy_out[6];
    assign wire_9435 = lut_tile_8_7_chanxy_out[7];
    assign wire_9437 = lut_tile_8_7_chanxy_out[8];
    assign wire_9439 = lut_tile_8_7_chanxy_out[9];
    assign wire_9441 = lut_tile_8_7_chanxy_out[10];
    assign wire_9443 = lut_tile_8_7_chanxy_out[11];
    assign wire_9445 = lut_tile_8_7_chanxy_out[12];
    assign wire_9447 = lut_tile_8_7_chanxy_out[13];
    assign wire_9449 = lut_tile_8_7_chanxy_out[14];
    assign wire_9510 = lut_tile_8_7_chanxy_out[15];
    assign wire_9512 = lut_tile_8_7_chanxy_out[16];
    assign wire_9514 = lut_tile_8_7_chanxy_out[17];
    assign wire_9516 = lut_tile_8_7_chanxy_out[18];
    assign wire_9518 = lut_tile_8_7_chanxy_out[19];
    assign wire_9520 = lut_tile_8_7_chanxy_out[20];
    assign wire_9522 = lut_tile_8_7_chanxy_out[21];
    assign wire_9524 = lut_tile_8_7_chanxy_out[22];
    assign wire_9526 = lut_tile_8_7_chanxy_out[23];
    assign wire_9528 = lut_tile_8_7_chanxy_out[24];
    assign wire_9530 = lut_tile_8_7_chanxy_out[25];
    assign wire_9532 = lut_tile_8_7_chanxy_out[26];
    assign wire_9534 = lut_tile_8_7_chanxy_out[27];
    assign wire_9536 = lut_tile_8_7_chanxy_out[28];
    assign wire_9538 = lut_tile_8_7_chanxy_out[29];
    assign wire_13351 = lut_tile_8_7_chanxy_out[30];
    assign wire_13353 = lut_tile_8_7_chanxy_out[31];
    assign wire_13355 = lut_tile_8_7_chanxy_out[32];
    assign wire_13357 = lut_tile_8_7_chanxy_out[33];
    assign wire_13359 = lut_tile_8_7_chanxy_out[34];
    assign wire_13361 = lut_tile_8_7_chanxy_out[35];
    assign wire_13363 = lut_tile_8_7_chanxy_out[36];
    assign wire_13365 = lut_tile_8_7_chanxy_out[37];
    assign wire_13367 = lut_tile_8_7_chanxy_out[38];
    assign wire_13369 = lut_tile_8_7_chanxy_out[39];
    assign wire_13371 = lut_tile_8_7_chanxy_out[40];
    assign wire_13373 = lut_tile_8_7_chanxy_out[41];
    assign wire_13375 = lut_tile_8_7_chanxy_out[42];
    assign wire_13377 = lut_tile_8_7_chanxy_out[43];
    assign wire_13379 = lut_tile_8_7_chanxy_out[44];
    assign wire_13440 = lut_tile_8_7_chanxy_out[45];
    assign wire_13442 = lut_tile_8_7_chanxy_out[46];
    assign wire_13444 = lut_tile_8_7_chanxy_out[47];
    assign wire_13446 = lut_tile_8_7_chanxy_out[48];
    assign wire_13448 = lut_tile_8_7_chanxy_out[49];
    assign wire_13450 = lut_tile_8_7_chanxy_out[50];
    assign wire_13452 = lut_tile_8_7_chanxy_out[51];
    assign wire_13454 = lut_tile_8_7_chanxy_out[52];
    assign wire_13456 = lut_tile_8_7_chanxy_out[53];
    assign wire_13458 = lut_tile_8_7_chanxy_out[54];
    assign wire_13460 = lut_tile_8_7_chanxy_out[55];
    assign wire_13462 = lut_tile_8_7_chanxy_out[56];
    assign wire_13464 = lut_tile_8_7_chanxy_out[57];
    assign wire_13466 = lut_tile_8_7_chanxy_out[58];
    assign wire_13468 = lut_tile_8_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_8_chanxy_in = {wire_13738, wire_9181, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9062, wire_4983, wire_13736, wire_9209, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9064, wire_4983, wire_13734, wire_9207, wire_9119, wire_9118, wire_9109, wire_9108, wire_9099, wire_9098, wire_9066, wire_4983, wire_13732, wire_9205, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9068, wire_4473, wire_13730, wire_9203, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9070, wire_4473, wire_13728, wire_9201, wire_9117, wire_9116, wire_9107, wire_9106, wire_9097, wire_9096, wire_9072, wire_4473, wire_13726, wire_9199, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9074, wire_4987, wire_4473, wire_13724, wire_9197, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9076, wire_4987, wire_4473, wire_13722, wire_9195, wire_9115, wire_9114, wire_9105, wire_9104, wire_9095, wire_9094, wire_9078, wire_4987, wire_4473, wire_13720, wire_9193, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9080, wire_4987, wire_4469, wire_13718, wire_9191, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9082, wire_4987, wire_4469, wire_13716, wire_9189, wire_9113, wire_9112, wire_9103, wire_9102, wire_9093, wire_9092, wire_9084, wire_4987, wire_4469, wire_13714, wire_9187, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9086, wire_4983, wire_4469, wire_13712, wire_9185, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9088, wire_4983, wire_4469, wire_13710, wire_9183, wire_9111, wire_9110, wire_9101, wire_9100, wire_9091, wire_9090, wire_9060, wire_4983, wire_4469, wire_13889, wire_9599, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9450, wire_4983, wire_13887, wire_9571, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9478, wire_4983, wire_13885, wire_9573, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9476, wire_4983, wire_13883, wire_9575, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9474, wire_4473, wire_13881, wire_9577, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9472, wire_4473, wire_13879, wire_9579, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9470, wire_4473, wire_13877, wire_9581, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9468, wire_4987, wire_4473, wire_13875, wire_9583, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9466, wire_4987, wire_4473, wire_13873, wire_9585, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9464, wire_4987, wire_4473, wire_13871, wire_9587, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9462, wire_4987, wire_4469, wire_13869, wire_9589, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9460, wire_4987, wire_4469, wire_13867, wire_9591, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9458, wire_4987, wire_4469, wire_13865, wire_9593, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9456, wire_4983, wire_4469, wire_13863, wire_9595, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9454, wire_4983, wire_4469, wire_13861, wire_9597, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9452, wire_4983, wire_4469, wire_13497, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13378, wire_9448, wire_4512, wire_13495, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13350, wire_9446, wire_4512, wire_13493, wire_13409, wire_13408, wire_13399, wire_13398, wire_13389, wire_13388, wire_13352, wire_9444, wire_4512, wire_13491, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13354, wire_9442, wire_4472, wire_13489, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13356, wire_9440, wire_4472, wire_13487, wire_13407, wire_13406, wire_13397, wire_13396, wire_13387, wire_13386, wire_13358, wire_9438, wire_4472, wire_13485, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13360, wire_9436, wire_4516, wire_4472, wire_13483, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13362, wire_9434, wire_4516, wire_4472, wire_13481, wire_13405, wire_13404, wire_13395, wire_13394, wire_13385, wire_13384, wire_13364, wire_9432, wire_4516, wire_4472, wire_13479, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13366, wire_9430, wire_4516, wire_4468, wire_13477, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13368, wire_9428, wire_4516, wire_4468, wire_13475, wire_13403, wire_13402, wire_13393, wire_13392, wire_13383, wire_13382, wire_13370, wire_9426, wire_4516, wire_4468, wire_13473, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13372, wire_9424, wire_4512, wire_4468, wire_13471, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13374, wire_9422, wire_4512, wire_4468, wire_13499, wire_13401, wire_13400, wire_13391, wire_13390, wire_13381, wire_13380, wire_13376, wire_9420, wire_4512, wire_4468, wire_13863, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13766, wire_9599, wire_4512, wire_13865, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13764, wire_9597, wire_4512, wire_13867, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13762, wire_9595, wire_4512, wire_13869, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13760, wire_9593, wire_4472, wire_13871, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13758, wire_9591, wire_4472, wire_13873, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13756, wire_9589, wire_4472, wire_13875, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13754, wire_9587, wire_4516, wire_4472, wire_13877, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13752, wire_9585, wire_4516, wire_4472, wire_13879, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13750, wire_9583, wire_4516, wire_4472, wire_13881, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13748, wire_9581, wire_4516, wire_4468, wire_13883, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13746, wire_9579, wire_4516, wire_4468, wire_13885, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13744, wire_9577, wire_4516, wire_4468, wire_13887, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13742, wire_9575, wire_4512, wire_4468, wire_13889, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13740, wire_9573, wire_4512, wire_4468, wire_13861, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13768, wire_9571, wire_4512, wire_4468};
    // CHNAXY TOTAL: 636
    assign wire_9451 = lut_tile_8_8_chanxy_out[0];
    assign wire_9453 = lut_tile_8_8_chanxy_out[1];
    assign wire_9455 = lut_tile_8_8_chanxy_out[2];
    assign wire_9457 = lut_tile_8_8_chanxy_out[3];
    assign wire_9459 = lut_tile_8_8_chanxy_out[4];
    assign wire_9461 = lut_tile_8_8_chanxy_out[5];
    assign wire_9463 = lut_tile_8_8_chanxy_out[6];
    assign wire_9465 = lut_tile_8_8_chanxy_out[7];
    assign wire_9467 = lut_tile_8_8_chanxy_out[8];
    assign wire_9469 = lut_tile_8_8_chanxy_out[9];
    assign wire_9471 = lut_tile_8_8_chanxy_out[10];
    assign wire_9473 = lut_tile_8_8_chanxy_out[11];
    assign wire_9475 = lut_tile_8_8_chanxy_out[12];
    assign wire_9477 = lut_tile_8_8_chanxy_out[13];
    assign wire_9479 = lut_tile_8_8_chanxy_out[14];
    assign wire_9540 = lut_tile_8_8_chanxy_out[15];
    assign wire_9542 = lut_tile_8_8_chanxy_out[16];
    assign wire_9544 = lut_tile_8_8_chanxy_out[17];
    assign wire_9546 = lut_tile_8_8_chanxy_out[18];
    assign wire_9548 = lut_tile_8_8_chanxy_out[19];
    assign wire_9550 = lut_tile_8_8_chanxy_out[20];
    assign wire_9552 = lut_tile_8_8_chanxy_out[21];
    assign wire_9554 = lut_tile_8_8_chanxy_out[22];
    assign wire_9556 = lut_tile_8_8_chanxy_out[23];
    assign wire_9558 = lut_tile_8_8_chanxy_out[24];
    assign wire_9560 = lut_tile_8_8_chanxy_out[25];
    assign wire_9562 = lut_tile_8_8_chanxy_out[26];
    assign wire_9564 = lut_tile_8_8_chanxy_out[27];
    assign wire_9566 = lut_tile_8_8_chanxy_out[28];
    assign wire_9568 = lut_tile_8_8_chanxy_out[29];
    assign wire_13741 = lut_tile_8_8_chanxy_out[30];
    assign wire_13743 = lut_tile_8_8_chanxy_out[31];
    assign wire_13745 = lut_tile_8_8_chanxy_out[32];
    assign wire_13747 = lut_tile_8_8_chanxy_out[33];
    assign wire_13749 = lut_tile_8_8_chanxy_out[34];
    assign wire_13751 = lut_tile_8_8_chanxy_out[35];
    assign wire_13753 = lut_tile_8_8_chanxy_out[36];
    assign wire_13755 = lut_tile_8_8_chanxy_out[37];
    assign wire_13757 = lut_tile_8_8_chanxy_out[38];
    assign wire_13759 = lut_tile_8_8_chanxy_out[39];
    assign wire_13761 = lut_tile_8_8_chanxy_out[40];
    assign wire_13763 = lut_tile_8_8_chanxy_out[41];
    assign wire_13765 = lut_tile_8_8_chanxy_out[42];
    assign wire_13767 = lut_tile_8_8_chanxy_out[43];
    assign wire_13769 = lut_tile_8_8_chanxy_out[44];
    assign wire_13830 = lut_tile_8_8_chanxy_out[45];
    assign wire_13832 = lut_tile_8_8_chanxy_out[46];
    assign wire_13834 = lut_tile_8_8_chanxy_out[47];
    assign wire_13836 = lut_tile_8_8_chanxy_out[48];
    assign wire_13838 = lut_tile_8_8_chanxy_out[49];
    assign wire_13840 = lut_tile_8_8_chanxy_out[50];
    assign wire_13842 = lut_tile_8_8_chanxy_out[51];
    assign wire_13844 = lut_tile_8_8_chanxy_out[52];
    assign wire_13846 = lut_tile_8_8_chanxy_out[53];
    assign wire_13848 = lut_tile_8_8_chanxy_out[54];
    assign wire_13850 = lut_tile_8_8_chanxy_out[55];
    assign wire_13852 = lut_tile_8_8_chanxy_out[56];
    assign wire_13854 = lut_tile_8_8_chanxy_out[57];
    assign wire_13856 = lut_tile_8_8_chanxy_out[58];
    assign wire_13858 = lut_tile_8_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_9_chanxy_in = {wire_14128, wire_9211, wire_9209, wire_9208, wire_9199, wire_9198, wire_9189, wire_9188, wire_9092, wire_5499, wire_14126, wire_9239, wire_9179, wire_9178, wire_9169, wire_9168, wire_9159, wire_9158, wire_9094, wire_5499, wire_14124, wire_9237, wire_9149, wire_9148, wire_9139, wire_9138, wire_9129, wire_9128, wire_9096, wire_5499, wire_14122, wire_9235, wire_9207, wire_9206, wire_9197, wire_9196, wire_9187, wire_9186, wire_9098, wire_4989, wire_14120, wire_9233, wire_9177, wire_9176, wire_9167, wire_9166, wire_9157, wire_9156, wire_9100, wire_4989, wire_14118, wire_9231, wire_9147, wire_9146, wire_9137, wire_9136, wire_9127, wire_9126, wire_9102, wire_4989, wire_14116, wire_9229, wire_9205, wire_9204, wire_9195, wire_9194, wire_9185, wire_9184, wire_9104, wire_5503, wire_4989, wire_14114, wire_9227, wire_9175, wire_9174, wire_9165, wire_9164, wire_9155, wire_9154, wire_9106, wire_5503, wire_4989, wire_14112, wire_9225, wire_9145, wire_9144, wire_9135, wire_9134, wire_9125, wire_9124, wire_9108, wire_5503, wire_4989, wire_14110, wire_9223, wire_9203, wire_9202, wire_9193, wire_9192, wire_9183, wire_9182, wire_9110, wire_5503, wire_4985, wire_14108, wire_9221, wire_9173, wire_9172, wire_9163, wire_9162, wire_9153, wire_9152, wire_9112, wire_5503, wire_4985, wire_14106, wire_9219, wire_9143, wire_9142, wire_9133, wire_9132, wire_9123, wire_9122, wire_9114, wire_5503, wire_4985, wire_14104, wire_9217, wire_9201, wire_9200, wire_9191, wire_9190, wire_9181, wire_9180, wire_9116, wire_5499, wire_4985, wire_14102, wire_9215, wire_9171, wire_9170, wire_9161, wire_9160, wire_9151, wire_9150, wire_9118, wire_5499, wire_4985, wire_14100, wire_9213, wire_9141, wire_9140, wire_9131, wire_9130, wire_9121, wire_9120, wire_9090, wire_5499, wire_4985, wire_14279, wire_9629, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9480, wire_5499, wire_14277, wire_9601, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9508, wire_5499, wire_14275, wire_9603, wire_9599, wire_9598, wire_9589, wire_9588, wire_9579, wire_9578, wire_9506, wire_5499, wire_14273, wire_9605, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9504, wire_4989, wire_14271, wire_9607, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9502, wire_4989, wire_14269, wire_9609, wire_9597, wire_9596, wire_9587, wire_9586, wire_9577, wire_9576, wire_9500, wire_4989, wire_14267, wire_9611, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9498, wire_5503, wire_4989, wire_14265, wire_9613, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9496, wire_5503, wire_4989, wire_14263, wire_9615, wire_9595, wire_9594, wire_9585, wire_9584, wire_9575, wire_9574, wire_9494, wire_5503, wire_4989, wire_14261, wire_9617, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9492, wire_5503, wire_4985, wire_14259, wire_9619, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9490, wire_5503, wire_4985, wire_14257, wire_9621, wire_9593, wire_9592, wire_9583, wire_9582, wire_9573, wire_9572, wire_9488, wire_5503, wire_4985, wire_14255, wire_9623, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9486, wire_5499, wire_4985, wire_14253, wire_9625, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9484, wire_5499, wire_4985, wire_14251, wire_9627, wire_9591, wire_9590, wire_9581, wire_9580, wire_9571, wire_9570, wire_9482, wire_5499, wire_4985, wire_13887, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13768, wire_9478, wire_5028, wire_13885, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13740, wire_9476, wire_5028, wire_13883, wire_13799, wire_13798, wire_13789, wire_13788, wire_13779, wire_13778, wire_13742, wire_9474, wire_5028, wire_13881, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13744, wire_9472, wire_4988, wire_13879, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13746, wire_9470, wire_4988, wire_13877, wire_13797, wire_13796, wire_13787, wire_13786, wire_13777, wire_13776, wire_13748, wire_9468, wire_4988, wire_13875, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13750, wire_9466, wire_5032, wire_4988, wire_13873, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13752, wire_9464, wire_5032, wire_4988, wire_13871, wire_13795, wire_13794, wire_13785, wire_13784, wire_13775, wire_13774, wire_13754, wire_9462, wire_5032, wire_4988, wire_13869, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13756, wire_9460, wire_5032, wire_4984, wire_13867, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13758, wire_9458, wire_5032, wire_4984, wire_13865, wire_13793, wire_13792, wire_13783, wire_13782, wire_13773, wire_13772, wire_13760, wire_9456, wire_5032, wire_4984, wire_13863, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13762, wire_9454, wire_5028, wire_4984, wire_13861, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13764, wire_9452, wire_5028, wire_4984, wire_13889, wire_13791, wire_13790, wire_13781, wire_13780, wire_13771, wire_13770, wire_13766, wire_9450, wire_5028, wire_4984, wire_14253, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14156, wire_9629, wire_5028, wire_14255, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14154, wire_9627, wire_5028, wire_14257, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14152, wire_9625, wire_5028, wire_14259, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14150, wire_9623, wire_4988, wire_14261, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14148, wire_9621, wire_4988, wire_14263, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14146, wire_9619, wire_4988, wire_14265, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14144, wire_9617, wire_5032, wire_4988, wire_14267, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14142, wire_9615, wire_5032, wire_4988, wire_14269, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14140, wire_9613, wire_5032, wire_4988, wire_14271, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14138, wire_9611, wire_5032, wire_4984, wire_14273, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14136, wire_9609, wire_5032, wire_4984, wire_14275, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14134, wire_9607, wire_5032, wire_4984, wire_14277, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14132, wire_9605, wire_5028, wire_4984, wire_14279, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14130, wire_9603, wire_5028, wire_4984, wire_14251, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14158, wire_9601, wire_5028, wire_4984};
    // CHNAXY TOTAL: 636
    assign wire_9481 = lut_tile_8_9_chanxy_out[0];
    assign wire_9483 = lut_tile_8_9_chanxy_out[1];
    assign wire_9485 = lut_tile_8_9_chanxy_out[2];
    assign wire_9487 = lut_tile_8_9_chanxy_out[3];
    assign wire_9489 = lut_tile_8_9_chanxy_out[4];
    assign wire_9491 = lut_tile_8_9_chanxy_out[5];
    assign wire_9493 = lut_tile_8_9_chanxy_out[6];
    assign wire_9495 = lut_tile_8_9_chanxy_out[7];
    assign wire_9497 = lut_tile_8_9_chanxy_out[8];
    assign wire_9499 = lut_tile_8_9_chanxy_out[9];
    assign wire_9501 = lut_tile_8_9_chanxy_out[10];
    assign wire_9503 = lut_tile_8_9_chanxy_out[11];
    assign wire_9505 = lut_tile_8_9_chanxy_out[12];
    assign wire_9507 = lut_tile_8_9_chanxy_out[13];
    assign wire_9509 = lut_tile_8_9_chanxy_out[14];
    assign wire_9570 = lut_tile_8_9_chanxy_out[15];
    assign wire_9572 = lut_tile_8_9_chanxy_out[16];
    assign wire_9574 = lut_tile_8_9_chanxy_out[17];
    assign wire_9576 = lut_tile_8_9_chanxy_out[18];
    assign wire_9578 = lut_tile_8_9_chanxy_out[19];
    assign wire_9580 = lut_tile_8_9_chanxy_out[20];
    assign wire_9582 = lut_tile_8_9_chanxy_out[21];
    assign wire_9584 = lut_tile_8_9_chanxy_out[22];
    assign wire_9586 = lut_tile_8_9_chanxy_out[23];
    assign wire_9588 = lut_tile_8_9_chanxy_out[24];
    assign wire_9590 = lut_tile_8_9_chanxy_out[25];
    assign wire_9592 = lut_tile_8_9_chanxy_out[26];
    assign wire_9594 = lut_tile_8_9_chanxy_out[27];
    assign wire_9596 = lut_tile_8_9_chanxy_out[28];
    assign wire_9598 = lut_tile_8_9_chanxy_out[29];
    assign wire_14131 = lut_tile_8_9_chanxy_out[30];
    assign wire_14133 = lut_tile_8_9_chanxy_out[31];
    assign wire_14135 = lut_tile_8_9_chanxy_out[32];
    assign wire_14137 = lut_tile_8_9_chanxy_out[33];
    assign wire_14139 = lut_tile_8_9_chanxy_out[34];
    assign wire_14141 = lut_tile_8_9_chanxy_out[35];
    assign wire_14143 = lut_tile_8_9_chanxy_out[36];
    assign wire_14145 = lut_tile_8_9_chanxy_out[37];
    assign wire_14147 = lut_tile_8_9_chanxy_out[38];
    assign wire_14149 = lut_tile_8_9_chanxy_out[39];
    assign wire_14151 = lut_tile_8_9_chanxy_out[40];
    assign wire_14153 = lut_tile_8_9_chanxy_out[41];
    assign wire_14155 = lut_tile_8_9_chanxy_out[42];
    assign wire_14157 = lut_tile_8_9_chanxy_out[43];
    assign wire_14159 = lut_tile_8_9_chanxy_out[44];
    assign wire_14220 = lut_tile_8_9_chanxy_out[45];
    assign wire_14222 = lut_tile_8_9_chanxy_out[46];
    assign wire_14224 = lut_tile_8_9_chanxy_out[47];
    assign wire_14226 = lut_tile_8_9_chanxy_out[48];
    assign wire_14228 = lut_tile_8_9_chanxy_out[49];
    assign wire_14230 = lut_tile_8_9_chanxy_out[50];
    assign wire_14232 = lut_tile_8_9_chanxy_out[51];
    assign wire_14234 = lut_tile_8_9_chanxy_out[52];
    assign wire_14236 = lut_tile_8_9_chanxy_out[53];
    assign wire_14238 = lut_tile_8_9_chanxy_out[54];
    assign wire_14240 = lut_tile_8_9_chanxy_out[55];
    assign wire_14242 = lut_tile_8_9_chanxy_out[56];
    assign wire_14244 = lut_tile_8_9_chanxy_out[57];
    assign wire_14246 = lut_tile_8_9_chanxy_out[58];
    assign wire_14248 = lut_tile_8_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_8_10_chanxy_in = {wire_14518, wire_9232, wire_9208, wire_9156, wire_9134, wire_6022, wire_6016, wire_6007, wire_6001, wire_14516, wire_9224, wire_9200, wire_9178, wire_9126, wire_6022, wire_6016, wire_6007, wire_6001, wire_14514, wire_9216, wire_9192, wire_9170, wire_9148, wire_6022, wire_6016, wire_6007, wire_6001, wire_14512, wire_9238, wire_9184, wire_9162, wire_9140, wire_6022, wire_6013, wire_6007, wire_5505, wire_14510, wire_9230, wire_9206, wire_9154, wire_9132, wire_6022, wire_6013, wire_6007, wire_5505, wire_14508, wire_9222, wire_9198, wire_9176, wire_9124, wire_6022, wire_6013, wire_6007, wire_5505, wire_14506, wire_9214, wire_9190, wire_9168, wire_9146, wire_6019, wire_6013, wire_6004, wire_5505, wire_14504, wire_9236, wire_9182, wire_9160, wire_9138, wire_6019, wire_6013, wire_6004, wire_5505, wire_14502, wire_9228, wire_9204, wire_9152, wire_9130, wire_6019, wire_6013, wire_6004, wire_5505, wire_14500, wire_9220, wire_9196, wire_9174, wire_9122, wire_6019, wire_6010, wire_6004, wire_5501, wire_14498, wire_9212, wire_9188, wire_9166, wire_9144, wire_6019, wire_6010, wire_6004, wire_5501, wire_14496, wire_9234, wire_9180, wire_9158, wire_9136, wire_6019, wire_6010, wire_6004, wire_5501, wire_14494, wire_9226, wire_9202, wire_9150, wire_9128, wire_6016, wire_6010, wire_6001, wire_5501, wire_14492, wire_9218, wire_9194, wire_9172, wire_9120, wire_6016, wire_6010, wire_6001, wire_5501, wire_14490, wire_9210, wire_9186, wire_9164, wire_9142, wire_6016, wire_6010, wire_6001, wire_5501, wire_14669, wire_9614, wire_9592, wire_9568, wire_9516, wire_6022, wire_6016, wire_6007, wire_6001, wire_14667, wire_9606, wire_9584, wire_9560, wire_9538, wire_6022, wire_6016, wire_6007, wire_6001, wire_14665, wire_9628, wire_9576, wire_9552, wire_9530, wire_6022, wire_6016, wire_6007, wire_6001, wire_14663, wire_9620, wire_9598, wire_9544, wire_9522, wire_6022, wire_6013, wire_6007, wire_5505, wire_14661, wire_9612, wire_9590, wire_9566, wire_9514, wire_6022, wire_6013, wire_6007, wire_5505, wire_14659, wire_9604, wire_9582, wire_9558, wire_9536, wire_6022, wire_6013, wire_6007, wire_5505, wire_14657, wire_9626, wire_9574, wire_9550, wire_9528, wire_6019, wire_6013, wire_6004, wire_5505, wire_14655, wire_9618, wire_9596, wire_9542, wire_9520, wire_6019, wire_6013, wire_6004, wire_5505, wire_14653, wire_9610, wire_9588, wire_9564, wire_9512, wire_6019, wire_6013, wire_6004, wire_5505, wire_14651, wire_9602, wire_9580, wire_9556, wire_9534, wire_6019, wire_6010, wire_6004, wire_5501, wire_14649, wire_9624, wire_9572, wire_9548, wire_9526, wire_6019, wire_6010, wire_6004, wire_5501, wire_14647, wire_9616, wire_9594, wire_9540, wire_9518, wire_6019, wire_6010, wire_6004, wire_5501, wire_14645, wire_9608, wire_9586, wire_9562, wire_9510, wire_6016, wire_6010, wire_6001, wire_5501, wire_14643, wire_9600, wire_9578, wire_9554, wire_9532, wire_6016, wire_6010, wire_6001, wire_5501, wire_14641, wire_9622, wire_9570, wire_9546, wire_9524, wire_6016, wire_6010, wire_6001, wire_5501, wire_14563, wire_14562, wire_14277, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14158, wire_9508, wire_5544, wire_14577, wire_14576, wire_14275, wire_14189, wire_14188, wire_14179, wire_14178, wire_14169, wire_14168, wire_14130, wire_9506, wire_5544, wire_14607, wire_14606, wire_14273, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14132, wire_9504, wire_5544, wire_14575, wire_14574, wire_14271, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14134, wire_9502, wire_5504, wire_14559, wire_14558, wire_14269, wire_14187, wire_14186, wire_14177, wire_14176, wire_14167, wire_14166, wire_14136, wire_9500, wire_5504, wire_14589, wire_14588, wire_14267, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14138, wire_9498, wire_5504, wire_14557, wire_14556, wire_14265, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14140, wire_9496, wire_5548, wire_5504, wire_14571, wire_14570, wire_14263, wire_14185, wire_14184, wire_14175, wire_14174, wire_14165, wire_14164, wire_14142, wire_9494, wire_5548, wire_5504, wire_14601, wire_14600, wire_14261, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14144, wire_9492, wire_5548, wire_5504, wire_14569, wire_14568, wire_5548, wire_14259, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14146, wire_9490, wire_5548, wire_5500, wire_14553, wire_14552, wire_5544, wire_14257, wire_14183, wire_14182, wire_14173, wire_14172, wire_14163, wire_14162, wire_14148, wire_9488, wire_5548, wire_5500, wire_14583, wire_14582, wire_5544, wire_14255, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14150, wire_9486, wire_5548, wire_5500, wire_14551, wire_14550, wire_5504, wire_14253, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14152, wire_9484, wire_5544, wire_5500, wire_14565, wire_14564, wire_5500, wire_14251, wire_14181, wire_14180, wire_14171, wire_14170, wire_14161, wire_14160, wire_14154, wire_9482, wire_5544, wire_5500, wire_14595, wire_14594, wire_5500, wire_14279, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14156, wire_9480, wire_5544, wire_5500, wire_14639, wire_14638, wire_14667, wire_14546, wire_14593, wire_14592, wire_14621, wire_14620, wire_14649, wire_14528, wire_14605, wire_14604, wire_14633, wire_14632, wire_14661, wire_14540, wire_14587, wire_14586, wire_14615, wire_14614, wire_5548, wire_14643, wire_14522, wire_5544, wire_14599, wire_14598, wire_5544, wire_14627, wire_14626, wire_5504, wire_14655, wire_14534, wire_5500, wire_14581, wire_14580, wire_5500, wire_14579, wire_14578, wire_14609, wire_14608, wire_14623, wire_14622, wire_14561, wire_14560, wire_14591, wire_14590, wire_14635, wire_14634, wire_14573, wire_14572, wire_14603, wire_14602, wire_14617, wire_14616, wire_14555, wire_14554, wire_5548, wire_14585, wire_14584, wire_5548, wire_14629, wire_14628, wire_5544, wire_14567, wire_14566, wire_5504, wire_14597, wire_14596, wire_5504, wire_14611, wire_14610, wire_5500, wire_14669, wire_14548, wire_14653, wire_14532, wire_14637, wire_14636, wire_14651, wire_14530, wire_14665, wire_14544, wire_14619, wire_14618, wire_14663, wire_14542, wire_14647, wire_14526, wire_14631, wire_14630, wire_14645, wire_14524, wire_5548, wire_14659, wire_14538, wire_5548, wire_14613, wire_14612, wire_5544, wire_14657, wire_14536, wire_5504, wire_14641, wire_14520, wire_5504, wire_14625, wire_14624, wire_5500};
    // CHNAXY TOTAL: 573
    assign wire_9511 = lut_tile_8_10_chanxy_out[0];
    assign wire_9513 = lut_tile_8_10_chanxy_out[1];
    assign wire_9515 = lut_tile_8_10_chanxy_out[2];
    assign wire_9517 = lut_tile_8_10_chanxy_out[3];
    assign wire_9519 = lut_tile_8_10_chanxy_out[4];
    assign wire_9521 = lut_tile_8_10_chanxy_out[5];
    assign wire_9523 = lut_tile_8_10_chanxy_out[6];
    assign wire_9525 = lut_tile_8_10_chanxy_out[7];
    assign wire_9527 = lut_tile_8_10_chanxy_out[8];
    assign wire_9529 = lut_tile_8_10_chanxy_out[9];
    assign wire_9531 = lut_tile_8_10_chanxy_out[10];
    assign wire_9533 = lut_tile_8_10_chanxy_out[11];
    assign wire_9535 = lut_tile_8_10_chanxy_out[12];
    assign wire_9537 = lut_tile_8_10_chanxy_out[13];
    assign wire_9539 = lut_tile_8_10_chanxy_out[14];
    assign wire_9541 = lut_tile_8_10_chanxy_out[15];
    assign wire_9543 = lut_tile_8_10_chanxy_out[16];
    assign wire_9545 = lut_tile_8_10_chanxy_out[17];
    assign wire_9547 = lut_tile_8_10_chanxy_out[18];
    assign wire_9549 = lut_tile_8_10_chanxy_out[19];
    assign wire_9551 = lut_tile_8_10_chanxy_out[20];
    assign wire_9553 = lut_tile_8_10_chanxy_out[21];
    assign wire_9555 = lut_tile_8_10_chanxy_out[22];
    assign wire_9557 = lut_tile_8_10_chanxy_out[23];
    assign wire_9559 = lut_tile_8_10_chanxy_out[24];
    assign wire_9561 = lut_tile_8_10_chanxy_out[25];
    assign wire_9563 = lut_tile_8_10_chanxy_out[26];
    assign wire_9565 = lut_tile_8_10_chanxy_out[27];
    assign wire_9567 = lut_tile_8_10_chanxy_out[28];
    assign wire_9569 = lut_tile_8_10_chanxy_out[29];
    assign wire_9571 = lut_tile_8_10_chanxy_out[30];
    assign wire_9573 = lut_tile_8_10_chanxy_out[31];
    assign wire_9575 = lut_tile_8_10_chanxy_out[32];
    assign wire_9577 = lut_tile_8_10_chanxy_out[33];
    assign wire_9579 = lut_tile_8_10_chanxy_out[34];
    assign wire_9581 = lut_tile_8_10_chanxy_out[35];
    assign wire_9583 = lut_tile_8_10_chanxy_out[36];
    assign wire_9585 = lut_tile_8_10_chanxy_out[37];
    assign wire_9587 = lut_tile_8_10_chanxy_out[38];
    assign wire_9589 = lut_tile_8_10_chanxy_out[39];
    assign wire_9591 = lut_tile_8_10_chanxy_out[40];
    assign wire_9593 = lut_tile_8_10_chanxy_out[41];
    assign wire_9595 = lut_tile_8_10_chanxy_out[42];
    assign wire_9597 = lut_tile_8_10_chanxy_out[43];
    assign wire_9599 = lut_tile_8_10_chanxy_out[44];
    assign wire_9600 = lut_tile_8_10_chanxy_out[45];
    assign wire_9601 = lut_tile_8_10_chanxy_out[46];
    assign wire_9602 = lut_tile_8_10_chanxy_out[47];
    assign wire_9603 = lut_tile_8_10_chanxy_out[48];
    assign wire_9604 = lut_tile_8_10_chanxy_out[49];
    assign wire_9605 = lut_tile_8_10_chanxy_out[50];
    assign wire_9606 = lut_tile_8_10_chanxy_out[51];
    assign wire_9607 = lut_tile_8_10_chanxy_out[52];
    assign wire_9608 = lut_tile_8_10_chanxy_out[53];
    assign wire_9609 = lut_tile_8_10_chanxy_out[54];
    assign wire_9610 = lut_tile_8_10_chanxy_out[55];
    assign wire_9611 = lut_tile_8_10_chanxy_out[56];
    assign wire_9612 = lut_tile_8_10_chanxy_out[57];
    assign wire_9613 = lut_tile_8_10_chanxy_out[58];
    assign wire_9614 = lut_tile_8_10_chanxy_out[59];
    assign wire_9615 = lut_tile_8_10_chanxy_out[60];
    assign wire_9616 = lut_tile_8_10_chanxy_out[61];
    assign wire_9617 = lut_tile_8_10_chanxy_out[62];
    assign wire_9618 = lut_tile_8_10_chanxy_out[63];
    assign wire_9619 = lut_tile_8_10_chanxy_out[64];
    assign wire_9620 = lut_tile_8_10_chanxy_out[65];
    assign wire_9621 = lut_tile_8_10_chanxy_out[66];
    assign wire_9622 = lut_tile_8_10_chanxy_out[67];
    assign wire_9623 = lut_tile_8_10_chanxy_out[68];
    assign wire_9624 = lut_tile_8_10_chanxy_out[69];
    assign wire_9625 = lut_tile_8_10_chanxy_out[70];
    assign wire_9626 = lut_tile_8_10_chanxy_out[71];
    assign wire_9627 = lut_tile_8_10_chanxy_out[72];
    assign wire_9628 = lut_tile_8_10_chanxy_out[73];
    assign wire_9629 = lut_tile_8_10_chanxy_out[74];
    assign wire_14521 = lut_tile_8_10_chanxy_out[75];
    assign wire_14523 = lut_tile_8_10_chanxy_out[76];
    assign wire_14525 = lut_tile_8_10_chanxy_out[77];
    assign wire_14527 = lut_tile_8_10_chanxy_out[78];
    assign wire_14529 = lut_tile_8_10_chanxy_out[79];
    assign wire_14531 = lut_tile_8_10_chanxy_out[80];
    assign wire_14533 = lut_tile_8_10_chanxy_out[81];
    assign wire_14535 = lut_tile_8_10_chanxy_out[82];
    assign wire_14537 = lut_tile_8_10_chanxy_out[83];
    assign wire_14539 = lut_tile_8_10_chanxy_out[84];
    assign wire_14541 = lut_tile_8_10_chanxy_out[85];
    assign wire_14543 = lut_tile_8_10_chanxy_out[86];
    assign wire_14545 = lut_tile_8_10_chanxy_out[87];
    assign wire_14547 = lut_tile_8_10_chanxy_out[88];
    assign wire_14549 = lut_tile_8_10_chanxy_out[89];
    assign wire_14610 = lut_tile_8_10_chanxy_out[90];
    assign wire_14612 = lut_tile_8_10_chanxy_out[91];
    assign wire_14614 = lut_tile_8_10_chanxy_out[92];
    assign wire_14616 = lut_tile_8_10_chanxy_out[93];
    assign wire_14618 = lut_tile_8_10_chanxy_out[94];
    assign wire_14620 = lut_tile_8_10_chanxy_out[95];
    assign wire_14622 = lut_tile_8_10_chanxy_out[96];
    assign wire_14624 = lut_tile_8_10_chanxy_out[97];
    assign wire_14626 = lut_tile_8_10_chanxy_out[98];
    assign wire_14628 = lut_tile_8_10_chanxy_out[99];
    assign wire_14630 = lut_tile_8_10_chanxy_out[100];
    assign wire_14632 = lut_tile_8_10_chanxy_out[101];
    assign wire_14634 = lut_tile_8_10_chanxy_out[102];
    assign wire_14636 = lut_tile_8_10_chanxy_out[103];
    assign wire_14638 = lut_tile_8_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_9_1_chanxy_in = {wire_11038, wire_9361, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_9250, wire_1413, wire_11036, wire_9389, wire_9357, wire_9356, wire_9317, wire_9316, wire_9277, wire_9276, wire_9258, wire_1413, wire_11034, wire_9387, wire_9353, wire_9352, wire_9313, wire_9312, wire_9273, wire_9272, wire_9266, wire_1413, wire_11032, wire_9385, wire_9351, wire_9350, wire_9311, wire_9310, wire_9274, wire_9271, wire_9270, wire_903, wire_11030, wire_9383, wire_9349, wire_9348, wire_9309, wire_9308, wire_9282, wire_9269, wire_9268, wire_903, wire_11028, wire_9381, wire_9345, wire_9344, wire_9305, wire_9304, wire_9290, wire_9265, wire_9264, wire_903, wire_11026, wire_9379, wire_9343, wire_9342, wire_9303, wire_9302, wire_9298, wire_9263, wire_9262, wire_1417, wire_903, wire_11024, wire_9377, wire_9341, wire_9340, wire_9306, wire_9301, wire_9300, wire_9261, wire_9260, wire_1417, wire_903, wire_11022, wire_9375, wire_9337, wire_9336, wire_9314, wire_9297, wire_9296, wire_9257, wire_9256, wire_1417, wire_903, wire_11020, wire_9373, wire_9335, wire_9334, wire_9322, wire_9295, wire_9294, wire_9255, wire_9254, wire_1417, wire_899, wire_11018, wire_9371, wire_9333, wire_9332, wire_9330, wire_9293, wire_9292, wire_9253, wire_9252, wire_1417, wire_899, wire_11016, wire_9369, wire_9338, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_1417, wire_899, wire_11014, wire_9367, wire_9346, wire_9327, wire_9326, wire_9287, wire_9286, wire_9247, wire_9246, wire_1413, wire_899, wire_11012, wire_9365, wire_9354, wire_9325, wire_9324, wire_9285, wire_9284, wire_9245, wire_9244, wire_1413, wire_899, wire_11010, wire_9363, wire_9321, wire_9320, wire_9281, wire_9280, wire_9242, wire_9241, wire_9240, wire_1413, wire_899, wire_11189, wire_9779, wire_9749, wire_9748, wire_9709, wire_9708, wire_9669, wire_9668, wire_9634, wire_1413, wire_11187, wire_9751, wire_9746, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_1413, wire_11185, wire_9753, wire_9743, wire_9742, wire_9738, wire_9703, wire_9702, wire_9663, wire_9662, wire_1413, wire_11183, wire_9755, wire_9741, wire_9740, wire_9730, wire_9701, wire_9700, wire_9661, wire_9660, wire_903, wire_11181, wire_9757, wire_9737, wire_9736, wire_9722, wire_9697, wire_9696, wire_9657, wire_9656, wire_903, wire_11179, wire_9759, wire_9735, wire_9734, wire_9714, wire_9695, wire_9694, wire_9655, wire_9654, wire_903, wire_11177, wire_9761, wire_9733, wire_9732, wire_9706, wire_9693, wire_9692, wire_9653, wire_9652, wire_1417, wire_903, wire_11175, wire_9763, wire_9729, wire_9728, wire_9698, wire_9689, wire_9688, wire_9649, wire_9648, wire_1417, wire_903, wire_11173, wire_9765, wire_9727, wire_9726, wire_9690, wire_9687, wire_9686, wire_9647, wire_9646, wire_1417, wire_903, wire_11171, wire_9767, wire_9725, wire_9724, wire_9685, wire_9684, wire_9682, wire_9645, wire_9644, wire_1417, wire_899, wire_11169, wire_9769, wire_9721, wire_9720, wire_9681, wire_9680, wire_9674, wire_9641, wire_9640, wire_1417, wire_899, wire_11167, wire_9771, wire_9719, wire_9718, wire_9679, wire_9678, wire_9666, wire_9639, wire_9638, wire_1417, wire_899, wire_11165, wire_9773, wire_9717, wire_9716, wire_9677, wire_9676, wire_9658, wire_9637, wire_9636, wire_1413, wire_899, wire_11163, wire_9775, wire_9713, wire_9712, wire_9673, wire_9672, wire_9650, wire_9633, wire_9632, wire_1413, wire_899, wire_11161, wire_9777, wire_9711, wire_9710, wire_9671, wire_9670, wire_9642, wire_9631, wire_9630, wire_1413, wire_899, wire_10723, wire_10722, wire_11163, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11066, wire_9779, wire_942, wire_10739, wire_10738, wire_10709, wire_10708, wire_10693, wire_10692, wire_10799, wire_10678, wire_11165, wire_11159, wire_11158, wire_11149, wire_11148, wire_11139, wire_11138, wire_11064, wire_9777, wire_942, wire_10769, wire_10768, wire_10783, wire_10662, wire_10737, wire_10736, wire_10707, wire_10706, wire_11167, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11062, wire_9775, wire_942, wire_10753, wire_10752, wire_10797, wire_10676, wire_10767, wire_10766, wire_10735, wire_10734, wire_11169, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11060, wire_9773, wire_902, wire_10721, wire_10720, wire_10691, wire_10690, wire_10705, wire_10704, wire_10781, wire_10660, wire_11171, wire_11157, wire_11156, wire_11147, wire_11146, wire_11137, wire_11136, wire_11058, wire_9771, wire_902, wire_10751, wire_10750, wire_10795, wire_10674, wire_10719, wire_10718, wire_10689, wire_10688, wire_11173, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11056, wire_9769, wire_902, wire_10765, wire_10764, wire_10779, wire_10658, wire_10749, wire_10748, wire_10717, wire_10716, wire_11175, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11054, wire_9767, wire_946, wire_902, wire_10733, wire_10732, wire_10703, wire_10702, wire_10687, wire_10686, wire_10793, wire_10672, wire_11177, wire_11155, wire_11154, wire_11145, wire_11144, wire_11135, wire_11134, wire_11052, wire_9765, wire_946, wire_902, wire_10763, wire_10762, wire_10777, wire_10656, wire_10731, wire_10730, wire_10701, wire_10700, wire_11179, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11050, wire_9763, wire_946, wire_902, wire_10747, wire_10746, wire_10791, wire_10670, wire_10761, wire_10760, wire_10729, wire_10728, wire_946, wire_11181, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11048, wire_9761, wire_946, wire_898, wire_10715, wire_10714, wire_946, wire_10685, wire_10684, wire_946, wire_10699, wire_10698, wire_946, wire_10775, wire_10654, wire_946, wire_11183, wire_11153, wire_11152, wire_11143, wire_11142, wire_11133, wire_11132, wire_11046, wire_9759, wire_946, wire_898, wire_10745, wire_10744, wire_946, wire_10789, wire_10668, wire_942, wire_10713, wire_10712, wire_942, wire_10683, wire_10682, wire_942, wire_11185, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11044, wire_9757, wire_946, wire_898, wire_10759, wire_10758, wire_942, wire_10773, wire_10652, wire_942, wire_10743, wire_10742, wire_942, wire_10711, wire_10710, wire_902, wire_11187, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11042, wire_9755, wire_942, wire_898, wire_10727, wire_10726, wire_902, wire_10697, wire_10696, wire_902, wire_10681, wire_10680, wire_902, wire_10787, wire_10666, wire_902, wire_11189, wire_11151, wire_11150, wire_11141, wire_11140, wire_11131, wire_11130, wire_11040, wire_9753, wire_942, wire_898, wire_10757, wire_10756, wire_902, wire_10771, wire_10650, wire_898, wire_10725, wire_10724, wire_898, wire_10695, wire_10694, wire_898, wire_11161, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11068, wire_9751, wire_942, wire_898, wire_10741, wire_10740, wire_898, wire_10785, wire_10664, wire_898, wire_10755, wire_10754, wire_898};
    // CHNAXY TOTAL: 621
    assign wire_9630 = lut_tile_9_1_chanxy_out[0];
    assign wire_9632 = lut_tile_9_1_chanxy_out[1];
    assign wire_9634 = lut_tile_9_1_chanxy_out[2];
    assign wire_9635 = lut_tile_9_1_chanxy_out[3];
    assign wire_9636 = lut_tile_9_1_chanxy_out[4];
    assign wire_9638 = lut_tile_9_1_chanxy_out[5];
    assign wire_9640 = lut_tile_9_1_chanxy_out[6];
    assign wire_9642 = lut_tile_9_1_chanxy_out[7];
    assign wire_9643 = lut_tile_9_1_chanxy_out[8];
    assign wire_9644 = lut_tile_9_1_chanxy_out[9];
    assign wire_9646 = lut_tile_9_1_chanxy_out[10];
    assign wire_9648 = lut_tile_9_1_chanxy_out[11];
    assign wire_9650 = lut_tile_9_1_chanxy_out[12];
    assign wire_9651 = lut_tile_9_1_chanxy_out[13];
    assign wire_9652 = lut_tile_9_1_chanxy_out[14];
    assign wire_9654 = lut_tile_9_1_chanxy_out[15];
    assign wire_9656 = lut_tile_9_1_chanxy_out[16];
    assign wire_9658 = lut_tile_9_1_chanxy_out[17];
    assign wire_9659 = lut_tile_9_1_chanxy_out[18];
    assign wire_9660 = lut_tile_9_1_chanxy_out[19];
    assign wire_9662 = lut_tile_9_1_chanxy_out[20];
    assign wire_9664 = lut_tile_9_1_chanxy_out[21];
    assign wire_9666 = lut_tile_9_1_chanxy_out[22];
    assign wire_9667 = lut_tile_9_1_chanxy_out[23];
    assign wire_9668 = lut_tile_9_1_chanxy_out[24];
    assign wire_9670 = lut_tile_9_1_chanxy_out[25];
    assign wire_9672 = lut_tile_9_1_chanxy_out[26];
    assign wire_9674 = lut_tile_9_1_chanxy_out[27];
    assign wire_9675 = lut_tile_9_1_chanxy_out[28];
    assign wire_9676 = lut_tile_9_1_chanxy_out[29];
    assign wire_9678 = lut_tile_9_1_chanxy_out[30];
    assign wire_9680 = lut_tile_9_1_chanxy_out[31];
    assign wire_9682 = lut_tile_9_1_chanxy_out[32];
    assign wire_9683 = lut_tile_9_1_chanxy_out[33];
    assign wire_9684 = lut_tile_9_1_chanxy_out[34];
    assign wire_9686 = lut_tile_9_1_chanxy_out[35];
    assign wire_9688 = lut_tile_9_1_chanxy_out[36];
    assign wire_9690 = lut_tile_9_1_chanxy_out[37];
    assign wire_9691 = lut_tile_9_1_chanxy_out[38];
    assign wire_9692 = lut_tile_9_1_chanxy_out[39];
    assign wire_9694 = lut_tile_9_1_chanxy_out[40];
    assign wire_9696 = lut_tile_9_1_chanxy_out[41];
    assign wire_9698 = lut_tile_9_1_chanxy_out[42];
    assign wire_9699 = lut_tile_9_1_chanxy_out[43];
    assign wire_9700 = lut_tile_9_1_chanxy_out[44];
    assign wire_9702 = lut_tile_9_1_chanxy_out[45];
    assign wire_9704 = lut_tile_9_1_chanxy_out[46];
    assign wire_9706 = lut_tile_9_1_chanxy_out[47];
    assign wire_9707 = lut_tile_9_1_chanxy_out[48];
    assign wire_9708 = lut_tile_9_1_chanxy_out[49];
    assign wire_9710 = lut_tile_9_1_chanxy_out[50];
    assign wire_9712 = lut_tile_9_1_chanxy_out[51];
    assign wire_9714 = lut_tile_9_1_chanxy_out[52];
    assign wire_9715 = lut_tile_9_1_chanxy_out[53];
    assign wire_9716 = lut_tile_9_1_chanxy_out[54];
    assign wire_9718 = lut_tile_9_1_chanxy_out[55];
    assign wire_9720 = lut_tile_9_1_chanxy_out[56];
    assign wire_9722 = lut_tile_9_1_chanxy_out[57];
    assign wire_9723 = lut_tile_9_1_chanxy_out[58];
    assign wire_9724 = lut_tile_9_1_chanxy_out[59];
    assign wire_9726 = lut_tile_9_1_chanxy_out[60];
    assign wire_9728 = lut_tile_9_1_chanxy_out[61];
    assign wire_9730 = lut_tile_9_1_chanxy_out[62];
    assign wire_9731 = lut_tile_9_1_chanxy_out[63];
    assign wire_9732 = lut_tile_9_1_chanxy_out[64];
    assign wire_9734 = lut_tile_9_1_chanxy_out[65];
    assign wire_9736 = lut_tile_9_1_chanxy_out[66];
    assign wire_9738 = lut_tile_9_1_chanxy_out[67];
    assign wire_9739 = lut_tile_9_1_chanxy_out[68];
    assign wire_9740 = lut_tile_9_1_chanxy_out[69];
    assign wire_9742 = lut_tile_9_1_chanxy_out[70];
    assign wire_9744 = lut_tile_9_1_chanxy_out[71];
    assign wire_9746 = lut_tile_9_1_chanxy_out[72];
    assign wire_9747 = lut_tile_9_1_chanxy_out[73];
    assign wire_9748 = lut_tile_9_1_chanxy_out[74];
    assign wire_11041 = lut_tile_9_1_chanxy_out[75];
    assign wire_11043 = lut_tile_9_1_chanxy_out[76];
    assign wire_11045 = lut_tile_9_1_chanxy_out[77];
    assign wire_11047 = lut_tile_9_1_chanxy_out[78];
    assign wire_11049 = lut_tile_9_1_chanxy_out[79];
    assign wire_11051 = lut_tile_9_1_chanxy_out[80];
    assign wire_11053 = lut_tile_9_1_chanxy_out[81];
    assign wire_11055 = lut_tile_9_1_chanxy_out[82];
    assign wire_11057 = lut_tile_9_1_chanxy_out[83];
    assign wire_11059 = lut_tile_9_1_chanxy_out[84];
    assign wire_11061 = lut_tile_9_1_chanxy_out[85];
    assign wire_11063 = lut_tile_9_1_chanxy_out[86];
    assign wire_11065 = lut_tile_9_1_chanxy_out[87];
    assign wire_11067 = lut_tile_9_1_chanxy_out[88];
    assign wire_11069 = lut_tile_9_1_chanxy_out[89];
    assign wire_11130 = lut_tile_9_1_chanxy_out[90];
    assign wire_11132 = lut_tile_9_1_chanxy_out[91];
    assign wire_11134 = lut_tile_9_1_chanxy_out[92];
    assign wire_11136 = lut_tile_9_1_chanxy_out[93];
    assign wire_11138 = lut_tile_9_1_chanxy_out[94];
    assign wire_11140 = lut_tile_9_1_chanxy_out[95];
    assign wire_11142 = lut_tile_9_1_chanxy_out[96];
    assign wire_11144 = lut_tile_9_1_chanxy_out[97];
    assign wire_11146 = lut_tile_9_1_chanxy_out[98];
    assign wire_11148 = lut_tile_9_1_chanxy_out[99];
    assign wire_11150 = lut_tile_9_1_chanxy_out[100];
    assign wire_11152 = lut_tile_9_1_chanxy_out[101];
    assign wire_11154 = lut_tile_9_1_chanxy_out[102];
    assign wire_11156 = lut_tile_9_1_chanxy_out[103];
    assign wire_11158 = lut_tile_9_1_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_9_2_chanxy_in = {wire_11428, wire_9391, wire_9359, wire_9358, wire_9319, wire_9318, wire_9279, wire_9278, wire_9252, wire_1929, wire_11426, wire_9419, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9260, wire_1929, wire_11424, wire_9417, wire_9353, wire_9352, wire_9313, wire_9312, wire_9273, wire_9272, wire_9268, wire_1929, wire_11422, wire_9415, wire_9351, wire_9350, wire_9311, wire_9310, wire_9276, wire_9271, wire_9270, wire_1419, wire_11420, wire_9413, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9284, wire_1419, wire_11418, wire_9411, wire_9345, wire_9344, wire_9305, wire_9304, wire_9292, wire_9265, wire_9264, wire_1419, wire_11416, wire_9409, wire_9343, wire_9342, wire_9303, wire_9302, wire_9300, wire_9263, wire_9262, wire_1933, wire_1419, wire_11414, wire_9407, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9308, wire_1933, wire_1419, wire_11412, wire_9405, wire_9337, wire_9336, wire_9316, wire_9297, wire_9296, wire_9257, wire_9256, wire_1933, wire_1419, wire_11410, wire_9403, wire_9335, wire_9334, wire_9324, wire_9295, wire_9294, wire_9255, wire_9254, wire_1933, wire_1415, wire_11408, wire_9401, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9332, wire_1933, wire_1415, wire_11406, wire_9399, wire_9340, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_1933, wire_1415, wire_11404, wire_9397, wire_9348, wire_9327, wire_9326, wire_9287, wire_9286, wire_9247, wire_9246, wire_1929, wire_1415, wire_11402, wire_9395, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9356, wire_1929, wire_1415, wire_11400, wire_9393, wire_9321, wire_9320, wire_9281, wire_9280, wire_9244, wire_9241, wire_9240, wire_1929, wire_1415, wire_11579, wire_9809, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9636, wire_1929, wire_11577, wire_9781, wire_9748, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_1929, wire_11575, wire_9783, wire_9743, wire_9742, wire_9740, wire_9703, wire_9702, wire_9663, wire_9662, wire_1929, wire_11573, wire_9785, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9732, wire_1419, wire_11571, wire_9787, wire_9737, wire_9736, wire_9724, wire_9697, wire_9696, wire_9657, wire_9656, wire_1419, wire_11569, wire_9789, wire_9735, wire_9734, wire_9716, wire_9695, wire_9694, wire_9655, wire_9654, wire_1419, wire_11567, wire_9791, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9708, wire_1933, wire_1419, wire_11565, wire_9793, wire_9729, wire_9728, wire_9700, wire_9689, wire_9688, wire_9649, wire_9648, wire_1933, wire_1419, wire_11563, wire_9795, wire_9727, wire_9726, wire_9692, wire_9687, wire_9686, wire_9647, wire_9646, wire_1933, wire_1419, wire_11561, wire_9797, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9684, wire_1933, wire_1415, wire_11559, wire_9799, wire_9721, wire_9720, wire_9681, wire_9680, wire_9676, wire_9641, wire_9640, wire_1933, wire_1415, wire_11557, wire_9801, wire_9719, wire_9718, wire_9679, wire_9678, wire_9668, wire_9639, wire_9638, wire_1933, wire_1415, wire_11555, wire_9803, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9660, wire_1929, wire_1415, wire_11553, wire_9805, wire_9713, wire_9712, wire_9673, wire_9672, wire_9652, wire_9633, wire_9632, wire_1929, wire_1415, wire_11551, wire_9807, wire_9711, wire_9710, wire_9671, wire_9670, wire_9644, wire_9631, wire_9630, wire_1929, wire_1415, wire_11187, wire_11099, wire_11098, wire_11089, wire_11088, wire_11079, wire_11078, wire_11068, wire_9746, wire_1458, wire_11185, wire_11159, wire_11158, wire_11149, wire_11148, wire_11139, wire_11138, wire_11040, wire_9738, wire_1458, wire_11183, wire_11129, wire_11128, wire_11119, wire_11118, wire_11109, wire_11108, wire_11042, wire_9730, wire_1458, wire_11181, wire_11097, wire_11096, wire_11087, wire_11086, wire_11077, wire_11076, wire_11044, wire_9722, wire_1418, wire_11179, wire_11157, wire_11156, wire_11147, wire_11146, wire_11137, wire_11136, wire_11046, wire_9714, wire_1418, wire_11177, wire_11127, wire_11126, wire_11117, wire_11116, wire_11107, wire_11106, wire_11048, wire_9706, wire_1418, wire_11175, wire_11095, wire_11094, wire_11085, wire_11084, wire_11075, wire_11074, wire_11050, wire_9698, wire_1462, wire_1418, wire_11173, wire_11155, wire_11154, wire_11145, wire_11144, wire_11135, wire_11134, wire_11052, wire_9690, wire_1462, wire_1418, wire_11171, wire_11125, wire_11124, wire_11115, wire_11114, wire_11105, wire_11104, wire_11054, wire_9682, wire_1462, wire_1418, wire_11169, wire_11093, wire_11092, wire_11083, wire_11082, wire_11073, wire_11072, wire_11056, wire_9674, wire_1462, wire_1414, wire_11167, wire_11153, wire_11152, wire_11143, wire_11142, wire_11133, wire_11132, wire_11058, wire_9666, wire_1462, wire_1414, wire_11165, wire_11123, wire_11122, wire_11113, wire_11112, wire_11103, wire_11102, wire_11060, wire_9658, wire_1462, wire_1414, wire_11163, wire_11091, wire_11090, wire_11081, wire_11080, wire_11071, wire_11070, wire_11062, wire_9650, wire_1458, wire_1414, wire_11161, wire_11151, wire_11150, wire_11141, wire_11140, wire_11131, wire_11130, wire_11064, wire_9642, wire_1458, wire_1414, wire_11189, wire_11121, wire_11120, wire_11111, wire_11110, wire_11101, wire_11100, wire_11066, wire_9634, wire_1458, wire_1414, wire_11553, wire_11549, wire_11548, wire_11539, wire_11538, wire_11529, wire_11528, wire_11456, wire_9809, wire_1458, wire_11555, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11454, wire_9807, wire_1458, wire_11557, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11452, wire_9805, wire_1458, wire_11559, wire_11547, wire_11546, wire_11537, wire_11536, wire_11527, wire_11526, wire_11450, wire_9803, wire_1418, wire_11561, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11448, wire_9801, wire_1418, wire_11563, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11446, wire_9799, wire_1418, wire_11565, wire_11545, wire_11544, wire_11535, wire_11534, wire_11525, wire_11524, wire_11444, wire_9797, wire_1462, wire_1418, wire_11567, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11442, wire_9795, wire_1462, wire_1418, wire_11569, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11440, wire_9793, wire_1462, wire_1418, wire_11571, wire_11543, wire_11542, wire_11533, wire_11532, wire_11523, wire_11522, wire_11438, wire_9791, wire_1462, wire_1414, wire_11573, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11436, wire_9789, wire_1462, wire_1414, wire_11575, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11434, wire_9787, wire_1462, wire_1414, wire_11577, wire_11541, wire_11540, wire_11531, wire_11530, wire_11521, wire_11520, wire_11432, wire_9785, wire_1458, wire_1414, wire_11579, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11430, wire_9783, wire_1458, wire_1414, wire_11551, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11458, wire_9781, wire_1458, wire_1414};
    // CHNAXY TOTAL: 636
    assign wire_9637 = lut_tile_9_2_chanxy_out[0];
    assign wire_9645 = lut_tile_9_2_chanxy_out[1];
    assign wire_9653 = lut_tile_9_2_chanxy_out[2];
    assign wire_9661 = lut_tile_9_2_chanxy_out[3];
    assign wire_9669 = lut_tile_9_2_chanxy_out[4];
    assign wire_9677 = lut_tile_9_2_chanxy_out[5];
    assign wire_9685 = lut_tile_9_2_chanxy_out[6];
    assign wire_9693 = lut_tile_9_2_chanxy_out[7];
    assign wire_9701 = lut_tile_9_2_chanxy_out[8];
    assign wire_9709 = lut_tile_9_2_chanxy_out[9];
    assign wire_9717 = lut_tile_9_2_chanxy_out[10];
    assign wire_9725 = lut_tile_9_2_chanxy_out[11];
    assign wire_9733 = lut_tile_9_2_chanxy_out[12];
    assign wire_9741 = lut_tile_9_2_chanxy_out[13];
    assign wire_9749 = lut_tile_9_2_chanxy_out[14];
    assign wire_9750 = lut_tile_9_2_chanxy_out[15];
    assign wire_9752 = lut_tile_9_2_chanxy_out[16];
    assign wire_9754 = lut_tile_9_2_chanxy_out[17];
    assign wire_9756 = lut_tile_9_2_chanxy_out[18];
    assign wire_9758 = lut_tile_9_2_chanxy_out[19];
    assign wire_9760 = lut_tile_9_2_chanxy_out[20];
    assign wire_9762 = lut_tile_9_2_chanxy_out[21];
    assign wire_9764 = lut_tile_9_2_chanxy_out[22];
    assign wire_9766 = lut_tile_9_2_chanxy_out[23];
    assign wire_9768 = lut_tile_9_2_chanxy_out[24];
    assign wire_9770 = lut_tile_9_2_chanxy_out[25];
    assign wire_9772 = lut_tile_9_2_chanxy_out[26];
    assign wire_9774 = lut_tile_9_2_chanxy_out[27];
    assign wire_9776 = lut_tile_9_2_chanxy_out[28];
    assign wire_9778 = lut_tile_9_2_chanxy_out[29];
    assign wire_11431 = lut_tile_9_2_chanxy_out[30];
    assign wire_11433 = lut_tile_9_2_chanxy_out[31];
    assign wire_11435 = lut_tile_9_2_chanxy_out[32];
    assign wire_11437 = lut_tile_9_2_chanxy_out[33];
    assign wire_11439 = lut_tile_9_2_chanxy_out[34];
    assign wire_11441 = lut_tile_9_2_chanxy_out[35];
    assign wire_11443 = lut_tile_9_2_chanxy_out[36];
    assign wire_11445 = lut_tile_9_2_chanxy_out[37];
    assign wire_11447 = lut_tile_9_2_chanxy_out[38];
    assign wire_11449 = lut_tile_9_2_chanxy_out[39];
    assign wire_11451 = lut_tile_9_2_chanxy_out[40];
    assign wire_11453 = lut_tile_9_2_chanxy_out[41];
    assign wire_11455 = lut_tile_9_2_chanxy_out[42];
    assign wire_11457 = lut_tile_9_2_chanxy_out[43];
    assign wire_11459 = lut_tile_9_2_chanxy_out[44];
    assign wire_11520 = lut_tile_9_2_chanxy_out[45];
    assign wire_11522 = lut_tile_9_2_chanxy_out[46];
    assign wire_11524 = lut_tile_9_2_chanxy_out[47];
    assign wire_11526 = lut_tile_9_2_chanxy_out[48];
    assign wire_11528 = lut_tile_9_2_chanxy_out[49];
    assign wire_11530 = lut_tile_9_2_chanxy_out[50];
    assign wire_11532 = lut_tile_9_2_chanxy_out[51];
    assign wire_11534 = lut_tile_9_2_chanxy_out[52];
    assign wire_11536 = lut_tile_9_2_chanxy_out[53];
    assign wire_11538 = lut_tile_9_2_chanxy_out[54];
    assign wire_11540 = lut_tile_9_2_chanxy_out[55];
    assign wire_11542 = lut_tile_9_2_chanxy_out[56];
    assign wire_11544 = lut_tile_9_2_chanxy_out[57];
    assign wire_11546 = lut_tile_9_2_chanxy_out[58];
    assign wire_11548 = lut_tile_9_2_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_3_chanxy_in = {wire_11818, wire_9421, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9254, wire_2445, wire_11816, wire_9449, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9262, wire_2445, wire_11814, wire_9447, wire_9353, wire_9352, wire_9313, wire_9312, wire_9273, wire_9272, wire_9270, wire_2445, wire_11812, wire_9445, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9278, wire_1935, wire_11810, wire_9443, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9286, wire_1935, wire_11808, wire_9441, wire_9345, wire_9344, wire_9305, wire_9304, wire_9294, wire_9265, wire_9264, wire_1935, wire_11806, wire_9439, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9302, wire_2449, wire_1935, wire_11804, wire_9437, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9310, wire_2449, wire_1935, wire_11802, wire_9435, wire_9337, wire_9336, wire_9318, wire_9297, wire_9296, wire_9257, wire_9256, wire_2449, wire_1935, wire_11800, wire_9433, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9326, wire_2449, wire_1931, wire_11798, wire_9431, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9334, wire_2449, wire_1931, wire_11796, wire_9429, wire_9342, wire_9329, wire_9328, wire_9289, wire_9288, wire_9249, wire_9248, wire_2449, wire_1931, wire_11794, wire_9427, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9350, wire_2445, wire_1931, wire_11792, wire_9425, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9358, wire_2445, wire_1931, wire_11790, wire_9423, wire_9321, wire_9320, wire_9281, wire_9280, wire_9246, wire_9241, wire_9240, wire_2445, wire_1931, wire_11969, wire_9839, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9630, wire_2445, wire_11967, wire_9811, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9742, wire_2445, wire_11965, wire_9813, wire_9745, wire_9744, wire_9734, wire_9705, wire_9704, wire_9665, wire_9664, wire_2445, wire_11963, wire_9815, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9726, wire_1935, wire_11961, wire_9817, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9718, wire_1935, wire_11959, wire_9819, wire_9737, wire_9736, wire_9710, wire_9697, wire_9696, wire_9657, wire_9656, wire_1935, wire_11957, wire_9821, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9702, wire_2449, wire_1935, wire_11955, wire_9823, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9694, wire_2449, wire_1935, wire_11953, wire_9825, wire_9729, wire_9728, wire_9689, wire_9688, wire_9686, wire_9649, wire_9648, wire_2449, wire_1935, wire_11951, wire_9827, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9678, wire_2449, wire_1931, wire_11949, wire_9829, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9670, wire_2449, wire_1931, wire_11947, wire_9831, wire_9721, wire_9720, wire_9681, wire_9680, wire_9662, wire_9641, wire_9640, wire_2449, wire_1931, wire_11945, wire_9833, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9654, wire_2445, wire_1931, wire_11943, wire_9835, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9646, wire_2445, wire_1931, wire_11941, wire_9837, wire_9713, wire_9712, wire_9673, wire_9672, wire_9638, wire_9633, wire_9632, wire_2445, wire_1931, wire_11577, wire_11549, wire_11548, wire_11539, wire_11538, wire_11529, wire_11528, wire_11458, wire_9748, wire_1974, wire_11575, wire_11519, wire_11518, wire_11509, wire_11508, wire_11499, wire_11498, wire_11430, wire_9740, wire_1974, wire_11573, wire_11489, wire_11488, wire_11479, wire_11478, wire_11469, wire_11468, wire_11432, wire_9732, wire_1974, wire_11571, wire_11547, wire_11546, wire_11537, wire_11536, wire_11527, wire_11526, wire_11434, wire_9724, wire_1934, wire_11569, wire_11517, wire_11516, wire_11507, wire_11506, wire_11497, wire_11496, wire_11436, wire_9716, wire_1934, wire_11567, wire_11487, wire_11486, wire_11477, wire_11476, wire_11467, wire_11466, wire_11438, wire_9708, wire_1934, wire_11565, wire_11545, wire_11544, wire_11535, wire_11534, wire_11525, wire_11524, wire_11440, wire_9700, wire_1978, wire_1934, wire_11563, wire_11515, wire_11514, wire_11505, wire_11504, wire_11495, wire_11494, wire_11442, wire_9692, wire_1978, wire_1934, wire_11561, wire_11485, wire_11484, wire_11475, wire_11474, wire_11465, wire_11464, wire_11444, wire_9684, wire_1978, wire_1934, wire_11559, wire_11543, wire_11542, wire_11533, wire_11532, wire_11523, wire_11522, wire_11446, wire_9676, wire_1978, wire_1930, wire_11557, wire_11513, wire_11512, wire_11503, wire_11502, wire_11493, wire_11492, wire_11448, wire_9668, wire_1978, wire_1930, wire_11555, wire_11483, wire_11482, wire_11473, wire_11472, wire_11463, wire_11462, wire_11450, wire_9660, wire_1978, wire_1930, wire_11553, wire_11541, wire_11540, wire_11531, wire_11530, wire_11521, wire_11520, wire_11452, wire_9652, wire_1974, wire_1930, wire_11551, wire_11511, wire_11510, wire_11501, wire_11500, wire_11491, wire_11490, wire_11454, wire_9644, wire_1974, wire_1930, wire_11579, wire_11481, wire_11480, wire_11471, wire_11470, wire_11461, wire_11460, wire_11456, wire_9636, wire_1974, wire_1930, wire_11943, wire_11939, wire_11938, wire_11929, wire_11928, wire_11919, wire_11918, wire_11846, wire_9839, wire_1974, wire_11945, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11844, wire_9837, wire_1974, wire_11947, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11842, wire_9835, wire_1974, wire_11949, wire_11937, wire_11936, wire_11927, wire_11926, wire_11917, wire_11916, wire_11840, wire_9833, wire_1934, wire_11951, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11838, wire_9831, wire_1934, wire_11953, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11836, wire_9829, wire_1934, wire_11955, wire_11935, wire_11934, wire_11925, wire_11924, wire_11915, wire_11914, wire_11834, wire_9827, wire_1978, wire_1934, wire_11957, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11832, wire_9825, wire_1978, wire_1934, wire_11959, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11830, wire_9823, wire_1978, wire_1934, wire_11961, wire_11933, wire_11932, wire_11923, wire_11922, wire_11913, wire_11912, wire_11828, wire_9821, wire_1978, wire_1930, wire_11963, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11826, wire_9819, wire_1978, wire_1930, wire_11965, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11824, wire_9817, wire_1978, wire_1930, wire_11967, wire_11931, wire_11930, wire_11921, wire_11920, wire_11911, wire_11910, wire_11822, wire_9815, wire_1974, wire_1930, wire_11969, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11820, wire_9813, wire_1974, wire_1930, wire_11941, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11848, wire_9811, wire_1974, wire_1930};
    // CHNAXY TOTAL: 636
    assign wire_9631 = lut_tile_9_3_chanxy_out[0];
    assign wire_9639 = lut_tile_9_3_chanxy_out[1];
    assign wire_9647 = lut_tile_9_3_chanxy_out[2];
    assign wire_9655 = lut_tile_9_3_chanxy_out[3];
    assign wire_9663 = lut_tile_9_3_chanxy_out[4];
    assign wire_9671 = lut_tile_9_3_chanxy_out[5];
    assign wire_9679 = lut_tile_9_3_chanxy_out[6];
    assign wire_9687 = lut_tile_9_3_chanxy_out[7];
    assign wire_9695 = lut_tile_9_3_chanxy_out[8];
    assign wire_9703 = lut_tile_9_3_chanxy_out[9];
    assign wire_9711 = lut_tile_9_3_chanxy_out[10];
    assign wire_9719 = lut_tile_9_3_chanxy_out[11];
    assign wire_9727 = lut_tile_9_3_chanxy_out[12];
    assign wire_9735 = lut_tile_9_3_chanxy_out[13];
    assign wire_9743 = lut_tile_9_3_chanxy_out[14];
    assign wire_9780 = lut_tile_9_3_chanxy_out[15];
    assign wire_9782 = lut_tile_9_3_chanxy_out[16];
    assign wire_9784 = lut_tile_9_3_chanxy_out[17];
    assign wire_9786 = lut_tile_9_3_chanxy_out[18];
    assign wire_9788 = lut_tile_9_3_chanxy_out[19];
    assign wire_9790 = lut_tile_9_3_chanxy_out[20];
    assign wire_9792 = lut_tile_9_3_chanxy_out[21];
    assign wire_9794 = lut_tile_9_3_chanxy_out[22];
    assign wire_9796 = lut_tile_9_3_chanxy_out[23];
    assign wire_9798 = lut_tile_9_3_chanxy_out[24];
    assign wire_9800 = lut_tile_9_3_chanxy_out[25];
    assign wire_9802 = lut_tile_9_3_chanxy_out[26];
    assign wire_9804 = lut_tile_9_3_chanxy_out[27];
    assign wire_9806 = lut_tile_9_3_chanxy_out[28];
    assign wire_9808 = lut_tile_9_3_chanxy_out[29];
    assign wire_11821 = lut_tile_9_3_chanxy_out[30];
    assign wire_11823 = lut_tile_9_3_chanxy_out[31];
    assign wire_11825 = lut_tile_9_3_chanxy_out[32];
    assign wire_11827 = lut_tile_9_3_chanxy_out[33];
    assign wire_11829 = lut_tile_9_3_chanxy_out[34];
    assign wire_11831 = lut_tile_9_3_chanxy_out[35];
    assign wire_11833 = lut_tile_9_3_chanxy_out[36];
    assign wire_11835 = lut_tile_9_3_chanxy_out[37];
    assign wire_11837 = lut_tile_9_3_chanxy_out[38];
    assign wire_11839 = lut_tile_9_3_chanxy_out[39];
    assign wire_11841 = lut_tile_9_3_chanxy_out[40];
    assign wire_11843 = lut_tile_9_3_chanxy_out[41];
    assign wire_11845 = lut_tile_9_3_chanxy_out[42];
    assign wire_11847 = lut_tile_9_3_chanxy_out[43];
    assign wire_11849 = lut_tile_9_3_chanxy_out[44];
    assign wire_11910 = lut_tile_9_3_chanxy_out[45];
    assign wire_11912 = lut_tile_9_3_chanxy_out[46];
    assign wire_11914 = lut_tile_9_3_chanxy_out[47];
    assign wire_11916 = lut_tile_9_3_chanxy_out[48];
    assign wire_11918 = lut_tile_9_3_chanxy_out[49];
    assign wire_11920 = lut_tile_9_3_chanxy_out[50];
    assign wire_11922 = lut_tile_9_3_chanxy_out[51];
    assign wire_11924 = lut_tile_9_3_chanxy_out[52];
    assign wire_11926 = lut_tile_9_3_chanxy_out[53];
    assign wire_11928 = lut_tile_9_3_chanxy_out[54];
    assign wire_11930 = lut_tile_9_3_chanxy_out[55];
    assign wire_11932 = lut_tile_9_3_chanxy_out[56];
    assign wire_11934 = lut_tile_9_3_chanxy_out[57];
    assign wire_11936 = lut_tile_9_3_chanxy_out[58];
    assign wire_11938 = lut_tile_9_3_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_4_chanxy_in = {wire_12208, wire_9451, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9248, wire_2961, wire_12206, wire_9479, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9256, wire_2961, wire_12204, wire_9477, wire_9389, wire_9388, wire_9379, wire_9378, wire_9369, wire_9368, wire_9264, wire_2961, wire_12202, wire_9475, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9272, wire_2451, wire_12200, wire_9473, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9280, wire_2451, wire_12198, wire_9471, wire_9387, wire_9386, wire_9377, wire_9376, wire_9367, wire_9366, wire_9288, wire_2451, wire_12196, wire_9469, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9296, wire_2965, wire_2451, wire_12194, wire_9467, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9304, wire_2965, wire_2451, wire_12192, wire_9465, wire_9385, wire_9384, wire_9375, wire_9374, wire_9365, wire_9364, wire_9312, wire_2965, wire_2451, wire_12190, wire_9463, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9320, wire_2965, wire_2447, wire_12188, wire_9461, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9328, wire_2965, wire_2447, wire_12186, wire_9459, wire_9383, wire_9382, wire_9373, wire_9372, wire_9363, wire_9362, wire_9336, wire_2965, wire_2447, wire_12184, wire_9457, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9344, wire_2961, wire_2447, wire_12182, wire_9455, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9352, wire_2961, wire_2447, wire_12180, wire_9453, wire_9381, wire_9380, wire_9371, wire_9370, wire_9361, wire_9360, wire_9240, wire_2961, wire_2447, wire_12359, wire_9869, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9632, wire_2961, wire_12357, wire_9841, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9744, wire_2961, wire_12355, wire_9843, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9736, wire_2961, wire_12353, wire_9845, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9728, wire_2451, wire_12351, wire_9847, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9720, wire_2451, wire_12349, wire_9849, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9712, wire_2451, wire_12347, wire_9851, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9704, wire_2965, wire_2451, wire_12345, wire_9853, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9696, wire_2965, wire_2451, wire_12343, wire_9855, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9688, wire_2965, wire_2451, wire_12341, wire_9857, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9680, wire_2965, wire_2447, wire_12339, wire_9859, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9672, wire_2965, wire_2447, wire_12337, wire_9861, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9664, wire_2965, wire_2447, wire_12335, wire_9863, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9656, wire_2961, wire_2447, wire_12333, wire_9865, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9648, wire_2961, wire_2447, wire_12331, wire_9867, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9640, wire_2961, wire_2447, wire_11967, wire_11939, wire_11938, wire_11929, wire_11928, wire_11919, wire_11918, wire_11848, wire_9742, wire_2490, wire_11965, wire_11909, wire_11908, wire_11899, wire_11898, wire_11889, wire_11888, wire_11820, wire_9734, wire_2490, wire_11963, wire_11879, wire_11878, wire_11869, wire_11868, wire_11859, wire_11858, wire_11822, wire_9726, wire_2490, wire_11961, wire_11937, wire_11936, wire_11927, wire_11926, wire_11917, wire_11916, wire_11824, wire_9718, wire_2450, wire_11959, wire_11907, wire_11906, wire_11897, wire_11896, wire_11887, wire_11886, wire_11826, wire_9710, wire_2450, wire_11957, wire_11877, wire_11876, wire_11867, wire_11866, wire_11857, wire_11856, wire_11828, wire_9702, wire_2450, wire_11955, wire_11935, wire_11934, wire_11925, wire_11924, wire_11915, wire_11914, wire_11830, wire_9694, wire_2494, wire_2450, wire_11953, wire_11905, wire_11904, wire_11895, wire_11894, wire_11885, wire_11884, wire_11832, wire_9686, wire_2494, wire_2450, wire_11951, wire_11875, wire_11874, wire_11865, wire_11864, wire_11855, wire_11854, wire_11834, wire_9678, wire_2494, wire_2450, wire_11949, wire_11933, wire_11932, wire_11923, wire_11922, wire_11913, wire_11912, wire_11836, wire_9670, wire_2494, wire_2446, wire_11947, wire_11903, wire_11902, wire_11893, wire_11892, wire_11883, wire_11882, wire_11838, wire_9662, wire_2494, wire_2446, wire_11945, wire_11873, wire_11872, wire_11863, wire_11862, wire_11853, wire_11852, wire_11840, wire_9654, wire_2494, wire_2446, wire_11943, wire_11931, wire_11930, wire_11921, wire_11920, wire_11911, wire_11910, wire_11842, wire_9646, wire_2490, wire_2446, wire_11941, wire_11901, wire_11900, wire_11891, wire_11890, wire_11881, wire_11880, wire_11844, wire_9638, wire_2490, wire_2446, wire_11969, wire_11871, wire_11870, wire_11861, wire_11860, wire_11851, wire_11850, wire_11846, wire_9630, wire_2490, wire_2446, wire_12333, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12236, wire_9869, wire_2490, wire_12335, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12234, wire_9867, wire_2490, wire_12337, wire_12329, wire_12328, wire_12319, wire_12318, wire_12309, wire_12308, wire_12232, wire_9865, wire_2490, wire_12339, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12230, wire_9863, wire_2450, wire_12341, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12228, wire_9861, wire_2450, wire_12343, wire_12327, wire_12326, wire_12317, wire_12316, wire_12307, wire_12306, wire_12226, wire_9859, wire_2450, wire_12345, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12224, wire_9857, wire_2494, wire_2450, wire_12347, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12222, wire_9855, wire_2494, wire_2450, wire_12349, wire_12325, wire_12324, wire_12315, wire_12314, wire_12305, wire_12304, wire_12220, wire_9853, wire_2494, wire_2450, wire_12351, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12218, wire_9851, wire_2494, wire_2446, wire_12353, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12216, wire_9849, wire_2494, wire_2446, wire_12355, wire_12323, wire_12322, wire_12313, wire_12312, wire_12303, wire_12302, wire_12214, wire_9847, wire_2494, wire_2446, wire_12357, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12212, wire_9845, wire_2490, wire_2446, wire_12359, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12210, wire_9843, wire_2490, wire_2446, wire_12331, wire_12321, wire_12320, wire_12311, wire_12310, wire_12301, wire_12300, wire_12238, wire_9841, wire_2490, wire_2446};
    // CHNAXY TOTAL: 636
    assign wire_9633 = lut_tile_9_4_chanxy_out[0];
    assign wire_9641 = lut_tile_9_4_chanxy_out[1];
    assign wire_9649 = lut_tile_9_4_chanxy_out[2];
    assign wire_9657 = lut_tile_9_4_chanxy_out[3];
    assign wire_9665 = lut_tile_9_4_chanxy_out[4];
    assign wire_9673 = lut_tile_9_4_chanxy_out[5];
    assign wire_9681 = lut_tile_9_4_chanxy_out[6];
    assign wire_9689 = lut_tile_9_4_chanxy_out[7];
    assign wire_9697 = lut_tile_9_4_chanxy_out[8];
    assign wire_9705 = lut_tile_9_4_chanxy_out[9];
    assign wire_9713 = lut_tile_9_4_chanxy_out[10];
    assign wire_9721 = lut_tile_9_4_chanxy_out[11];
    assign wire_9729 = lut_tile_9_4_chanxy_out[12];
    assign wire_9737 = lut_tile_9_4_chanxy_out[13];
    assign wire_9745 = lut_tile_9_4_chanxy_out[14];
    assign wire_9810 = lut_tile_9_4_chanxy_out[15];
    assign wire_9812 = lut_tile_9_4_chanxy_out[16];
    assign wire_9814 = lut_tile_9_4_chanxy_out[17];
    assign wire_9816 = lut_tile_9_4_chanxy_out[18];
    assign wire_9818 = lut_tile_9_4_chanxy_out[19];
    assign wire_9820 = lut_tile_9_4_chanxy_out[20];
    assign wire_9822 = lut_tile_9_4_chanxy_out[21];
    assign wire_9824 = lut_tile_9_4_chanxy_out[22];
    assign wire_9826 = lut_tile_9_4_chanxy_out[23];
    assign wire_9828 = lut_tile_9_4_chanxy_out[24];
    assign wire_9830 = lut_tile_9_4_chanxy_out[25];
    assign wire_9832 = lut_tile_9_4_chanxy_out[26];
    assign wire_9834 = lut_tile_9_4_chanxy_out[27];
    assign wire_9836 = lut_tile_9_4_chanxy_out[28];
    assign wire_9838 = lut_tile_9_4_chanxy_out[29];
    assign wire_12211 = lut_tile_9_4_chanxy_out[30];
    assign wire_12213 = lut_tile_9_4_chanxy_out[31];
    assign wire_12215 = lut_tile_9_4_chanxy_out[32];
    assign wire_12217 = lut_tile_9_4_chanxy_out[33];
    assign wire_12219 = lut_tile_9_4_chanxy_out[34];
    assign wire_12221 = lut_tile_9_4_chanxy_out[35];
    assign wire_12223 = lut_tile_9_4_chanxy_out[36];
    assign wire_12225 = lut_tile_9_4_chanxy_out[37];
    assign wire_12227 = lut_tile_9_4_chanxy_out[38];
    assign wire_12229 = lut_tile_9_4_chanxy_out[39];
    assign wire_12231 = lut_tile_9_4_chanxy_out[40];
    assign wire_12233 = lut_tile_9_4_chanxy_out[41];
    assign wire_12235 = lut_tile_9_4_chanxy_out[42];
    assign wire_12237 = lut_tile_9_4_chanxy_out[43];
    assign wire_12239 = lut_tile_9_4_chanxy_out[44];
    assign wire_12300 = lut_tile_9_4_chanxy_out[45];
    assign wire_12302 = lut_tile_9_4_chanxy_out[46];
    assign wire_12304 = lut_tile_9_4_chanxy_out[47];
    assign wire_12306 = lut_tile_9_4_chanxy_out[48];
    assign wire_12308 = lut_tile_9_4_chanxy_out[49];
    assign wire_12310 = lut_tile_9_4_chanxy_out[50];
    assign wire_12312 = lut_tile_9_4_chanxy_out[51];
    assign wire_12314 = lut_tile_9_4_chanxy_out[52];
    assign wire_12316 = lut_tile_9_4_chanxy_out[53];
    assign wire_12318 = lut_tile_9_4_chanxy_out[54];
    assign wire_12320 = lut_tile_9_4_chanxy_out[55];
    assign wire_12322 = lut_tile_9_4_chanxy_out[56];
    assign wire_12324 = lut_tile_9_4_chanxy_out[57];
    assign wire_12326 = lut_tile_9_4_chanxy_out[58];
    assign wire_12328 = lut_tile_9_4_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_5_chanxy_in = {wire_12598, wire_9481, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9362, wire_3477, wire_12596, wire_9509, wire_9419, wire_9418, wire_9409, wire_9408, wire_9399, wire_9398, wire_9364, wire_3477, wire_12594, wire_9507, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9366, wire_3477, wire_12592, wire_9505, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9368, wire_2967, wire_12590, wire_9503, wire_9417, wire_9416, wire_9407, wire_9406, wire_9397, wire_9396, wire_9370, wire_2967, wire_12588, wire_9501, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9372, wire_2967, wire_12586, wire_9499, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9374, wire_3481, wire_2967, wire_12584, wire_9497, wire_9415, wire_9414, wire_9405, wire_9404, wire_9395, wire_9394, wire_9376, wire_3481, wire_2967, wire_12582, wire_9495, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9378, wire_3481, wire_2967, wire_12580, wire_9493, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9380, wire_3481, wire_2963, wire_12578, wire_9491, wire_9413, wire_9412, wire_9403, wire_9402, wire_9393, wire_9392, wire_9382, wire_3481, wire_2963, wire_12576, wire_9489, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9384, wire_3481, wire_2963, wire_12574, wire_9487, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9386, wire_3477, wire_2963, wire_12572, wire_9485, wire_9411, wire_9410, wire_9401, wire_9400, wire_9391, wire_9390, wire_9388, wire_3477, wire_2963, wire_12570, wire_9483, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9360, wire_3477, wire_2963, wire_12749, wire_9899, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9750, wire_3477, wire_12747, wire_9871, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9778, wire_3477, wire_12745, wire_9873, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9776, wire_3477, wire_12743, wire_9875, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9774, wire_2967, wire_12741, wire_9877, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9772, wire_2967, wire_12739, wire_9879, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9770, wire_2967, wire_12737, wire_9881, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9768, wire_3481, wire_2967, wire_12735, wire_9883, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9766, wire_3481, wire_2967, wire_12733, wire_9885, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9764, wire_3481, wire_2967, wire_12731, wire_9887, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9762, wire_3481, wire_2963, wire_12729, wire_9889, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9760, wire_3481, wire_2963, wire_12727, wire_9891, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9758, wire_3481, wire_2963, wire_12725, wire_9893, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9756, wire_3477, wire_2963, wire_12723, wire_9895, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9754, wire_3477, wire_2963, wire_12721, wire_9897, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9752, wire_3477, wire_2963, wire_12357, wire_12299, wire_12298, wire_12289, wire_12288, wire_12279, wire_12278, wire_12238, wire_9744, wire_3006, wire_12355, wire_12269, wire_12268, wire_12259, wire_12258, wire_12249, wire_12248, wire_12210, wire_9736, wire_3006, wire_12353, wire_12329, wire_12328, wire_12319, wire_12318, wire_12309, wire_12308, wire_12212, wire_9728, wire_3006, wire_12351, wire_12297, wire_12296, wire_12287, wire_12286, wire_12277, wire_12276, wire_12214, wire_9720, wire_2966, wire_12349, wire_12267, wire_12266, wire_12257, wire_12256, wire_12247, wire_12246, wire_12216, wire_9712, wire_2966, wire_12347, wire_12327, wire_12326, wire_12317, wire_12316, wire_12307, wire_12306, wire_12218, wire_9704, wire_2966, wire_12345, wire_12295, wire_12294, wire_12285, wire_12284, wire_12275, wire_12274, wire_12220, wire_9696, wire_3010, wire_2966, wire_12343, wire_12265, wire_12264, wire_12255, wire_12254, wire_12245, wire_12244, wire_12222, wire_9688, wire_3010, wire_2966, wire_12341, wire_12325, wire_12324, wire_12315, wire_12314, wire_12305, wire_12304, wire_12224, wire_9680, wire_3010, wire_2966, wire_12339, wire_12293, wire_12292, wire_12283, wire_12282, wire_12273, wire_12272, wire_12226, wire_9672, wire_3010, wire_2962, wire_12337, wire_12263, wire_12262, wire_12253, wire_12252, wire_12243, wire_12242, wire_12228, wire_9664, wire_3010, wire_2962, wire_12335, wire_12323, wire_12322, wire_12313, wire_12312, wire_12303, wire_12302, wire_12230, wire_9656, wire_3010, wire_2962, wire_12333, wire_12291, wire_12290, wire_12281, wire_12280, wire_12271, wire_12270, wire_12232, wire_9648, wire_3006, wire_2962, wire_12331, wire_12261, wire_12260, wire_12251, wire_12250, wire_12241, wire_12240, wire_12234, wire_9640, wire_3006, wire_2962, wire_12359, wire_12321, wire_12320, wire_12311, wire_12310, wire_12301, wire_12300, wire_12236, wire_9632, wire_3006, wire_2962, wire_12723, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12626, wire_9899, wire_3006, wire_12725, wire_12719, wire_12718, wire_12709, wire_12708, wire_12699, wire_12698, wire_12624, wire_9897, wire_3006, wire_12727, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12622, wire_9895, wire_3006, wire_12729, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12620, wire_9893, wire_2966, wire_12731, wire_12717, wire_12716, wire_12707, wire_12706, wire_12697, wire_12696, wire_12618, wire_9891, wire_2966, wire_12733, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12616, wire_9889, wire_2966, wire_12735, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12614, wire_9887, wire_3010, wire_2966, wire_12737, wire_12715, wire_12714, wire_12705, wire_12704, wire_12695, wire_12694, wire_12612, wire_9885, wire_3010, wire_2966, wire_12739, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12610, wire_9883, wire_3010, wire_2966, wire_12741, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12608, wire_9881, wire_3010, wire_2962, wire_12743, wire_12713, wire_12712, wire_12703, wire_12702, wire_12693, wire_12692, wire_12606, wire_9879, wire_3010, wire_2962, wire_12745, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12604, wire_9877, wire_3010, wire_2962, wire_12747, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12602, wire_9875, wire_3006, wire_2962, wire_12749, wire_12711, wire_12710, wire_12701, wire_12700, wire_12691, wire_12690, wire_12600, wire_9873, wire_3006, wire_2962, wire_12721, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12628, wire_9871, wire_3006, wire_2962};
    // CHNAXY TOTAL: 636
    assign wire_9751 = lut_tile_9_5_chanxy_out[0];
    assign wire_9753 = lut_tile_9_5_chanxy_out[1];
    assign wire_9755 = lut_tile_9_5_chanxy_out[2];
    assign wire_9757 = lut_tile_9_5_chanxy_out[3];
    assign wire_9759 = lut_tile_9_5_chanxy_out[4];
    assign wire_9761 = lut_tile_9_5_chanxy_out[5];
    assign wire_9763 = lut_tile_9_5_chanxy_out[6];
    assign wire_9765 = lut_tile_9_5_chanxy_out[7];
    assign wire_9767 = lut_tile_9_5_chanxy_out[8];
    assign wire_9769 = lut_tile_9_5_chanxy_out[9];
    assign wire_9771 = lut_tile_9_5_chanxy_out[10];
    assign wire_9773 = lut_tile_9_5_chanxy_out[11];
    assign wire_9775 = lut_tile_9_5_chanxy_out[12];
    assign wire_9777 = lut_tile_9_5_chanxy_out[13];
    assign wire_9779 = lut_tile_9_5_chanxy_out[14];
    assign wire_9840 = lut_tile_9_5_chanxy_out[15];
    assign wire_9842 = lut_tile_9_5_chanxy_out[16];
    assign wire_9844 = lut_tile_9_5_chanxy_out[17];
    assign wire_9846 = lut_tile_9_5_chanxy_out[18];
    assign wire_9848 = lut_tile_9_5_chanxy_out[19];
    assign wire_9850 = lut_tile_9_5_chanxy_out[20];
    assign wire_9852 = lut_tile_9_5_chanxy_out[21];
    assign wire_9854 = lut_tile_9_5_chanxy_out[22];
    assign wire_9856 = lut_tile_9_5_chanxy_out[23];
    assign wire_9858 = lut_tile_9_5_chanxy_out[24];
    assign wire_9860 = lut_tile_9_5_chanxy_out[25];
    assign wire_9862 = lut_tile_9_5_chanxy_out[26];
    assign wire_9864 = lut_tile_9_5_chanxy_out[27];
    assign wire_9866 = lut_tile_9_5_chanxy_out[28];
    assign wire_9868 = lut_tile_9_5_chanxy_out[29];
    assign wire_12601 = lut_tile_9_5_chanxy_out[30];
    assign wire_12603 = lut_tile_9_5_chanxy_out[31];
    assign wire_12605 = lut_tile_9_5_chanxy_out[32];
    assign wire_12607 = lut_tile_9_5_chanxy_out[33];
    assign wire_12609 = lut_tile_9_5_chanxy_out[34];
    assign wire_12611 = lut_tile_9_5_chanxy_out[35];
    assign wire_12613 = lut_tile_9_5_chanxy_out[36];
    assign wire_12615 = lut_tile_9_5_chanxy_out[37];
    assign wire_12617 = lut_tile_9_5_chanxy_out[38];
    assign wire_12619 = lut_tile_9_5_chanxy_out[39];
    assign wire_12621 = lut_tile_9_5_chanxy_out[40];
    assign wire_12623 = lut_tile_9_5_chanxy_out[41];
    assign wire_12625 = lut_tile_9_5_chanxy_out[42];
    assign wire_12627 = lut_tile_9_5_chanxy_out[43];
    assign wire_12629 = lut_tile_9_5_chanxy_out[44];
    assign wire_12690 = lut_tile_9_5_chanxy_out[45];
    assign wire_12692 = lut_tile_9_5_chanxy_out[46];
    assign wire_12694 = lut_tile_9_5_chanxy_out[47];
    assign wire_12696 = lut_tile_9_5_chanxy_out[48];
    assign wire_12698 = lut_tile_9_5_chanxy_out[49];
    assign wire_12700 = lut_tile_9_5_chanxy_out[50];
    assign wire_12702 = lut_tile_9_5_chanxy_out[51];
    assign wire_12704 = lut_tile_9_5_chanxy_out[52];
    assign wire_12706 = lut_tile_9_5_chanxy_out[53];
    assign wire_12708 = lut_tile_9_5_chanxy_out[54];
    assign wire_12710 = lut_tile_9_5_chanxy_out[55];
    assign wire_12712 = lut_tile_9_5_chanxy_out[56];
    assign wire_12714 = lut_tile_9_5_chanxy_out[57];
    assign wire_12716 = lut_tile_9_5_chanxy_out[58];
    assign wire_12718 = lut_tile_9_5_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_6_chanxy_in = {wire_12988, wire_9511, wire_9449, wire_9448, wire_9439, wire_9438, wire_9429, wire_9428, wire_9392, wire_3993, wire_12986, wire_9539, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9394, wire_3993, wire_12984, wire_9537, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9396, wire_3993, wire_12982, wire_9535, wire_9447, wire_9446, wire_9437, wire_9436, wire_9427, wire_9426, wire_9398, wire_3483, wire_12980, wire_9533, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9400, wire_3483, wire_12978, wire_9531, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9402, wire_3483, wire_12976, wire_9529, wire_9445, wire_9444, wire_9435, wire_9434, wire_9425, wire_9424, wire_9404, wire_3997, wire_3483, wire_12974, wire_9527, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9406, wire_3997, wire_3483, wire_12972, wire_9525, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9408, wire_3997, wire_3483, wire_12970, wire_9523, wire_9443, wire_9442, wire_9433, wire_9432, wire_9423, wire_9422, wire_9410, wire_3997, wire_3479, wire_12968, wire_9521, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9412, wire_3997, wire_3479, wire_12966, wire_9519, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9414, wire_3997, wire_3479, wire_12964, wire_9517, wire_9441, wire_9440, wire_9431, wire_9430, wire_9421, wire_9420, wire_9416, wire_3993, wire_3479, wire_12962, wire_9515, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9418, wire_3993, wire_3479, wire_12960, wire_9513, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9390, wire_3993, wire_3479, wire_13139, wire_9929, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9780, wire_3993, wire_13137, wire_9901, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9808, wire_3993, wire_13135, wire_9903, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9806, wire_3993, wire_13133, wire_9905, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9804, wire_3483, wire_13131, wire_9907, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9802, wire_3483, wire_13129, wire_9909, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9800, wire_3483, wire_13127, wire_9911, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9798, wire_3997, wire_3483, wire_13125, wire_9913, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9796, wire_3997, wire_3483, wire_13123, wire_9915, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9794, wire_3997, wire_3483, wire_13121, wire_9917, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9792, wire_3997, wire_3479, wire_13119, wire_9919, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9790, wire_3997, wire_3479, wire_13117, wire_9921, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9788, wire_3997, wire_3479, wire_13115, wire_9923, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9786, wire_3993, wire_3479, wire_13113, wire_9925, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9784, wire_3993, wire_3479, wire_13111, wire_9927, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9782, wire_3993, wire_3479, wire_12747, wire_12659, wire_12658, wire_12649, wire_12648, wire_12639, wire_12638, wire_12628, wire_9778, wire_3522, wire_12745, wire_12719, wire_12718, wire_12709, wire_12708, wire_12699, wire_12698, wire_12600, wire_9776, wire_3522, wire_12743, wire_12689, wire_12688, wire_12679, wire_12678, wire_12669, wire_12668, wire_12602, wire_9774, wire_3522, wire_12741, wire_12657, wire_12656, wire_12647, wire_12646, wire_12637, wire_12636, wire_12604, wire_9772, wire_3482, wire_12739, wire_12717, wire_12716, wire_12707, wire_12706, wire_12697, wire_12696, wire_12606, wire_9770, wire_3482, wire_12737, wire_12687, wire_12686, wire_12677, wire_12676, wire_12667, wire_12666, wire_12608, wire_9768, wire_3482, wire_12735, wire_12655, wire_12654, wire_12645, wire_12644, wire_12635, wire_12634, wire_12610, wire_9766, wire_3526, wire_3482, wire_12733, wire_12715, wire_12714, wire_12705, wire_12704, wire_12695, wire_12694, wire_12612, wire_9764, wire_3526, wire_3482, wire_12731, wire_12685, wire_12684, wire_12675, wire_12674, wire_12665, wire_12664, wire_12614, wire_9762, wire_3526, wire_3482, wire_12729, wire_12653, wire_12652, wire_12643, wire_12642, wire_12633, wire_12632, wire_12616, wire_9760, wire_3526, wire_3478, wire_12727, wire_12713, wire_12712, wire_12703, wire_12702, wire_12693, wire_12692, wire_12618, wire_9758, wire_3526, wire_3478, wire_12725, wire_12683, wire_12682, wire_12673, wire_12672, wire_12663, wire_12662, wire_12620, wire_9756, wire_3526, wire_3478, wire_12723, wire_12651, wire_12650, wire_12641, wire_12640, wire_12631, wire_12630, wire_12622, wire_9754, wire_3522, wire_3478, wire_12721, wire_12711, wire_12710, wire_12701, wire_12700, wire_12691, wire_12690, wire_12624, wire_9752, wire_3522, wire_3478, wire_12749, wire_12681, wire_12680, wire_12671, wire_12670, wire_12661, wire_12660, wire_12626, wire_9750, wire_3522, wire_3478, wire_13113, wire_13109, wire_13108, wire_13099, wire_13098, wire_13089, wire_13088, wire_13016, wire_9929, wire_3522, wire_13115, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_13014, wire_9927, wire_3522, wire_13117, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_13012, wire_9925, wire_3522, wire_13119, wire_13107, wire_13106, wire_13097, wire_13096, wire_13087, wire_13086, wire_13010, wire_9923, wire_3482, wire_13121, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_13008, wire_9921, wire_3482, wire_13123, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_13006, wire_9919, wire_3482, wire_13125, wire_13105, wire_13104, wire_13095, wire_13094, wire_13085, wire_13084, wire_13004, wire_9917, wire_3526, wire_3482, wire_13127, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_13002, wire_9915, wire_3526, wire_3482, wire_13129, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_13000, wire_9913, wire_3526, wire_3482, wire_13131, wire_13103, wire_13102, wire_13093, wire_13092, wire_13083, wire_13082, wire_12998, wire_9911, wire_3526, wire_3478, wire_13133, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_12996, wire_9909, wire_3526, wire_3478, wire_13135, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_12994, wire_9907, wire_3526, wire_3478, wire_13137, wire_13101, wire_13100, wire_13091, wire_13090, wire_13081, wire_13080, wire_12992, wire_9905, wire_3522, wire_3478, wire_13139, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_12990, wire_9903, wire_3522, wire_3478, wire_13111, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_13018, wire_9901, wire_3522, wire_3478};
    // CHNAXY TOTAL: 636
    assign wire_9781 = lut_tile_9_6_chanxy_out[0];
    assign wire_9783 = lut_tile_9_6_chanxy_out[1];
    assign wire_9785 = lut_tile_9_6_chanxy_out[2];
    assign wire_9787 = lut_tile_9_6_chanxy_out[3];
    assign wire_9789 = lut_tile_9_6_chanxy_out[4];
    assign wire_9791 = lut_tile_9_6_chanxy_out[5];
    assign wire_9793 = lut_tile_9_6_chanxy_out[6];
    assign wire_9795 = lut_tile_9_6_chanxy_out[7];
    assign wire_9797 = lut_tile_9_6_chanxy_out[8];
    assign wire_9799 = lut_tile_9_6_chanxy_out[9];
    assign wire_9801 = lut_tile_9_6_chanxy_out[10];
    assign wire_9803 = lut_tile_9_6_chanxy_out[11];
    assign wire_9805 = lut_tile_9_6_chanxy_out[12];
    assign wire_9807 = lut_tile_9_6_chanxy_out[13];
    assign wire_9809 = lut_tile_9_6_chanxy_out[14];
    assign wire_9870 = lut_tile_9_6_chanxy_out[15];
    assign wire_9872 = lut_tile_9_6_chanxy_out[16];
    assign wire_9874 = lut_tile_9_6_chanxy_out[17];
    assign wire_9876 = lut_tile_9_6_chanxy_out[18];
    assign wire_9878 = lut_tile_9_6_chanxy_out[19];
    assign wire_9880 = lut_tile_9_6_chanxy_out[20];
    assign wire_9882 = lut_tile_9_6_chanxy_out[21];
    assign wire_9884 = lut_tile_9_6_chanxy_out[22];
    assign wire_9886 = lut_tile_9_6_chanxy_out[23];
    assign wire_9888 = lut_tile_9_6_chanxy_out[24];
    assign wire_9890 = lut_tile_9_6_chanxy_out[25];
    assign wire_9892 = lut_tile_9_6_chanxy_out[26];
    assign wire_9894 = lut_tile_9_6_chanxy_out[27];
    assign wire_9896 = lut_tile_9_6_chanxy_out[28];
    assign wire_9898 = lut_tile_9_6_chanxy_out[29];
    assign wire_12991 = lut_tile_9_6_chanxy_out[30];
    assign wire_12993 = lut_tile_9_6_chanxy_out[31];
    assign wire_12995 = lut_tile_9_6_chanxy_out[32];
    assign wire_12997 = lut_tile_9_6_chanxy_out[33];
    assign wire_12999 = lut_tile_9_6_chanxy_out[34];
    assign wire_13001 = lut_tile_9_6_chanxy_out[35];
    assign wire_13003 = lut_tile_9_6_chanxy_out[36];
    assign wire_13005 = lut_tile_9_6_chanxy_out[37];
    assign wire_13007 = lut_tile_9_6_chanxy_out[38];
    assign wire_13009 = lut_tile_9_6_chanxy_out[39];
    assign wire_13011 = lut_tile_9_6_chanxy_out[40];
    assign wire_13013 = lut_tile_9_6_chanxy_out[41];
    assign wire_13015 = lut_tile_9_6_chanxy_out[42];
    assign wire_13017 = lut_tile_9_6_chanxy_out[43];
    assign wire_13019 = lut_tile_9_6_chanxy_out[44];
    assign wire_13080 = lut_tile_9_6_chanxy_out[45];
    assign wire_13082 = lut_tile_9_6_chanxy_out[46];
    assign wire_13084 = lut_tile_9_6_chanxy_out[47];
    assign wire_13086 = lut_tile_9_6_chanxy_out[48];
    assign wire_13088 = lut_tile_9_6_chanxy_out[49];
    assign wire_13090 = lut_tile_9_6_chanxy_out[50];
    assign wire_13092 = lut_tile_9_6_chanxy_out[51];
    assign wire_13094 = lut_tile_9_6_chanxy_out[52];
    assign wire_13096 = lut_tile_9_6_chanxy_out[53];
    assign wire_13098 = lut_tile_9_6_chanxy_out[54];
    assign wire_13100 = lut_tile_9_6_chanxy_out[55];
    assign wire_13102 = lut_tile_9_6_chanxy_out[56];
    assign wire_13104 = lut_tile_9_6_chanxy_out[57];
    assign wire_13106 = lut_tile_9_6_chanxy_out[58];
    assign wire_13108 = lut_tile_9_6_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_7_chanxy_in = {wire_13378, wire_9541, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9422, wire_4509, wire_13376, wire_9569, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9424, wire_4509, wire_13374, wire_9567, wire_9479, wire_9478, wire_9469, wire_9468, wire_9459, wire_9458, wire_9426, wire_4509, wire_13372, wire_9565, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9428, wire_3999, wire_13370, wire_9563, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9430, wire_3999, wire_13368, wire_9561, wire_9477, wire_9476, wire_9467, wire_9466, wire_9457, wire_9456, wire_9432, wire_3999, wire_13366, wire_9559, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9434, wire_4513, wire_3999, wire_13364, wire_9557, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9436, wire_4513, wire_3999, wire_13362, wire_9555, wire_9475, wire_9474, wire_9465, wire_9464, wire_9455, wire_9454, wire_9438, wire_4513, wire_3999, wire_13360, wire_9553, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9440, wire_4513, wire_3995, wire_13358, wire_9551, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9442, wire_4513, wire_3995, wire_13356, wire_9549, wire_9473, wire_9472, wire_9463, wire_9462, wire_9453, wire_9452, wire_9444, wire_4513, wire_3995, wire_13354, wire_9547, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9446, wire_4509, wire_3995, wire_13352, wire_9545, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9448, wire_4509, wire_3995, wire_13350, wire_9543, wire_9471, wire_9470, wire_9461, wire_9460, wire_9451, wire_9450, wire_9420, wire_4509, wire_3995, wire_13529, wire_9959, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9810, wire_4509, wire_13527, wire_9931, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9838, wire_4509, wire_13525, wire_9933, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9836, wire_4509, wire_13523, wire_9935, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9834, wire_3999, wire_13521, wire_9937, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9832, wire_3999, wire_13519, wire_9939, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9830, wire_3999, wire_13517, wire_9941, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9828, wire_4513, wire_3999, wire_13515, wire_9943, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9826, wire_4513, wire_3999, wire_13513, wire_9945, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9824, wire_4513, wire_3999, wire_13511, wire_9947, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9822, wire_4513, wire_3995, wire_13509, wire_9949, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9820, wire_4513, wire_3995, wire_13507, wire_9951, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9818, wire_4513, wire_3995, wire_13505, wire_9953, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9816, wire_4509, wire_3995, wire_13503, wire_9955, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9814, wire_4509, wire_3995, wire_13501, wire_9957, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9812, wire_4509, wire_3995, wire_13137, wire_13109, wire_13108, wire_13099, wire_13098, wire_13089, wire_13088, wire_13018, wire_9808, wire_4038, wire_13135, wire_13079, wire_13078, wire_13069, wire_13068, wire_13059, wire_13058, wire_12990, wire_9806, wire_4038, wire_13133, wire_13049, wire_13048, wire_13039, wire_13038, wire_13029, wire_13028, wire_12992, wire_9804, wire_4038, wire_13131, wire_13107, wire_13106, wire_13097, wire_13096, wire_13087, wire_13086, wire_12994, wire_9802, wire_3998, wire_13129, wire_13077, wire_13076, wire_13067, wire_13066, wire_13057, wire_13056, wire_12996, wire_9800, wire_3998, wire_13127, wire_13047, wire_13046, wire_13037, wire_13036, wire_13027, wire_13026, wire_12998, wire_9798, wire_3998, wire_13125, wire_13105, wire_13104, wire_13095, wire_13094, wire_13085, wire_13084, wire_13000, wire_9796, wire_4042, wire_3998, wire_13123, wire_13075, wire_13074, wire_13065, wire_13064, wire_13055, wire_13054, wire_13002, wire_9794, wire_4042, wire_3998, wire_13121, wire_13045, wire_13044, wire_13035, wire_13034, wire_13025, wire_13024, wire_13004, wire_9792, wire_4042, wire_3998, wire_13119, wire_13103, wire_13102, wire_13093, wire_13092, wire_13083, wire_13082, wire_13006, wire_9790, wire_4042, wire_3994, wire_13117, wire_13073, wire_13072, wire_13063, wire_13062, wire_13053, wire_13052, wire_13008, wire_9788, wire_4042, wire_3994, wire_13115, wire_13043, wire_13042, wire_13033, wire_13032, wire_13023, wire_13022, wire_13010, wire_9786, wire_4042, wire_3994, wire_13113, wire_13101, wire_13100, wire_13091, wire_13090, wire_13081, wire_13080, wire_13012, wire_9784, wire_4038, wire_3994, wire_13111, wire_13071, wire_13070, wire_13061, wire_13060, wire_13051, wire_13050, wire_13014, wire_9782, wire_4038, wire_3994, wire_13139, wire_13041, wire_13040, wire_13031, wire_13030, wire_13021, wire_13020, wire_13016, wire_9780, wire_4038, wire_3994, wire_13503, wire_13499, wire_13498, wire_13489, wire_13488, wire_13479, wire_13478, wire_13406, wire_9959, wire_4038, wire_13505, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13404, wire_9957, wire_4038, wire_13507, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13402, wire_9955, wire_4038, wire_13509, wire_13497, wire_13496, wire_13487, wire_13486, wire_13477, wire_13476, wire_13400, wire_9953, wire_3998, wire_13511, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13398, wire_9951, wire_3998, wire_13513, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13396, wire_9949, wire_3998, wire_13515, wire_13495, wire_13494, wire_13485, wire_13484, wire_13475, wire_13474, wire_13394, wire_9947, wire_4042, wire_3998, wire_13517, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13392, wire_9945, wire_4042, wire_3998, wire_13519, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13390, wire_9943, wire_4042, wire_3998, wire_13521, wire_13493, wire_13492, wire_13483, wire_13482, wire_13473, wire_13472, wire_13388, wire_9941, wire_4042, wire_3994, wire_13523, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13386, wire_9939, wire_4042, wire_3994, wire_13525, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13384, wire_9937, wire_4042, wire_3994, wire_13527, wire_13491, wire_13490, wire_13481, wire_13480, wire_13471, wire_13470, wire_13382, wire_9935, wire_4038, wire_3994, wire_13529, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13380, wire_9933, wire_4038, wire_3994, wire_13501, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13408, wire_9931, wire_4038, wire_3994};
    // CHNAXY TOTAL: 636
    assign wire_9811 = lut_tile_9_7_chanxy_out[0];
    assign wire_9813 = lut_tile_9_7_chanxy_out[1];
    assign wire_9815 = lut_tile_9_7_chanxy_out[2];
    assign wire_9817 = lut_tile_9_7_chanxy_out[3];
    assign wire_9819 = lut_tile_9_7_chanxy_out[4];
    assign wire_9821 = lut_tile_9_7_chanxy_out[5];
    assign wire_9823 = lut_tile_9_7_chanxy_out[6];
    assign wire_9825 = lut_tile_9_7_chanxy_out[7];
    assign wire_9827 = lut_tile_9_7_chanxy_out[8];
    assign wire_9829 = lut_tile_9_7_chanxy_out[9];
    assign wire_9831 = lut_tile_9_7_chanxy_out[10];
    assign wire_9833 = lut_tile_9_7_chanxy_out[11];
    assign wire_9835 = lut_tile_9_7_chanxy_out[12];
    assign wire_9837 = lut_tile_9_7_chanxy_out[13];
    assign wire_9839 = lut_tile_9_7_chanxy_out[14];
    assign wire_9900 = lut_tile_9_7_chanxy_out[15];
    assign wire_9902 = lut_tile_9_7_chanxy_out[16];
    assign wire_9904 = lut_tile_9_7_chanxy_out[17];
    assign wire_9906 = lut_tile_9_7_chanxy_out[18];
    assign wire_9908 = lut_tile_9_7_chanxy_out[19];
    assign wire_9910 = lut_tile_9_7_chanxy_out[20];
    assign wire_9912 = lut_tile_9_7_chanxy_out[21];
    assign wire_9914 = lut_tile_9_7_chanxy_out[22];
    assign wire_9916 = lut_tile_9_7_chanxy_out[23];
    assign wire_9918 = lut_tile_9_7_chanxy_out[24];
    assign wire_9920 = lut_tile_9_7_chanxy_out[25];
    assign wire_9922 = lut_tile_9_7_chanxy_out[26];
    assign wire_9924 = lut_tile_9_7_chanxy_out[27];
    assign wire_9926 = lut_tile_9_7_chanxy_out[28];
    assign wire_9928 = lut_tile_9_7_chanxy_out[29];
    assign wire_13381 = lut_tile_9_7_chanxy_out[30];
    assign wire_13383 = lut_tile_9_7_chanxy_out[31];
    assign wire_13385 = lut_tile_9_7_chanxy_out[32];
    assign wire_13387 = lut_tile_9_7_chanxy_out[33];
    assign wire_13389 = lut_tile_9_7_chanxy_out[34];
    assign wire_13391 = lut_tile_9_7_chanxy_out[35];
    assign wire_13393 = lut_tile_9_7_chanxy_out[36];
    assign wire_13395 = lut_tile_9_7_chanxy_out[37];
    assign wire_13397 = lut_tile_9_7_chanxy_out[38];
    assign wire_13399 = lut_tile_9_7_chanxy_out[39];
    assign wire_13401 = lut_tile_9_7_chanxy_out[40];
    assign wire_13403 = lut_tile_9_7_chanxy_out[41];
    assign wire_13405 = lut_tile_9_7_chanxy_out[42];
    assign wire_13407 = lut_tile_9_7_chanxy_out[43];
    assign wire_13409 = lut_tile_9_7_chanxy_out[44];
    assign wire_13470 = lut_tile_9_7_chanxy_out[45];
    assign wire_13472 = lut_tile_9_7_chanxy_out[46];
    assign wire_13474 = lut_tile_9_7_chanxy_out[47];
    assign wire_13476 = lut_tile_9_7_chanxy_out[48];
    assign wire_13478 = lut_tile_9_7_chanxy_out[49];
    assign wire_13480 = lut_tile_9_7_chanxy_out[50];
    assign wire_13482 = lut_tile_9_7_chanxy_out[51];
    assign wire_13484 = lut_tile_9_7_chanxy_out[52];
    assign wire_13486 = lut_tile_9_7_chanxy_out[53];
    assign wire_13488 = lut_tile_9_7_chanxy_out[54];
    assign wire_13490 = lut_tile_9_7_chanxy_out[55];
    assign wire_13492 = lut_tile_9_7_chanxy_out[56];
    assign wire_13494 = lut_tile_9_7_chanxy_out[57];
    assign wire_13496 = lut_tile_9_7_chanxy_out[58];
    assign wire_13498 = lut_tile_9_7_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_8_chanxy_in = {wire_13768, wire_9571, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9452, wire_5025, wire_13766, wire_9599, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9454, wire_5025, wire_13764, wire_9597, wire_9509, wire_9508, wire_9499, wire_9498, wire_9489, wire_9488, wire_9456, wire_5025, wire_13762, wire_9595, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9458, wire_4515, wire_13760, wire_9593, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9460, wire_4515, wire_13758, wire_9591, wire_9507, wire_9506, wire_9497, wire_9496, wire_9487, wire_9486, wire_9462, wire_4515, wire_13756, wire_9589, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9464, wire_5029, wire_4515, wire_13754, wire_9587, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9466, wire_5029, wire_4515, wire_13752, wire_9585, wire_9505, wire_9504, wire_9495, wire_9494, wire_9485, wire_9484, wire_9468, wire_5029, wire_4515, wire_13750, wire_9583, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9470, wire_5029, wire_4511, wire_13748, wire_9581, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9472, wire_5029, wire_4511, wire_13746, wire_9579, wire_9503, wire_9502, wire_9493, wire_9492, wire_9483, wire_9482, wire_9474, wire_5029, wire_4511, wire_13744, wire_9577, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9476, wire_5025, wire_4511, wire_13742, wire_9575, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9478, wire_5025, wire_4511, wire_13740, wire_9573, wire_9501, wire_9500, wire_9491, wire_9490, wire_9481, wire_9480, wire_9450, wire_5025, wire_4511, wire_13919, wire_9989, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9840, wire_5025, wire_13917, wire_9961, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9868, wire_5025, wire_13915, wire_9963, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9866, wire_5025, wire_13913, wire_9965, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9864, wire_4515, wire_13911, wire_9967, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9862, wire_4515, wire_13909, wire_9969, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9860, wire_4515, wire_13907, wire_9971, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9858, wire_5029, wire_4515, wire_13905, wire_9973, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9856, wire_5029, wire_4515, wire_13903, wire_9975, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9854, wire_5029, wire_4515, wire_13901, wire_9977, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9852, wire_5029, wire_4511, wire_13899, wire_9979, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9850, wire_5029, wire_4511, wire_13897, wire_9981, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9848, wire_5029, wire_4511, wire_13895, wire_9983, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9846, wire_5025, wire_4511, wire_13893, wire_9985, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9844, wire_5025, wire_4511, wire_13891, wire_9987, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9842, wire_5025, wire_4511, wire_13527, wire_13499, wire_13498, wire_13489, wire_13488, wire_13479, wire_13478, wire_13408, wire_9838, wire_4554, wire_13525, wire_13469, wire_13468, wire_13459, wire_13458, wire_13449, wire_13448, wire_13380, wire_9836, wire_4554, wire_13523, wire_13439, wire_13438, wire_13429, wire_13428, wire_13419, wire_13418, wire_13382, wire_9834, wire_4554, wire_13521, wire_13497, wire_13496, wire_13487, wire_13486, wire_13477, wire_13476, wire_13384, wire_9832, wire_4514, wire_13519, wire_13467, wire_13466, wire_13457, wire_13456, wire_13447, wire_13446, wire_13386, wire_9830, wire_4514, wire_13517, wire_13437, wire_13436, wire_13427, wire_13426, wire_13417, wire_13416, wire_13388, wire_9828, wire_4514, wire_13515, wire_13495, wire_13494, wire_13485, wire_13484, wire_13475, wire_13474, wire_13390, wire_9826, wire_4558, wire_4514, wire_13513, wire_13465, wire_13464, wire_13455, wire_13454, wire_13445, wire_13444, wire_13392, wire_9824, wire_4558, wire_4514, wire_13511, wire_13435, wire_13434, wire_13425, wire_13424, wire_13415, wire_13414, wire_13394, wire_9822, wire_4558, wire_4514, wire_13509, wire_13493, wire_13492, wire_13483, wire_13482, wire_13473, wire_13472, wire_13396, wire_9820, wire_4558, wire_4510, wire_13507, wire_13463, wire_13462, wire_13453, wire_13452, wire_13443, wire_13442, wire_13398, wire_9818, wire_4558, wire_4510, wire_13505, wire_13433, wire_13432, wire_13423, wire_13422, wire_13413, wire_13412, wire_13400, wire_9816, wire_4558, wire_4510, wire_13503, wire_13491, wire_13490, wire_13481, wire_13480, wire_13471, wire_13470, wire_13402, wire_9814, wire_4554, wire_4510, wire_13501, wire_13461, wire_13460, wire_13451, wire_13450, wire_13441, wire_13440, wire_13404, wire_9812, wire_4554, wire_4510, wire_13529, wire_13431, wire_13430, wire_13421, wire_13420, wire_13411, wire_13410, wire_13406, wire_9810, wire_4554, wire_4510, wire_13893, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13796, wire_9989, wire_4554, wire_13895, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13794, wire_9987, wire_4554, wire_13897, wire_13889, wire_13888, wire_13879, wire_13878, wire_13869, wire_13868, wire_13792, wire_9985, wire_4554, wire_13899, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13790, wire_9983, wire_4514, wire_13901, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13788, wire_9981, wire_4514, wire_13903, wire_13887, wire_13886, wire_13877, wire_13876, wire_13867, wire_13866, wire_13786, wire_9979, wire_4514, wire_13905, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13784, wire_9977, wire_4558, wire_4514, wire_13907, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13782, wire_9975, wire_4558, wire_4514, wire_13909, wire_13885, wire_13884, wire_13875, wire_13874, wire_13865, wire_13864, wire_13780, wire_9973, wire_4558, wire_4514, wire_13911, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13778, wire_9971, wire_4558, wire_4510, wire_13913, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13776, wire_9969, wire_4558, wire_4510, wire_13915, wire_13883, wire_13882, wire_13873, wire_13872, wire_13863, wire_13862, wire_13774, wire_9967, wire_4558, wire_4510, wire_13917, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13772, wire_9965, wire_4554, wire_4510, wire_13919, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13770, wire_9963, wire_4554, wire_4510, wire_13891, wire_13881, wire_13880, wire_13871, wire_13870, wire_13861, wire_13860, wire_13798, wire_9961, wire_4554, wire_4510};
    // CHNAXY TOTAL: 636
    assign wire_9841 = lut_tile_9_8_chanxy_out[0];
    assign wire_9843 = lut_tile_9_8_chanxy_out[1];
    assign wire_9845 = lut_tile_9_8_chanxy_out[2];
    assign wire_9847 = lut_tile_9_8_chanxy_out[3];
    assign wire_9849 = lut_tile_9_8_chanxy_out[4];
    assign wire_9851 = lut_tile_9_8_chanxy_out[5];
    assign wire_9853 = lut_tile_9_8_chanxy_out[6];
    assign wire_9855 = lut_tile_9_8_chanxy_out[7];
    assign wire_9857 = lut_tile_9_8_chanxy_out[8];
    assign wire_9859 = lut_tile_9_8_chanxy_out[9];
    assign wire_9861 = lut_tile_9_8_chanxy_out[10];
    assign wire_9863 = lut_tile_9_8_chanxy_out[11];
    assign wire_9865 = lut_tile_9_8_chanxy_out[12];
    assign wire_9867 = lut_tile_9_8_chanxy_out[13];
    assign wire_9869 = lut_tile_9_8_chanxy_out[14];
    assign wire_9930 = lut_tile_9_8_chanxy_out[15];
    assign wire_9932 = lut_tile_9_8_chanxy_out[16];
    assign wire_9934 = lut_tile_9_8_chanxy_out[17];
    assign wire_9936 = lut_tile_9_8_chanxy_out[18];
    assign wire_9938 = lut_tile_9_8_chanxy_out[19];
    assign wire_9940 = lut_tile_9_8_chanxy_out[20];
    assign wire_9942 = lut_tile_9_8_chanxy_out[21];
    assign wire_9944 = lut_tile_9_8_chanxy_out[22];
    assign wire_9946 = lut_tile_9_8_chanxy_out[23];
    assign wire_9948 = lut_tile_9_8_chanxy_out[24];
    assign wire_9950 = lut_tile_9_8_chanxy_out[25];
    assign wire_9952 = lut_tile_9_8_chanxy_out[26];
    assign wire_9954 = lut_tile_9_8_chanxy_out[27];
    assign wire_9956 = lut_tile_9_8_chanxy_out[28];
    assign wire_9958 = lut_tile_9_8_chanxy_out[29];
    assign wire_13771 = lut_tile_9_8_chanxy_out[30];
    assign wire_13773 = lut_tile_9_8_chanxy_out[31];
    assign wire_13775 = lut_tile_9_8_chanxy_out[32];
    assign wire_13777 = lut_tile_9_8_chanxy_out[33];
    assign wire_13779 = lut_tile_9_8_chanxy_out[34];
    assign wire_13781 = lut_tile_9_8_chanxy_out[35];
    assign wire_13783 = lut_tile_9_8_chanxy_out[36];
    assign wire_13785 = lut_tile_9_8_chanxy_out[37];
    assign wire_13787 = lut_tile_9_8_chanxy_out[38];
    assign wire_13789 = lut_tile_9_8_chanxy_out[39];
    assign wire_13791 = lut_tile_9_8_chanxy_out[40];
    assign wire_13793 = lut_tile_9_8_chanxy_out[41];
    assign wire_13795 = lut_tile_9_8_chanxy_out[42];
    assign wire_13797 = lut_tile_9_8_chanxy_out[43];
    assign wire_13799 = lut_tile_9_8_chanxy_out[44];
    assign wire_13860 = lut_tile_9_8_chanxy_out[45];
    assign wire_13862 = lut_tile_9_8_chanxy_out[46];
    assign wire_13864 = lut_tile_9_8_chanxy_out[47];
    assign wire_13866 = lut_tile_9_8_chanxy_out[48];
    assign wire_13868 = lut_tile_9_8_chanxy_out[49];
    assign wire_13870 = lut_tile_9_8_chanxy_out[50];
    assign wire_13872 = lut_tile_9_8_chanxy_out[51];
    assign wire_13874 = lut_tile_9_8_chanxy_out[52];
    assign wire_13876 = lut_tile_9_8_chanxy_out[53];
    assign wire_13878 = lut_tile_9_8_chanxy_out[54];
    assign wire_13880 = lut_tile_9_8_chanxy_out[55];
    assign wire_13882 = lut_tile_9_8_chanxy_out[56];
    assign wire_13884 = lut_tile_9_8_chanxy_out[57];
    assign wire_13886 = lut_tile_9_8_chanxy_out[58];
    assign wire_13888 = lut_tile_9_8_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_9_chanxy_in = {wire_14158, wire_9601, wire_9569, wire_9568, wire_9559, wire_9558, wire_9549, wire_9548, wire_9482, wire_5541, wire_14156, wire_9629, wire_9539, wire_9538, wire_9529, wire_9528, wire_9519, wire_9518, wire_9484, wire_5541, wire_14154, wire_9627, wire_9599, wire_9598, wire_9589, wire_9588, wire_9579, wire_9578, wire_9486, wire_5541, wire_14152, wire_9625, wire_9567, wire_9566, wire_9557, wire_9556, wire_9547, wire_9546, wire_9488, wire_5031, wire_14150, wire_9623, wire_9537, wire_9536, wire_9527, wire_9526, wire_9517, wire_9516, wire_9490, wire_5031, wire_14148, wire_9621, wire_9597, wire_9596, wire_9587, wire_9586, wire_9577, wire_9576, wire_9492, wire_5031, wire_14146, wire_9619, wire_9565, wire_9564, wire_9555, wire_9554, wire_9545, wire_9544, wire_9494, wire_5545, wire_5031, wire_14144, wire_9617, wire_9535, wire_9534, wire_9525, wire_9524, wire_9515, wire_9514, wire_9496, wire_5545, wire_5031, wire_14142, wire_9615, wire_9595, wire_9594, wire_9585, wire_9584, wire_9575, wire_9574, wire_9498, wire_5545, wire_5031, wire_14140, wire_9613, wire_9563, wire_9562, wire_9553, wire_9552, wire_9543, wire_9542, wire_9500, wire_5545, wire_5027, wire_14138, wire_9611, wire_9533, wire_9532, wire_9523, wire_9522, wire_9513, wire_9512, wire_9502, wire_5545, wire_5027, wire_14136, wire_9609, wire_9593, wire_9592, wire_9583, wire_9582, wire_9573, wire_9572, wire_9504, wire_5545, wire_5027, wire_14134, wire_9607, wire_9561, wire_9560, wire_9551, wire_9550, wire_9541, wire_9540, wire_9506, wire_5541, wire_5027, wire_14132, wire_9605, wire_9531, wire_9530, wire_9521, wire_9520, wire_9511, wire_9510, wire_9508, wire_5541, wire_5027, wire_14130, wire_9603, wire_9591, wire_9590, wire_9581, wire_9580, wire_9571, wire_9570, wire_9480, wire_5541, wire_5027, wire_14309, wire_10019, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9870, wire_5541, wire_14307, wire_9991, wire_9989, wire_9988, wire_9979, wire_9978, wire_9969, wire_9968, wire_9898, wire_5541, wire_14305, wire_9993, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9896, wire_5541, wire_14303, wire_9995, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9894, wire_5031, wire_14301, wire_9997, wire_9987, wire_9986, wire_9977, wire_9976, wire_9967, wire_9966, wire_9892, wire_5031, wire_14299, wire_9999, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9890, wire_5031, wire_14297, wire_10001, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9888, wire_5545, wire_5031, wire_14295, wire_10003, wire_9985, wire_9984, wire_9975, wire_9974, wire_9965, wire_9964, wire_9886, wire_5545, wire_5031, wire_14293, wire_10005, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9884, wire_5545, wire_5031, wire_14291, wire_10007, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9882, wire_5545, wire_5027, wire_14289, wire_10009, wire_9983, wire_9982, wire_9973, wire_9972, wire_9963, wire_9962, wire_9880, wire_5545, wire_5027, wire_14287, wire_10011, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9878, wire_5545, wire_5027, wire_14285, wire_10013, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9876, wire_5541, wire_5027, wire_14283, wire_10015, wire_9981, wire_9980, wire_9971, wire_9970, wire_9961, wire_9960, wire_9874, wire_5541, wire_5027, wire_14281, wire_10017, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9872, wire_5541, wire_5027, wire_13917, wire_13859, wire_13858, wire_13849, wire_13848, wire_13839, wire_13838, wire_13798, wire_9868, wire_5070, wire_13915, wire_13829, wire_13828, wire_13819, wire_13818, wire_13809, wire_13808, wire_13770, wire_9866, wire_5070, wire_13913, wire_13889, wire_13888, wire_13879, wire_13878, wire_13869, wire_13868, wire_13772, wire_9864, wire_5070, wire_13911, wire_13857, wire_13856, wire_13847, wire_13846, wire_13837, wire_13836, wire_13774, wire_9862, wire_5030, wire_13909, wire_13827, wire_13826, wire_13817, wire_13816, wire_13807, wire_13806, wire_13776, wire_9860, wire_5030, wire_13907, wire_13887, wire_13886, wire_13877, wire_13876, wire_13867, wire_13866, wire_13778, wire_9858, wire_5030, wire_13905, wire_13855, wire_13854, wire_13845, wire_13844, wire_13835, wire_13834, wire_13780, wire_9856, wire_5074, wire_5030, wire_13903, wire_13825, wire_13824, wire_13815, wire_13814, wire_13805, wire_13804, wire_13782, wire_9854, wire_5074, wire_5030, wire_13901, wire_13885, wire_13884, wire_13875, wire_13874, wire_13865, wire_13864, wire_13784, wire_9852, wire_5074, wire_5030, wire_13899, wire_13853, wire_13852, wire_13843, wire_13842, wire_13833, wire_13832, wire_13786, wire_9850, wire_5074, wire_5026, wire_13897, wire_13823, wire_13822, wire_13813, wire_13812, wire_13803, wire_13802, wire_13788, wire_9848, wire_5074, wire_5026, wire_13895, wire_13883, wire_13882, wire_13873, wire_13872, wire_13863, wire_13862, wire_13790, wire_9846, wire_5074, wire_5026, wire_13893, wire_13851, wire_13850, wire_13841, wire_13840, wire_13831, wire_13830, wire_13792, wire_9844, wire_5070, wire_5026, wire_13891, wire_13821, wire_13820, wire_13811, wire_13810, wire_13801, wire_13800, wire_13794, wire_9842, wire_5070, wire_5026, wire_13919, wire_13881, wire_13880, wire_13871, wire_13870, wire_13861, wire_13860, wire_13796, wire_9840, wire_5070, wire_5026, wire_14283, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14186, wire_10019, wire_5070, wire_14285, wire_14279, wire_14278, wire_14269, wire_14268, wire_14259, wire_14258, wire_14184, wire_10017, wire_5070, wire_14287, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14182, wire_10015, wire_5070, wire_14289, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14180, wire_10013, wire_5030, wire_14291, wire_14277, wire_14276, wire_14267, wire_14266, wire_14257, wire_14256, wire_14178, wire_10011, wire_5030, wire_14293, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14176, wire_10009, wire_5030, wire_14295, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14174, wire_10007, wire_5074, wire_5030, wire_14297, wire_14275, wire_14274, wire_14265, wire_14264, wire_14255, wire_14254, wire_14172, wire_10005, wire_5074, wire_5030, wire_14299, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14170, wire_10003, wire_5074, wire_5030, wire_14301, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14168, wire_10001, wire_5074, wire_5026, wire_14303, wire_14273, wire_14272, wire_14263, wire_14262, wire_14253, wire_14252, wire_14166, wire_9999, wire_5074, wire_5026, wire_14305, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14164, wire_9997, wire_5074, wire_5026, wire_14307, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14162, wire_9995, wire_5070, wire_5026, wire_14309, wire_14271, wire_14270, wire_14261, wire_14260, wire_14251, wire_14250, wire_14160, wire_9993, wire_5070, wire_5026, wire_14281, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14188, wire_9991, wire_5070, wire_5026};
    // CHNAXY TOTAL: 636
    assign wire_9871 = lut_tile_9_9_chanxy_out[0];
    assign wire_9873 = lut_tile_9_9_chanxy_out[1];
    assign wire_9875 = lut_tile_9_9_chanxy_out[2];
    assign wire_9877 = lut_tile_9_9_chanxy_out[3];
    assign wire_9879 = lut_tile_9_9_chanxy_out[4];
    assign wire_9881 = lut_tile_9_9_chanxy_out[5];
    assign wire_9883 = lut_tile_9_9_chanxy_out[6];
    assign wire_9885 = lut_tile_9_9_chanxy_out[7];
    assign wire_9887 = lut_tile_9_9_chanxy_out[8];
    assign wire_9889 = lut_tile_9_9_chanxy_out[9];
    assign wire_9891 = lut_tile_9_9_chanxy_out[10];
    assign wire_9893 = lut_tile_9_9_chanxy_out[11];
    assign wire_9895 = lut_tile_9_9_chanxy_out[12];
    assign wire_9897 = lut_tile_9_9_chanxy_out[13];
    assign wire_9899 = lut_tile_9_9_chanxy_out[14];
    assign wire_9960 = lut_tile_9_9_chanxy_out[15];
    assign wire_9962 = lut_tile_9_9_chanxy_out[16];
    assign wire_9964 = lut_tile_9_9_chanxy_out[17];
    assign wire_9966 = lut_tile_9_9_chanxy_out[18];
    assign wire_9968 = lut_tile_9_9_chanxy_out[19];
    assign wire_9970 = lut_tile_9_9_chanxy_out[20];
    assign wire_9972 = lut_tile_9_9_chanxy_out[21];
    assign wire_9974 = lut_tile_9_9_chanxy_out[22];
    assign wire_9976 = lut_tile_9_9_chanxy_out[23];
    assign wire_9978 = lut_tile_9_9_chanxy_out[24];
    assign wire_9980 = lut_tile_9_9_chanxy_out[25];
    assign wire_9982 = lut_tile_9_9_chanxy_out[26];
    assign wire_9984 = lut_tile_9_9_chanxy_out[27];
    assign wire_9986 = lut_tile_9_9_chanxy_out[28];
    assign wire_9988 = lut_tile_9_9_chanxy_out[29];
    assign wire_14161 = lut_tile_9_9_chanxy_out[30];
    assign wire_14163 = lut_tile_9_9_chanxy_out[31];
    assign wire_14165 = lut_tile_9_9_chanxy_out[32];
    assign wire_14167 = lut_tile_9_9_chanxy_out[33];
    assign wire_14169 = lut_tile_9_9_chanxy_out[34];
    assign wire_14171 = lut_tile_9_9_chanxy_out[35];
    assign wire_14173 = lut_tile_9_9_chanxy_out[36];
    assign wire_14175 = lut_tile_9_9_chanxy_out[37];
    assign wire_14177 = lut_tile_9_9_chanxy_out[38];
    assign wire_14179 = lut_tile_9_9_chanxy_out[39];
    assign wire_14181 = lut_tile_9_9_chanxy_out[40];
    assign wire_14183 = lut_tile_9_9_chanxy_out[41];
    assign wire_14185 = lut_tile_9_9_chanxy_out[42];
    assign wire_14187 = lut_tile_9_9_chanxy_out[43];
    assign wire_14189 = lut_tile_9_9_chanxy_out[44];
    assign wire_14250 = lut_tile_9_9_chanxy_out[45];
    assign wire_14252 = lut_tile_9_9_chanxy_out[46];
    assign wire_14254 = lut_tile_9_9_chanxy_out[47];
    assign wire_14256 = lut_tile_9_9_chanxy_out[48];
    assign wire_14258 = lut_tile_9_9_chanxy_out[49];
    assign wire_14260 = lut_tile_9_9_chanxy_out[50];
    assign wire_14262 = lut_tile_9_9_chanxy_out[51];
    assign wire_14264 = lut_tile_9_9_chanxy_out[52];
    assign wire_14266 = lut_tile_9_9_chanxy_out[53];
    assign wire_14268 = lut_tile_9_9_chanxy_out[54];
    assign wire_14270 = lut_tile_9_9_chanxy_out[55];
    assign wire_14272 = lut_tile_9_9_chanxy_out[56];
    assign wire_14274 = lut_tile_9_9_chanxy_out[57];
    assign wire_14276 = lut_tile_9_9_chanxy_out[58];
    assign wire_14278 = lut_tile_9_9_chanxy_out[59];
   // CHANXY OUT
    assign lut_tile_9_10_chanxy_in = {wire_14548, wire_9614, wire_9592, wire_9568, wire_9516, wire_6070, wire_6064, wire_6055, wire_6049, wire_14546, wire_9606, wire_9584, wire_9560, wire_9538, wire_6070, wire_6064, wire_6055, wire_6049, wire_14544, wire_9628, wire_9576, wire_9552, wire_9530, wire_6070, wire_6064, wire_6055, wire_6049, wire_14542, wire_9620, wire_9598, wire_9544, wire_9522, wire_6070, wire_6061, wire_6055, wire_5547, wire_14540, wire_9612, wire_9590, wire_9566, wire_9514, wire_6070, wire_6061, wire_6055, wire_5547, wire_14538, wire_9604, wire_9582, wire_9558, wire_9536, wire_6070, wire_6061, wire_6055, wire_5547, wire_14536, wire_9626, wire_9574, wire_9550, wire_9528, wire_6067, wire_6061, wire_6052, wire_5547, wire_14534, wire_9618, wire_9596, wire_9542, wire_9520, wire_6067, wire_6061, wire_6052, wire_5547, wire_14532, wire_9610, wire_9588, wire_9564, wire_9512, wire_6067, wire_6061, wire_6052, wire_5547, wire_14530, wire_9602, wire_9580, wire_9556, wire_9534, wire_6067, wire_6058, wire_6052, wire_5543, wire_14528, wire_9624, wire_9572, wire_9548, wire_9526, wire_6067, wire_6058, wire_6052, wire_5543, wire_14526, wire_9616, wire_9594, wire_9540, wire_9518, wire_6067, wire_6058, wire_6052, wire_5543, wire_14524, wire_9608, wire_9586, wire_9562, wire_9510, wire_6064, wire_6058, wire_6049, wire_5543, wire_14522, wire_9600, wire_9578, wire_9554, wire_9532, wire_6064, wire_6058, wire_6049, wire_5543, wire_14520, wire_9622, wire_9570, wire_9546, wire_9524, wire_6064, wire_6058, wire_6049, wire_5543, wire_14699, wire_9996, wire_9974, wire_9952, wire_9928, wire_6070, wire_6064, wire_6055, wire_6049, wire_14697, wire_10018, wire_9966, wire_9944, wire_9920, wire_6070, wire_6064, wire_6055, wire_6049, wire_14695, wire_10010, wire_9988, wire_9936, wire_9912, wire_6070, wire_6064, wire_6055, wire_6049, wire_14693, wire_10002, wire_9980, wire_9958, wire_9904, wire_6070, wire_6061, wire_6055, wire_5547, wire_14691, wire_9994, wire_9972, wire_9950, wire_9926, wire_6070, wire_6061, wire_6055, wire_5547, wire_14689, wire_10016, wire_9964, wire_9942, wire_9918, wire_6070, wire_6061, wire_6055, wire_5547, wire_14687, wire_10008, wire_9986, wire_9934, wire_9910, wire_6067, wire_6061, wire_6052, wire_5547, wire_14685, wire_10000, wire_9978, wire_9956, wire_9902, wire_6067, wire_6061, wire_6052, wire_5547, wire_14683, wire_9992, wire_9970, wire_9948, wire_9924, wire_6067, wire_6061, wire_6052, wire_5547, wire_14681, wire_10014, wire_9962, wire_9940, wire_9916, wire_6067, wire_6058, wire_6052, wire_5543, wire_14679, wire_10006, wire_9984, wire_9932, wire_9908, wire_6067, wire_6058, wire_6052, wire_5543, wire_14677, wire_9998, wire_9976, wire_9954, wire_9900, wire_6067, wire_6058, wire_6052, wire_5543, wire_14675, wire_9990, wire_9968, wire_9946, wire_9922, wire_6064, wire_6058, wire_6049, wire_5543, wire_14673, wire_10012, wire_9960, wire_9938, wire_9914, wire_6064, wire_6058, wire_6049, wire_5543, wire_14671, wire_10004, wire_9982, wire_9930, wire_9906, wire_6064, wire_6058, wire_6049, wire_5543, wire_14669, wire_14668, wire_14307, wire_14219, wire_14218, wire_14209, wire_14208, wire_14199, wire_14198, wire_14188, wire_9898, wire_5586, wire_14653, wire_14652, wire_14305, wire_14279, wire_14278, wire_14269, wire_14268, wire_14259, wire_14258, wire_14160, wire_9896, wire_5586, wire_14637, wire_14636, wire_14303, wire_14249, wire_14248, wire_14239, wire_14238, wire_14229, wire_14228, wire_14162, wire_9894, wire_5586, wire_14651, wire_14650, wire_14301, wire_14217, wire_14216, wire_14207, wire_14206, wire_14197, wire_14196, wire_14164, wire_9892, wire_5546, wire_14665, wire_14664, wire_14299, wire_14277, wire_14276, wire_14267, wire_14266, wire_14257, wire_14256, wire_14166, wire_9890, wire_5546, wire_14619, wire_14618, wire_14297, wire_14247, wire_14246, wire_14237, wire_14236, wire_14227, wire_14226, wire_14168, wire_9888, wire_5546, wire_14663, wire_14662, wire_14295, wire_14215, wire_14214, wire_14205, wire_14204, wire_14195, wire_14194, wire_14170, wire_9886, wire_5590, wire_5546, wire_14647, wire_14646, wire_14293, wire_14275, wire_14274, wire_14265, wire_14264, wire_14255, wire_14254, wire_14172, wire_9884, wire_5590, wire_5546, wire_14631, wire_14630, wire_14291, wire_14245, wire_14244, wire_14235, wire_14234, wire_14225, wire_14224, wire_14174, wire_9882, wire_5590, wire_5546, wire_14645, wire_14644, wire_5590, wire_14289, wire_14213, wire_14212, wire_14203, wire_14202, wire_14193, wire_14192, wire_14176, wire_9880, wire_5590, wire_5542, wire_14659, wire_14658, wire_5590, wire_14287, wire_14273, wire_14272, wire_14263, wire_14262, wire_14253, wire_14252, wire_14178, wire_9878, wire_5590, wire_5542, wire_14613, wire_14612, wire_5586, wire_14285, wire_14243, wire_14242, wire_14233, wire_14232, wire_14223, wire_14222, wire_14180, wire_9876, wire_5590, wire_5542, wire_14657, wire_14656, wire_5546, wire_14283, wire_14211, wire_14210, wire_14201, wire_14200, wire_14191, wire_14190, wire_14182, wire_9874, wire_5586, wire_5542, wire_14641, wire_14640, wire_5546, wire_14281, wire_14271, wire_14270, wire_14261, wire_14260, wire_14251, wire_14250, wire_14184, wire_9872, wire_5586, wire_5542, wire_14625, wire_14624, wire_5542, wire_14309, wire_14241, wire_14240, wire_14231, wire_14230, wire_14221, wire_14220, wire_14186, wire_9870, wire_5586, wire_5542, wire_14683, wire_14562, wire_14697, wire_14576, wire_14607, wire_14606, wire_14695, wire_14574, wire_14679, wire_14558, wire_14589, wire_14588, wire_14677, wire_14556, wire_14691, wire_14570, wire_14601, wire_14600, wire_14689, wire_14568, wire_5590, wire_14673, wire_14552, wire_5586, wire_14583, wire_14582, wire_5586, wire_14671, wire_14550, wire_5546, wire_14685, wire_14564, wire_5542, wire_14595, wire_14594, wire_5542, wire_14639, wire_14638, wire_14667, wire_14666, wire_14593, wire_14592, wire_14621, wire_14620, wire_14649, wire_14648, wire_14605, wire_14604, wire_14633, wire_14632, wire_14661, wire_14660, wire_14587, wire_14586, wire_14615, wire_14614, wire_5590, wire_14643, wire_14642, wire_5586, wire_14599, wire_14598, wire_5586, wire_14627, wire_14626, wire_5546, wire_14655, wire_14654, wire_5542, wire_14581, wire_14580, wire_5542, wire_14699, wire_14578, wire_14609, wire_14608, wire_14623, wire_14622, wire_14681, wire_14560, wire_14591, wire_14590, wire_14635, wire_14634, wire_14693, wire_14572, wire_14603, wire_14602, wire_14617, wire_14616, wire_14675, wire_14554, wire_5590, wire_14585, wire_14584, wire_5590, wire_14629, wire_14628, wire_5586, wire_14687, wire_14566, wire_5546, wire_14597, wire_14596, wire_5546, wire_14611, wire_14610, wire_5542};
    // CHNAXY TOTAL: 573
    assign wire_9901 = lut_tile_9_10_chanxy_out[0];
    assign wire_9903 = lut_tile_9_10_chanxy_out[1];
    assign wire_9905 = lut_tile_9_10_chanxy_out[2];
    assign wire_9907 = lut_tile_9_10_chanxy_out[3];
    assign wire_9909 = lut_tile_9_10_chanxy_out[4];
    assign wire_9911 = lut_tile_9_10_chanxy_out[5];
    assign wire_9913 = lut_tile_9_10_chanxy_out[6];
    assign wire_9915 = lut_tile_9_10_chanxy_out[7];
    assign wire_9917 = lut_tile_9_10_chanxy_out[8];
    assign wire_9919 = lut_tile_9_10_chanxy_out[9];
    assign wire_9921 = lut_tile_9_10_chanxy_out[10];
    assign wire_9923 = lut_tile_9_10_chanxy_out[11];
    assign wire_9925 = lut_tile_9_10_chanxy_out[12];
    assign wire_9927 = lut_tile_9_10_chanxy_out[13];
    assign wire_9929 = lut_tile_9_10_chanxy_out[14];
    assign wire_9931 = lut_tile_9_10_chanxy_out[15];
    assign wire_9933 = lut_tile_9_10_chanxy_out[16];
    assign wire_9935 = lut_tile_9_10_chanxy_out[17];
    assign wire_9937 = lut_tile_9_10_chanxy_out[18];
    assign wire_9939 = lut_tile_9_10_chanxy_out[19];
    assign wire_9941 = lut_tile_9_10_chanxy_out[20];
    assign wire_9943 = lut_tile_9_10_chanxy_out[21];
    assign wire_9945 = lut_tile_9_10_chanxy_out[22];
    assign wire_9947 = lut_tile_9_10_chanxy_out[23];
    assign wire_9949 = lut_tile_9_10_chanxy_out[24];
    assign wire_9951 = lut_tile_9_10_chanxy_out[25];
    assign wire_9953 = lut_tile_9_10_chanxy_out[26];
    assign wire_9955 = lut_tile_9_10_chanxy_out[27];
    assign wire_9957 = lut_tile_9_10_chanxy_out[28];
    assign wire_9959 = lut_tile_9_10_chanxy_out[29];
    assign wire_9961 = lut_tile_9_10_chanxy_out[30];
    assign wire_9963 = lut_tile_9_10_chanxy_out[31];
    assign wire_9965 = lut_tile_9_10_chanxy_out[32];
    assign wire_9967 = lut_tile_9_10_chanxy_out[33];
    assign wire_9969 = lut_tile_9_10_chanxy_out[34];
    assign wire_9971 = lut_tile_9_10_chanxy_out[35];
    assign wire_9973 = lut_tile_9_10_chanxy_out[36];
    assign wire_9975 = lut_tile_9_10_chanxy_out[37];
    assign wire_9977 = lut_tile_9_10_chanxy_out[38];
    assign wire_9979 = lut_tile_9_10_chanxy_out[39];
    assign wire_9981 = lut_tile_9_10_chanxy_out[40];
    assign wire_9983 = lut_tile_9_10_chanxy_out[41];
    assign wire_9985 = lut_tile_9_10_chanxy_out[42];
    assign wire_9987 = lut_tile_9_10_chanxy_out[43];
    assign wire_9989 = lut_tile_9_10_chanxy_out[44];
    assign wire_9990 = lut_tile_9_10_chanxy_out[45];
    assign wire_9991 = lut_tile_9_10_chanxy_out[46];
    assign wire_9992 = lut_tile_9_10_chanxy_out[47];
    assign wire_9993 = lut_tile_9_10_chanxy_out[48];
    assign wire_9994 = lut_tile_9_10_chanxy_out[49];
    assign wire_9995 = lut_tile_9_10_chanxy_out[50];
    assign wire_9996 = lut_tile_9_10_chanxy_out[51];
    assign wire_9997 = lut_tile_9_10_chanxy_out[52];
    assign wire_9998 = lut_tile_9_10_chanxy_out[53];
    assign wire_9999 = lut_tile_9_10_chanxy_out[54];
    assign wire_10000 = lut_tile_9_10_chanxy_out[55];
    assign wire_10001 = lut_tile_9_10_chanxy_out[56];
    assign wire_10002 = lut_tile_9_10_chanxy_out[57];
    assign wire_10003 = lut_tile_9_10_chanxy_out[58];
    assign wire_10004 = lut_tile_9_10_chanxy_out[59];
    assign wire_10005 = lut_tile_9_10_chanxy_out[60];
    assign wire_10006 = lut_tile_9_10_chanxy_out[61];
    assign wire_10007 = lut_tile_9_10_chanxy_out[62];
    assign wire_10008 = lut_tile_9_10_chanxy_out[63];
    assign wire_10009 = lut_tile_9_10_chanxy_out[64];
    assign wire_10010 = lut_tile_9_10_chanxy_out[65];
    assign wire_10011 = lut_tile_9_10_chanxy_out[66];
    assign wire_10012 = lut_tile_9_10_chanxy_out[67];
    assign wire_10013 = lut_tile_9_10_chanxy_out[68];
    assign wire_10014 = lut_tile_9_10_chanxy_out[69];
    assign wire_10015 = lut_tile_9_10_chanxy_out[70];
    assign wire_10016 = lut_tile_9_10_chanxy_out[71];
    assign wire_10017 = lut_tile_9_10_chanxy_out[72];
    assign wire_10018 = lut_tile_9_10_chanxy_out[73];
    assign wire_10019 = lut_tile_9_10_chanxy_out[74];
    assign wire_14551 = lut_tile_9_10_chanxy_out[75];
    assign wire_14553 = lut_tile_9_10_chanxy_out[76];
    assign wire_14555 = lut_tile_9_10_chanxy_out[77];
    assign wire_14557 = lut_tile_9_10_chanxy_out[78];
    assign wire_14559 = lut_tile_9_10_chanxy_out[79];
    assign wire_14561 = lut_tile_9_10_chanxy_out[80];
    assign wire_14563 = lut_tile_9_10_chanxy_out[81];
    assign wire_14565 = lut_tile_9_10_chanxy_out[82];
    assign wire_14567 = lut_tile_9_10_chanxy_out[83];
    assign wire_14569 = lut_tile_9_10_chanxy_out[84];
    assign wire_14571 = lut_tile_9_10_chanxy_out[85];
    assign wire_14573 = lut_tile_9_10_chanxy_out[86];
    assign wire_14575 = lut_tile_9_10_chanxy_out[87];
    assign wire_14577 = lut_tile_9_10_chanxy_out[88];
    assign wire_14579 = lut_tile_9_10_chanxy_out[89];
    assign wire_14640 = lut_tile_9_10_chanxy_out[90];
    assign wire_14642 = lut_tile_9_10_chanxy_out[91];
    assign wire_14644 = lut_tile_9_10_chanxy_out[92];
    assign wire_14646 = lut_tile_9_10_chanxy_out[93];
    assign wire_14648 = lut_tile_9_10_chanxy_out[94];
    assign wire_14650 = lut_tile_9_10_chanxy_out[95];
    assign wire_14652 = lut_tile_9_10_chanxy_out[96];
    assign wire_14654 = lut_tile_9_10_chanxy_out[97];
    assign wire_14656 = lut_tile_9_10_chanxy_out[98];
    assign wire_14658 = lut_tile_9_10_chanxy_out[99];
    assign wire_14660 = lut_tile_9_10_chanxy_out[100];
    assign wire_14662 = lut_tile_9_10_chanxy_out[101];
    assign wire_14664 = lut_tile_9_10_chanxy_out[102];
    assign wire_14666 = lut_tile_9_10_chanxy_out[103];
    assign wire_14668 = lut_tile_9_10_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_1_chanxy_in = {wire_10137, wire_10136, wire_11068, wire_9751, wire_9749, wire_9748, wire_9709, wire_9708, wire_9669, wire_9668, wire_9642, wire_1455, wire_10073, wire_10072, wire_11066, wire_9779, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_9650, wire_1455, wire_10127, wire_10126, wire_11064, wire_9777, wire_9743, wire_9742, wire_9703, wire_9702, wire_9663, wire_9662, wire_9658, wire_1455, wire_10065, wire_10064, wire_11062, wire_9775, wire_9741, wire_9740, wire_9701, wire_9700, wire_9666, wire_9661, wire_9660, wire_945, wire_10121, wire_10120, wire_11060, wire_9773, wire_9737, wire_9736, wire_9697, wire_9696, wire_9674, wire_9657, wire_9656, wire_945, wire_10055, wire_10054, wire_11058, wire_9771, wire_9735, wire_9734, wire_9695, wire_9694, wire_9682, wire_9655, wire_9654, wire_945, wire_10113, wire_10112, wire_11056, wire_9769, wire_9733, wire_9732, wire_9693, wire_9692, wire_9690, wire_9653, wire_9652, wire_1459, wire_945, wire_10049, wire_10048, wire_11054, wire_9767, wire_9729, wire_9728, wire_9698, wire_9689, wire_9688, wire_9649, wire_9648, wire_1459, wire_945, wire_10103, wire_10102, wire_11052, wire_9765, wire_9727, wire_9726, wire_9706, wire_9687, wire_9686, wire_9647, wire_9646, wire_1459, wire_945, wire_10041, wire_10040, wire_1459, wire_11050, wire_9763, wire_9725, wire_9724, wire_9714, wire_9685, wire_9684, wire_9645, wire_9644, wire_1459, wire_941, wire_10097, wire_10096, wire_1459, wire_11048, wire_9761, wire_9722, wire_9721, wire_9720, wire_9681, wire_9680, wire_9641, wire_9640, wire_1459, wire_941, wire_10031, wire_10030, wire_1455, wire_11046, wire_9759, wire_9730, wire_9719, wire_9718, wire_9679, wire_9678, wire_9639, wire_9638, wire_1459, wire_941, wire_10089, wire_10088, wire_945, wire_11044, wire_9757, wire_9738, wire_9717, wire_9716, wire_9677, wire_9676, wire_9637, wire_9636, wire_1455, wire_941, wire_10025, wire_10024, wire_945, wire_11042, wire_9755, wire_9746, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632, wire_1455, wire_941, wire_10079, wire_10078, wire_941, wire_11040, wire_9753, wire_9711, wire_9710, wire_9671, wire_9670, wire_9634, wire_9631, wire_9630, wire_1455, wire_941, wire_10153, wire_10074, wire_10167, wire_10130, wire_10125, wire_10124, wire_10165, wire_10122, wire_10149, wire_10058, wire_10053, wire_10052, wire_10147, wire_10050, wire_10161, wire_10106, wire_10101, wire_10100, wire_10159, wire_10098, wire_1459, wire_10143, wire_10034, wire_1455, wire_10029, wire_10028, wire_1455, wire_10141, wire_10026, wire_945, wire_10155, wire_10082, wire_941, wire_10077, wire_10076, wire_941, wire_10135, wire_10134, wire_10129, wire_10128, wire_10069, wire_10068, wire_10063, wire_10062, wire_10057, wire_10056, wire_10117, wire_10116, wire_10111, wire_10110, wire_10105, wire_10104, wire_10045, wire_10044, wire_10039, wire_10038, wire_1459, wire_10033, wire_10032, wire_1455, wire_10093, wire_10092, wire_1455, wire_10087, wire_10086, wire_945, wire_10081, wire_10080, wire_941, wire_10021, wire_10020, wire_941, wire_10169, wire_10138, wire_10133, wire_10132, wire_10071, wire_10070, wire_10151, wire_10066, wire_10061, wire_10060, wire_10119, wire_10118, wire_10163, wire_10114, wire_10109, wire_10108, wire_10047, wire_10046, wire_10145, wire_10042, wire_1459, wire_10037, wire_10036, wire_1459, wire_10095, wire_10094, wire_1455, wire_10157, wire_10090, wire_945, wire_10085, wire_10084, wire_945, wire_10023, wire_10022, wire_941, wire_11166, wire_11144, wire_11122, wire_11098, wire_10169, wire_994, wire_988, wire_979, wire_973, wire_10738, wire_994, wire_10740, wire_994, wire_10770, wire_994, wire_10680, wire_994, wire_11188, wire_11136, wire_11114, wire_11090, wire_10167, wire_994, wire_988, wire_979, wire_973, wire_10710, wire_994, wire_10742, wire_994, wire_10772, wire_991, wire_10682, wire_991, wire_11180, wire_11158, wire_11106, wire_11082, wire_10165, wire_994, wire_988, wire_979, wire_973, wire_10712, wire_991, wire_10744, wire_991, wire_10774, wire_991, wire_10684, wire_991, wire_11172, wire_11150, wire_11128, wire_11074, wire_10163, wire_994, wire_985, wire_979, wire_944, wire_10714, wire_988, wire_10746, wire_988, wire_10776, wire_988, wire_10686, wire_988, wire_11164, wire_11142, wire_11120, wire_11096, wire_10161, wire_994, wire_985, wire_979, wire_944, wire_10716, wire_988, wire_10748, wire_988, wire_10778, wire_985, wire_10688, wire_985, wire_11186, wire_11134, wire_11112, wire_11088, wire_10159, wire_994, wire_985, wire_979, wire_944, wire_10718, wire_985, wire_10750, wire_985, wire_10780, wire_985, wire_10690, wire_985, wire_11178, wire_11156, wire_11104, wire_11080, wire_10157, wire_991, wire_985, wire_976, wire_944, wire_10720, wire_982, wire_10752, wire_982, wire_10782, wire_982, wire_10692, wire_982, wire_11170, wire_11148, wire_11126, wire_11072, wire_10155, wire_991, wire_985, wire_976, wire_944, wire_10722, wire_982, wire_10754, wire_982, wire_10784, wire_979, wire_10694, wire_979, wire_11162, wire_11140, wire_11118, wire_11094, wire_10153, wire_991, wire_985, wire_976, wire_944, wire_10724, wire_979, wire_10756, wire_979, wire_10786, wire_979, wire_10696, wire_979, wire_11184, wire_11132, wire_11110, wire_11086, wire_10151, wire_991, wire_982, wire_976, wire_940, wire_10726, wire_976, wire_10758, wire_976, wire_10788, wire_976, wire_10698, wire_976, wire_11176, wire_11154, wire_11102, wire_11078, wire_10149, wire_991, wire_982, wire_976, wire_940, wire_10728, wire_976, wire_10760, wire_976, wire_10790, wire_973, wire_10700, wire_973, wire_11168, wire_11146, wire_11124, wire_11070, wire_10147, wire_991, wire_982, wire_976, wire_940, wire_10730, wire_973, wire_10762, wire_973, wire_10792, wire_973, wire_10702, wire_973, wire_11160, wire_11138, wire_11116, wire_11092, wire_10145, wire_988, wire_982, wire_973, wire_940, wire_10732, wire_944, wire_10764, wire_944, wire_10794, wire_944, wire_10704, wire_944, wire_11182, wire_11130, wire_11108, wire_11084, wire_10143, wire_988, wire_982, wire_973, wire_940, wire_10734, wire_944, wire_10766, wire_944, wire_10796, wire_940, wire_10706, wire_940, wire_11174, wire_11152, wire_11100, wire_11076, wire_10141, wire_988, wire_982, wire_973, wire_940, wire_10736, wire_940, wire_10768, wire_940, wire_10798, wire_940, wire_10708, wire_940};
    // CHNAXY TOTAL: 558
    assign wire_10020 = lut_tile_10_1_chanxy_out[0];
    assign wire_10022 = lut_tile_10_1_chanxy_out[1];
    assign wire_10024 = lut_tile_10_1_chanxy_out[2];
    assign wire_10026 = lut_tile_10_1_chanxy_out[3];
    assign wire_10027 = lut_tile_10_1_chanxy_out[4];
    assign wire_10028 = lut_tile_10_1_chanxy_out[5];
    assign wire_10030 = lut_tile_10_1_chanxy_out[6];
    assign wire_10032 = lut_tile_10_1_chanxy_out[7];
    assign wire_10034 = lut_tile_10_1_chanxy_out[8];
    assign wire_10035 = lut_tile_10_1_chanxy_out[9];
    assign wire_10036 = lut_tile_10_1_chanxy_out[10];
    assign wire_10038 = lut_tile_10_1_chanxy_out[11];
    assign wire_10040 = lut_tile_10_1_chanxy_out[12];
    assign wire_10042 = lut_tile_10_1_chanxy_out[13];
    assign wire_10043 = lut_tile_10_1_chanxy_out[14];
    assign wire_10044 = lut_tile_10_1_chanxy_out[15];
    assign wire_10046 = lut_tile_10_1_chanxy_out[16];
    assign wire_10048 = lut_tile_10_1_chanxy_out[17];
    assign wire_10050 = lut_tile_10_1_chanxy_out[18];
    assign wire_10051 = lut_tile_10_1_chanxy_out[19];
    assign wire_10052 = lut_tile_10_1_chanxy_out[20];
    assign wire_10054 = lut_tile_10_1_chanxy_out[21];
    assign wire_10056 = lut_tile_10_1_chanxy_out[22];
    assign wire_10058 = lut_tile_10_1_chanxy_out[23];
    assign wire_10059 = lut_tile_10_1_chanxy_out[24];
    assign wire_10060 = lut_tile_10_1_chanxy_out[25];
    assign wire_10062 = lut_tile_10_1_chanxy_out[26];
    assign wire_10064 = lut_tile_10_1_chanxy_out[27];
    assign wire_10066 = lut_tile_10_1_chanxy_out[28];
    assign wire_10067 = lut_tile_10_1_chanxy_out[29];
    assign wire_10068 = lut_tile_10_1_chanxy_out[30];
    assign wire_10070 = lut_tile_10_1_chanxy_out[31];
    assign wire_10072 = lut_tile_10_1_chanxy_out[32];
    assign wire_10074 = lut_tile_10_1_chanxy_out[33];
    assign wire_10075 = lut_tile_10_1_chanxy_out[34];
    assign wire_10076 = lut_tile_10_1_chanxy_out[35];
    assign wire_10078 = lut_tile_10_1_chanxy_out[36];
    assign wire_10080 = lut_tile_10_1_chanxy_out[37];
    assign wire_10082 = lut_tile_10_1_chanxy_out[38];
    assign wire_10083 = lut_tile_10_1_chanxy_out[39];
    assign wire_10084 = lut_tile_10_1_chanxy_out[40];
    assign wire_10086 = lut_tile_10_1_chanxy_out[41];
    assign wire_10088 = lut_tile_10_1_chanxy_out[42];
    assign wire_10090 = lut_tile_10_1_chanxy_out[43];
    assign wire_10091 = lut_tile_10_1_chanxy_out[44];
    assign wire_10092 = lut_tile_10_1_chanxy_out[45];
    assign wire_10094 = lut_tile_10_1_chanxy_out[46];
    assign wire_10096 = lut_tile_10_1_chanxy_out[47];
    assign wire_10098 = lut_tile_10_1_chanxy_out[48];
    assign wire_10099 = lut_tile_10_1_chanxy_out[49];
    assign wire_10100 = lut_tile_10_1_chanxy_out[50];
    assign wire_10102 = lut_tile_10_1_chanxy_out[51];
    assign wire_10104 = lut_tile_10_1_chanxy_out[52];
    assign wire_10106 = lut_tile_10_1_chanxy_out[53];
    assign wire_10107 = lut_tile_10_1_chanxy_out[54];
    assign wire_10108 = lut_tile_10_1_chanxy_out[55];
    assign wire_10110 = lut_tile_10_1_chanxy_out[56];
    assign wire_10112 = lut_tile_10_1_chanxy_out[57];
    assign wire_10114 = lut_tile_10_1_chanxy_out[58];
    assign wire_10115 = lut_tile_10_1_chanxy_out[59];
    assign wire_10116 = lut_tile_10_1_chanxy_out[60];
    assign wire_10118 = lut_tile_10_1_chanxy_out[61];
    assign wire_10120 = lut_tile_10_1_chanxy_out[62];
    assign wire_10122 = lut_tile_10_1_chanxy_out[63];
    assign wire_10123 = lut_tile_10_1_chanxy_out[64];
    assign wire_10124 = lut_tile_10_1_chanxy_out[65];
    assign wire_10126 = lut_tile_10_1_chanxy_out[66];
    assign wire_10128 = lut_tile_10_1_chanxy_out[67];
    assign wire_10130 = lut_tile_10_1_chanxy_out[68];
    assign wire_10131 = lut_tile_10_1_chanxy_out[69];
    assign wire_10132 = lut_tile_10_1_chanxy_out[70];
    assign wire_10134 = lut_tile_10_1_chanxy_out[71];
    assign wire_10136 = lut_tile_10_1_chanxy_out[72];
    assign wire_10138 = lut_tile_10_1_chanxy_out[73];
    assign wire_10139 = lut_tile_10_1_chanxy_out[74];
    assign wire_11071 = lut_tile_10_1_chanxy_out[75];
    assign wire_11073 = lut_tile_10_1_chanxy_out[76];
    assign wire_11075 = lut_tile_10_1_chanxy_out[77];
    assign wire_11077 = lut_tile_10_1_chanxy_out[78];
    assign wire_11079 = lut_tile_10_1_chanxy_out[79];
    assign wire_11081 = lut_tile_10_1_chanxy_out[80];
    assign wire_11083 = lut_tile_10_1_chanxy_out[81];
    assign wire_11085 = lut_tile_10_1_chanxy_out[82];
    assign wire_11087 = lut_tile_10_1_chanxy_out[83];
    assign wire_11089 = lut_tile_10_1_chanxy_out[84];
    assign wire_11091 = lut_tile_10_1_chanxy_out[85];
    assign wire_11093 = lut_tile_10_1_chanxy_out[86];
    assign wire_11095 = lut_tile_10_1_chanxy_out[87];
    assign wire_11097 = lut_tile_10_1_chanxy_out[88];
    assign wire_11099 = lut_tile_10_1_chanxy_out[89];
    assign wire_11101 = lut_tile_10_1_chanxy_out[90];
    assign wire_11103 = lut_tile_10_1_chanxy_out[91];
    assign wire_11105 = lut_tile_10_1_chanxy_out[92];
    assign wire_11107 = lut_tile_10_1_chanxy_out[93];
    assign wire_11109 = lut_tile_10_1_chanxy_out[94];
    assign wire_11111 = lut_tile_10_1_chanxy_out[95];
    assign wire_11113 = lut_tile_10_1_chanxy_out[96];
    assign wire_11115 = lut_tile_10_1_chanxy_out[97];
    assign wire_11117 = lut_tile_10_1_chanxy_out[98];
    assign wire_11119 = lut_tile_10_1_chanxy_out[99];
    assign wire_11121 = lut_tile_10_1_chanxy_out[100];
    assign wire_11123 = lut_tile_10_1_chanxy_out[101];
    assign wire_11125 = lut_tile_10_1_chanxy_out[102];
    assign wire_11127 = lut_tile_10_1_chanxy_out[103];
    assign wire_11129 = lut_tile_10_1_chanxy_out[104];
    assign wire_11131 = lut_tile_10_1_chanxy_out[105];
    assign wire_11133 = lut_tile_10_1_chanxy_out[106];
    assign wire_11135 = lut_tile_10_1_chanxy_out[107];
    assign wire_11137 = lut_tile_10_1_chanxy_out[108];
    assign wire_11139 = lut_tile_10_1_chanxy_out[109];
    assign wire_11141 = lut_tile_10_1_chanxy_out[110];
    assign wire_11143 = lut_tile_10_1_chanxy_out[111];
    assign wire_11145 = lut_tile_10_1_chanxy_out[112];
    assign wire_11147 = lut_tile_10_1_chanxy_out[113];
    assign wire_11149 = lut_tile_10_1_chanxy_out[114];
    assign wire_11151 = lut_tile_10_1_chanxy_out[115];
    assign wire_11153 = lut_tile_10_1_chanxy_out[116];
    assign wire_11155 = lut_tile_10_1_chanxy_out[117];
    assign wire_11157 = lut_tile_10_1_chanxy_out[118];
    assign wire_11159 = lut_tile_10_1_chanxy_out[119];
    assign wire_11160 = lut_tile_10_1_chanxy_out[120];
    assign wire_11161 = lut_tile_10_1_chanxy_out[121];
    assign wire_11162 = lut_tile_10_1_chanxy_out[122];
    assign wire_11163 = lut_tile_10_1_chanxy_out[123];
    assign wire_11164 = lut_tile_10_1_chanxy_out[124];
    assign wire_11165 = lut_tile_10_1_chanxy_out[125];
    assign wire_11166 = lut_tile_10_1_chanxy_out[126];
    assign wire_11167 = lut_tile_10_1_chanxy_out[127];
    assign wire_11168 = lut_tile_10_1_chanxy_out[128];
    assign wire_11169 = lut_tile_10_1_chanxy_out[129];
    assign wire_11170 = lut_tile_10_1_chanxy_out[130];
    assign wire_11171 = lut_tile_10_1_chanxy_out[131];
    assign wire_11172 = lut_tile_10_1_chanxy_out[132];
    assign wire_11173 = lut_tile_10_1_chanxy_out[133];
    assign wire_11174 = lut_tile_10_1_chanxy_out[134];
    assign wire_11175 = lut_tile_10_1_chanxy_out[135];
    assign wire_11176 = lut_tile_10_1_chanxy_out[136];
    assign wire_11177 = lut_tile_10_1_chanxy_out[137];
    assign wire_11178 = lut_tile_10_1_chanxy_out[138];
    assign wire_11179 = lut_tile_10_1_chanxy_out[139];
    assign wire_11180 = lut_tile_10_1_chanxy_out[140];
    assign wire_11181 = lut_tile_10_1_chanxy_out[141];
    assign wire_11182 = lut_tile_10_1_chanxy_out[142];
    assign wire_11183 = lut_tile_10_1_chanxy_out[143];
    assign wire_11184 = lut_tile_10_1_chanxy_out[144];
    assign wire_11185 = lut_tile_10_1_chanxy_out[145];
    assign wire_11186 = lut_tile_10_1_chanxy_out[146];
    assign wire_11187 = lut_tile_10_1_chanxy_out[147];
    assign wire_11188 = lut_tile_10_1_chanxy_out[148];
    assign wire_11189 = lut_tile_10_1_chanxy_out[149];
   // CHANXY OUT
    assign lut_tile_10_2_chanxy_in = {wire_10169, wire_10168, wire_11458, wire_9781, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9644, wire_1971, wire_10199, wire_10132, wire_11456, wire_9809, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_9652, wire_1971, wire_10071, wire_10070, wire_11454, wire_9807, wire_9743, wire_9742, wire_9703, wire_9702, wire_9663, wire_9662, wire_9660, wire_1971, wire_10151, wire_10150, wire_11452, wire_9805, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9668, wire_1461, wire_10181, wire_10060, wire_11450, wire_9803, wire_9737, wire_9736, wire_9697, wire_9696, wire_9676, wire_9657, wire_9656, wire_1461, wire_10119, wire_10118, wire_11448, wire_9801, wire_9735, wire_9734, wire_9695, wire_9694, wire_9684, wire_9655, wire_9654, wire_1461, wire_10163, wire_10162, wire_11446, wire_9799, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9692, wire_1975, wire_1461, wire_10193, wire_10108, wire_11444, wire_9797, wire_9729, wire_9728, wire_9700, wire_9689, wire_9688, wire_9649, wire_9648, wire_1975, wire_1461, wire_10047, wire_10046, wire_11442, wire_9795, wire_9727, wire_9726, wire_9708, wire_9687, wire_9686, wire_9647, wire_9646, wire_1975, wire_1461, wire_10145, wire_10144, wire_1975, wire_11440, wire_9793, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9716, wire_1975, wire_1457, wire_10175, wire_10036, wire_1975, wire_11438, wire_9791, wire_9724, wire_9721, wire_9720, wire_9681, wire_9680, wire_9641, wire_9640, wire_1975, wire_1457, wire_10095, wire_10094, wire_1971, wire_11436, wire_9789, wire_9732, wire_9719, wire_9718, wire_9679, wire_9678, wire_9639, wire_9638, wire_1975, wire_1457, wire_10157, wire_10156, wire_1461, wire_11434, wire_9787, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9740, wire_1971, wire_1457, wire_10187, wire_10084, wire_1461, wire_11432, wire_9785, wire_9748, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632, wire_1971, wire_1457, wire_10023, wire_10022, wire_1457, wire_11430, wire_9783, wire_9711, wire_9710, wire_9671, wire_9670, wire_9636, wire_9631, wire_9630, wire_1971, wire_1457, wire_10137, wire_10136, wire_10073, wire_10072, wire_10127, wire_10126, wire_10065, wire_10064, wire_10121, wire_10120, wire_10055, wire_10054, wire_10113, wire_10112, wire_10049, wire_10048, wire_10103, wire_10102, wire_10041, wire_10040, wire_1975, wire_10097, wire_10096, wire_1975, wire_10031, wire_10030, wire_1971, wire_10089, wire_10088, wire_1461, wire_10025, wire_10024, wire_1461, wire_10079, wire_10078, wire_1457, wire_10153, wire_10152, wire_10167, wire_10166, wire_10197, wire_10124, wire_10165, wire_10164, wire_10149, wire_10148, wire_10179, wire_10052, wire_10147, wire_10146, wire_10161, wire_10160, wire_10191, wire_10100, wire_10159, wire_10158, wire_1975, wire_10143, wire_10142, wire_1971, wire_10173, wire_10028, wire_1971, wire_10141, wire_10140, wire_1461, wire_10155, wire_10154, wire_1457, wire_10185, wire_10076, wire_1457, wire_10135, wire_10134, wire_10129, wire_10128, wire_10183, wire_10068, wire_10063, wire_10062, wire_10057, wire_10056, wire_10195, wire_10116, wire_10111, wire_10110, wire_10105, wire_10104, wire_10177, wire_10044, wire_10039, wire_10038, wire_1975, wire_10033, wire_10032, wire_1971, wire_10189, wire_10092, wire_1971, wire_10087, wire_10086, wire_1461, wire_10081, wire_10080, wire_1457, wire_10171, wire_10020, wire_1457, wire_11166, wire_11144, wire_11122, wire_11098, wire_10138, wire_1510, wire_1504, wire_1495, wire_1489, wire_11188, wire_11136, wire_11114, wire_11090, wire_10130, wire_1510, wire_1504, wire_1495, wire_1489, wire_11180, wire_11158, wire_11106, wire_11082, wire_10122, wire_1510, wire_1504, wire_1495, wire_1489, wire_11172, wire_11150, wire_11128, wire_11074, wire_10114, wire_1510, wire_1501, wire_1495, wire_1460, wire_11164, wire_11142, wire_11120, wire_11096, wire_10106, wire_1510, wire_1501, wire_1495, wire_1460, wire_11186, wire_11134, wire_11112, wire_11088, wire_10098, wire_1510, wire_1501, wire_1495, wire_1460, wire_11178, wire_11156, wire_11104, wire_11080, wire_10090, wire_1507, wire_1501, wire_1492, wire_1460, wire_11170, wire_11148, wire_11126, wire_11072, wire_10082, wire_1507, wire_1501, wire_1492, wire_1460, wire_11162, wire_11140, wire_11118, wire_11094, wire_10074, wire_1507, wire_1501, wire_1492, wire_1460, wire_11184, wire_11132, wire_11110, wire_11086, wire_10066, wire_1507, wire_1498, wire_1492, wire_1456, wire_11176, wire_11154, wire_11102, wire_11078, wire_10058, wire_1507, wire_1498, wire_1492, wire_1456, wire_11168, wire_11146, wire_11124, wire_11070, wire_10050, wire_1507, wire_1498, wire_1492, wire_1456, wire_11160, wire_11138, wire_11116, wire_11092, wire_10042, wire_1504, wire_1498, wire_1489, wire_1456, wire_11182, wire_11130, wire_11108, wire_11084, wire_10034, wire_1504, wire_1498, wire_1489, wire_1456, wire_11174, wire_11152, wire_11100, wire_11076, wire_10026, wire_1504, wire_1498, wire_1489, wire_1456, wire_11578, wire_11526, wire_11504, wire_11482, wire_10199, wire_1510, wire_1504, wire_1495, wire_1489, wire_11570, wire_11548, wire_11496, wire_11474, wire_10197, wire_1510, wire_1504, wire_1495, wire_1489, wire_11562, wire_11540, wire_11518, wire_11466, wire_10195, wire_1510, wire_1504, wire_1495, wire_1489, wire_11554, wire_11532, wire_11510, wire_11488, wire_10193, wire_1510, wire_1501, wire_1495, wire_1460, wire_11576, wire_11524, wire_11502, wire_11480, wire_10191, wire_1510, wire_1501, wire_1495, wire_1460, wire_11568, wire_11546, wire_11494, wire_11472, wire_10189, wire_1510, wire_1501, wire_1495, wire_1460, wire_11560, wire_11538, wire_11516, wire_11464, wire_10187, wire_1507, wire_1501, wire_1492, wire_1460, wire_11552, wire_11530, wire_11508, wire_11486, wire_10185, wire_1507, wire_1501, wire_1492, wire_1460, wire_11574, wire_11522, wire_11500, wire_11478, wire_10183, wire_1507, wire_1501, wire_1492, wire_1460, wire_11566, wire_11544, wire_11492, wire_11470, wire_10181, wire_1507, wire_1498, wire_1492, wire_1456, wire_11558, wire_11536, wire_11514, wire_11462, wire_10179, wire_1507, wire_1498, wire_1492, wire_1456, wire_11550, wire_11528, wire_11506, wire_11484, wire_10177, wire_1507, wire_1498, wire_1492, wire_1456, wire_11572, wire_11520, wire_11498, wire_11476, wire_10175, wire_1504, wire_1498, wire_1489, wire_1456, wire_11564, wire_11542, wire_11490, wire_11468, wire_10173, wire_1504, wire_1498, wire_1489, wire_1456, wire_11556, wire_11534, wire_11512, wire_11460, wire_10171, wire_1504, wire_1498, wire_1489, wire_1456};
    // CHNAXY TOTAL: 573
    assign wire_10021 = lut_tile_10_2_chanxy_out[0];
    assign wire_10029 = lut_tile_10_2_chanxy_out[1];
    assign wire_10037 = lut_tile_10_2_chanxy_out[2];
    assign wire_10045 = lut_tile_10_2_chanxy_out[3];
    assign wire_10053 = lut_tile_10_2_chanxy_out[4];
    assign wire_10061 = lut_tile_10_2_chanxy_out[5];
    assign wire_10069 = lut_tile_10_2_chanxy_out[6];
    assign wire_10077 = lut_tile_10_2_chanxy_out[7];
    assign wire_10085 = lut_tile_10_2_chanxy_out[8];
    assign wire_10093 = lut_tile_10_2_chanxy_out[9];
    assign wire_10101 = lut_tile_10_2_chanxy_out[10];
    assign wire_10109 = lut_tile_10_2_chanxy_out[11];
    assign wire_10117 = lut_tile_10_2_chanxy_out[12];
    assign wire_10125 = lut_tile_10_2_chanxy_out[13];
    assign wire_10133 = lut_tile_10_2_chanxy_out[14];
    assign wire_10140 = lut_tile_10_2_chanxy_out[15];
    assign wire_10142 = lut_tile_10_2_chanxy_out[16];
    assign wire_10144 = lut_tile_10_2_chanxy_out[17];
    assign wire_10146 = lut_tile_10_2_chanxy_out[18];
    assign wire_10148 = lut_tile_10_2_chanxy_out[19];
    assign wire_10150 = lut_tile_10_2_chanxy_out[20];
    assign wire_10152 = lut_tile_10_2_chanxy_out[21];
    assign wire_10154 = lut_tile_10_2_chanxy_out[22];
    assign wire_10156 = lut_tile_10_2_chanxy_out[23];
    assign wire_10158 = lut_tile_10_2_chanxy_out[24];
    assign wire_10160 = lut_tile_10_2_chanxy_out[25];
    assign wire_10162 = lut_tile_10_2_chanxy_out[26];
    assign wire_10164 = lut_tile_10_2_chanxy_out[27];
    assign wire_10166 = lut_tile_10_2_chanxy_out[28];
    assign wire_10168 = lut_tile_10_2_chanxy_out[29];
    assign wire_11461 = lut_tile_10_2_chanxy_out[30];
    assign wire_11463 = lut_tile_10_2_chanxy_out[31];
    assign wire_11465 = lut_tile_10_2_chanxy_out[32];
    assign wire_11467 = lut_tile_10_2_chanxy_out[33];
    assign wire_11469 = lut_tile_10_2_chanxy_out[34];
    assign wire_11471 = lut_tile_10_2_chanxy_out[35];
    assign wire_11473 = lut_tile_10_2_chanxy_out[36];
    assign wire_11475 = lut_tile_10_2_chanxy_out[37];
    assign wire_11477 = lut_tile_10_2_chanxy_out[38];
    assign wire_11479 = lut_tile_10_2_chanxy_out[39];
    assign wire_11481 = lut_tile_10_2_chanxy_out[40];
    assign wire_11483 = lut_tile_10_2_chanxy_out[41];
    assign wire_11485 = lut_tile_10_2_chanxy_out[42];
    assign wire_11487 = lut_tile_10_2_chanxy_out[43];
    assign wire_11489 = lut_tile_10_2_chanxy_out[44];
    assign wire_11491 = lut_tile_10_2_chanxy_out[45];
    assign wire_11493 = lut_tile_10_2_chanxy_out[46];
    assign wire_11495 = lut_tile_10_2_chanxy_out[47];
    assign wire_11497 = lut_tile_10_2_chanxy_out[48];
    assign wire_11499 = lut_tile_10_2_chanxy_out[49];
    assign wire_11501 = lut_tile_10_2_chanxy_out[50];
    assign wire_11503 = lut_tile_10_2_chanxy_out[51];
    assign wire_11505 = lut_tile_10_2_chanxy_out[52];
    assign wire_11507 = lut_tile_10_2_chanxy_out[53];
    assign wire_11509 = lut_tile_10_2_chanxy_out[54];
    assign wire_11511 = lut_tile_10_2_chanxy_out[55];
    assign wire_11513 = lut_tile_10_2_chanxy_out[56];
    assign wire_11515 = lut_tile_10_2_chanxy_out[57];
    assign wire_11517 = lut_tile_10_2_chanxy_out[58];
    assign wire_11519 = lut_tile_10_2_chanxy_out[59];
    assign wire_11521 = lut_tile_10_2_chanxy_out[60];
    assign wire_11523 = lut_tile_10_2_chanxy_out[61];
    assign wire_11525 = lut_tile_10_2_chanxy_out[62];
    assign wire_11527 = lut_tile_10_2_chanxy_out[63];
    assign wire_11529 = lut_tile_10_2_chanxy_out[64];
    assign wire_11531 = lut_tile_10_2_chanxy_out[65];
    assign wire_11533 = lut_tile_10_2_chanxy_out[66];
    assign wire_11535 = lut_tile_10_2_chanxy_out[67];
    assign wire_11537 = lut_tile_10_2_chanxy_out[68];
    assign wire_11539 = lut_tile_10_2_chanxy_out[69];
    assign wire_11541 = lut_tile_10_2_chanxy_out[70];
    assign wire_11543 = lut_tile_10_2_chanxy_out[71];
    assign wire_11545 = lut_tile_10_2_chanxy_out[72];
    assign wire_11547 = lut_tile_10_2_chanxy_out[73];
    assign wire_11549 = lut_tile_10_2_chanxy_out[74];
    assign wire_11550 = lut_tile_10_2_chanxy_out[75];
    assign wire_11551 = lut_tile_10_2_chanxy_out[76];
    assign wire_11552 = lut_tile_10_2_chanxy_out[77];
    assign wire_11553 = lut_tile_10_2_chanxy_out[78];
    assign wire_11554 = lut_tile_10_2_chanxy_out[79];
    assign wire_11555 = lut_tile_10_2_chanxy_out[80];
    assign wire_11556 = lut_tile_10_2_chanxy_out[81];
    assign wire_11557 = lut_tile_10_2_chanxy_out[82];
    assign wire_11558 = lut_tile_10_2_chanxy_out[83];
    assign wire_11559 = lut_tile_10_2_chanxy_out[84];
    assign wire_11560 = lut_tile_10_2_chanxy_out[85];
    assign wire_11561 = lut_tile_10_2_chanxy_out[86];
    assign wire_11562 = lut_tile_10_2_chanxy_out[87];
    assign wire_11563 = lut_tile_10_2_chanxy_out[88];
    assign wire_11564 = lut_tile_10_2_chanxy_out[89];
    assign wire_11565 = lut_tile_10_2_chanxy_out[90];
    assign wire_11566 = lut_tile_10_2_chanxy_out[91];
    assign wire_11567 = lut_tile_10_2_chanxy_out[92];
    assign wire_11568 = lut_tile_10_2_chanxy_out[93];
    assign wire_11569 = lut_tile_10_2_chanxy_out[94];
    assign wire_11570 = lut_tile_10_2_chanxy_out[95];
    assign wire_11571 = lut_tile_10_2_chanxy_out[96];
    assign wire_11572 = lut_tile_10_2_chanxy_out[97];
    assign wire_11573 = lut_tile_10_2_chanxy_out[98];
    assign wire_11574 = lut_tile_10_2_chanxy_out[99];
    assign wire_11575 = lut_tile_10_2_chanxy_out[100];
    assign wire_11576 = lut_tile_10_2_chanxy_out[101];
    assign wire_11577 = lut_tile_10_2_chanxy_out[102];
    assign wire_11578 = lut_tile_10_2_chanxy_out[103];
    assign wire_11579 = lut_tile_10_2_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_3_chanxy_in = {wire_10229, wire_10134, wire_11848, wire_9811, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9638, wire_2487, wire_10129, wire_10128, wire_11846, wire_9839, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9646, wire_2487, wire_10183, wire_10182, wire_11844, wire_9837, wire_9745, wire_9744, wire_9705, wire_9704, wire_9665, wire_9664, wire_9654, wire_2487, wire_10211, wire_10062, wire_11842, wire_9835, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9662, wire_1977, wire_10057, wire_10056, wire_11840, wire_9833, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9670, wire_1977, wire_10195, wire_10194, wire_11838, wire_9831, wire_9737, wire_9736, wire_9697, wire_9696, wire_9678, wire_9657, wire_9656, wire_1977, wire_10223, wire_10110, wire_11836, wire_9829, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9686, wire_2491, wire_1977, wire_10105, wire_10104, wire_11834, wire_9827, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9694, wire_2491, wire_1977, wire_10177, wire_10176, wire_11832, wire_9825, wire_9729, wire_9728, wire_9702, wire_9689, wire_9688, wire_9649, wire_9648, wire_2491, wire_1977, wire_10205, wire_10038, wire_2491, wire_11830, wire_9823, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9710, wire_2491, wire_1973, wire_10033, wire_10032, wire_2487, wire_11828, wire_9821, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9718, wire_2491, wire_1973, wire_10189, wire_10188, wire_2487, wire_11826, wire_9819, wire_9726, wire_9721, wire_9720, wire_9681, wire_9680, wire_9641, wire_9640, wire_2491, wire_1973, wire_10217, wire_10086, wire_1977, wire_11824, wire_9817, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9734, wire_2487, wire_1973, wire_10081, wire_10080, wire_1973, wire_11822, wire_9815, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9742, wire_2487, wire_1973, wire_10171, wire_10170, wire_1973, wire_11820, wire_9813, wire_9713, wire_9712, wire_9673, wire_9672, wire_9633, wire_9632, wire_9630, wire_2487, wire_1973, wire_10169, wire_10168, wire_10199, wire_10198, wire_10213, wire_10070, wire_10151, wire_10150, wire_10181, wire_10180, wire_10225, wire_10118, wire_10163, wire_10162, wire_10193, wire_10192, wire_10207, wire_10046, wire_10145, wire_10144, wire_2491, wire_10175, wire_10174, wire_2491, wire_10219, wire_10094, wire_2487, wire_10157, wire_10156, wire_1977, wire_10187, wire_10186, wire_1977, wire_10201, wire_10022, wire_1973, wire_10137, wire_10136, wire_10073, wire_10072, wire_10227, wire_10126, wire_10065, wire_10064, wire_10121, wire_10120, wire_10209, wire_10054, wire_10113, wire_10112, wire_10049, wire_10048, wire_10221, wire_10102, wire_10041, wire_10040, wire_2491, wire_10097, wire_10096, wire_2491, wire_10203, wire_10030, wire_2487, wire_10089, wire_10088, wire_1977, wire_10025, wire_10024, wire_1977, wire_10215, wire_10078, wire_1973, wire_10153, wire_10152, wire_10167, wire_10166, wire_10197, wire_10196, wire_10165, wire_10164, wire_10149, wire_10148, wire_10179, wire_10178, wire_10147, wire_10146, wire_10161, wire_10160, wire_10191, wire_10190, wire_10159, wire_10158, wire_2491, wire_10143, wire_10142, wire_2487, wire_10173, wire_10172, wire_2487, wire_10141, wire_10140, wire_1977, wire_10155, wire_10154, wire_1973, wire_10185, wire_10184, wire_1973, wire_11578, wire_11526, wire_11504, wire_11482, wire_10132, wire_2026, wire_2020, wire_2011, wire_2005, wire_11570, wire_11548, wire_11496, wire_11474, wire_10124, wire_2026, wire_2020, wire_2011, wire_2005, wire_11562, wire_11540, wire_11518, wire_11466, wire_10116, wire_2026, wire_2020, wire_2011, wire_2005, wire_11554, wire_11532, wire_11510, wire_11488, wire_10108, wire_2026, wire_2017, wire_2011, wire_1976, wire_11576, wire_11524, wire_11502, wire_11480, wire_10100, wire_2026, wire_2017, wire_2011, wire_1976, wire_11568, wire_11546, wire_11494, wire_11472, wire_10092, wire_2026, wire_2017, wire_2011, wire_1976, wire_11560, wire_11538, wire_11516, wire_11464, wire_10084, wire_2023, wire_2017, wire_2008, wire_1976, wire_11552, wire_11530, wire_11508, wire_11486, wire_10076, wire_2023, wire_2017, wire_2008, wire_1976, wire_11574, wire_11522, wire_11500, wire_11478, wire_10068, wire_2023, wire_2017, wire_2008, wire_1976, wire_11566, wire_11544, wire_11492, wire_11470, wire_10060, wire_2023, wire_2014, wire_2008, wire_1972, wire_11558, wire_11536, wire_11514, wire_11462, wire_10052, wire_2023, wire_2014, wire_2008, wire_1972, wire_11550, wire_11528, wire_11506, wire_11484, wire_10044, wire_2023, wire_2014, wire_2008, wire_1972, wire_11572, wire_11520, wire_11498, wire_11476, wire_10036, wire_2020, wire_2014, wire_2005, wire_1972, wire_11564, wire_11542, wire_11490, wire_11468, wire_10028, wire_2020, wire_2014, wire_2005, wire_1972, wire_11556, wire_11534, wire_11512, wire_11460, wire_10020, wire_2020, wire_2014, wire_2005, wire_1972, wire_11962, wire_11938, wire_11886, wire_11864, wire_10229, wire_2026, wire_2020, wire_2011, wire_2005, wire_11954, wire_11930, wire_11908, wire_11856, wire_10227, wire_2026, wire_2020, wire_2011, wire_2005, wire_11946, wire_11922, wire_11900, wire_11878, wire_10225, wire_2026, wire_2020, wire_2011, wire_2005, wire_11968, wire_11914, wire_11892, wire_11870, wire_10223, wire_2026, wire_2017, wire_2011, wire_1976, wire_11960, wire_11936, wire_11884, wire_11862, wire_10221, wire_2026, wire_2017, wire_2011, wire_1976, wire_11952, wire_11928, wire_11906, wire_11854, wire_10219, wire_2026, wire_2017, wire_2011, wire_1976, wire_11944, wire_11920, wire_11898, wire_11876, wire_10217, wire_2023, wire_2017, wire_2008, wire_1976, wire_11966, wire_11912, wire_11890, wire_11868, wire_10215, wire_2023, wire_2017, wire_2008, wire_1976, wire_11958, wire_11934, wire_11882, wire_11860, wire_10213, wire_2023, wire_2017, wire_2008, wire_1976, wire_11950, wire_11926, wire_11904, wire_11852, wire_10211, wire_2023, wire_2014, wire_2008, wire_1972, wire_11942, wire_11918, wire_11896, wire_11874, wire_10209, wire_2023, wire_2014, wire_2008, wire_1972, wire_11964, wire_11910, wire_11888, wire_11866, wire_10207, wire_2023, wire_2014, wire_2008, wire_1972, wire_11956, wire_11932, wire_11880, wire_11858, wire_10205, wire_2020, wire_2014, wire_2005, wire_1972, wire_11948, wire_11924, wire_11902, wire_11850, wire_10203, wire_2020, wire_2014, wire_2005, wire_1972, wire_11940, wire_11916, wire_11894, wire_11872, wire_10201, wire_2020, wire_2014, wire_2005, wire_1972};
    // CHNAXY TOTAL: 573
    assign wire_10023 = lut_tile_10_3_chanxy_out[0];
    assign wire_10031 = lut_tile_10_3_chanxy_out[1];
    assign wire_10039 = lut_tile_10_3_chanxy_out[2];
    assign wire_10047 = lut_tile_10_3_chanxy_out[3];
    assign wire_10055 = lut_tile_10_3_chanxy_out[4];
    assign wire_10063 = lut_tile_10_3_chanxy_out[5];
    assign wire_10071 = lut_tile_10_3_chanxy_out[6];
    assign wire_10079 = lut_tile_10_3_chanxy_out[7];
    assign wire_10087 = lut_tile_10_3_chanxy_out[8];
    assign wire_10095 = lut_tile_10_3_chanxy_out[9];
    assign wire_10103 = lut_tile_10_3_chanxy_out[10];
    assign wire_10111 = lut_tile_10_3_chanxy_out[11];
    assign wire_10119 = lut_tile_10_3_chanxy_out[12];
    assign wire_10127 = lut_tile_10_3_chanxy_out[13];
    assign wire_10135 = lut_tile_10_3_chanxy_out[14];
    assign wire_10170 = lut_tile_10_3_chanxy_out[15];
    assign wire_10172 = lut_tile_10_3_chanxy_out[16];
    assign wire_10174 = lut_tile_10_3_chanxy_out[17];
    assign wire_10176 = lut_tile_10_3_chanxy_out[18];
    assign wire_10178 = lut_tile_10_3_chanxy_out[19];
    assign wire_10180 = lut_tile_10_3_chanxy_out[20];
    assign wire_10182 = lut_tile_10_3_chanxy_out[21];
    assign wire_10184 = lut_tile_10_3_chanxy_out[22];
    assign wire_10186 = lut_tile_10_3_chanxy_out[23];
    assign wire_10188 = lut_tile_10_3_chanxy_out[24];
    assign wire_10190 = lut_tile_10_3_chanxy_out[25];
    assign wire_10192 = lut_tile_10_3_chanxy_out[26];
    assign wire_10194 = lut_tile_10_3_chanxy_out[27];
    assign wire_10196 = lut_tile_10_3_chanxy_out[28];
    assign wire_10198 = lut_tile_10_3_chanxy_out[29];
    assign wire_11851 = lut_tile_10_3_chanxy_out[30];
    assign wire_11853 = lut_tile_10_3_chanxy_out[31];
    assign wire_11855 = lut_tile_10_3_chanxy_out[32];
    assign wire_11857 = lut_tile_10_3_chanxy_out[33];
    assign wire_11859 = lut_tile_10_3_chanxy_out[34];
    assign wire_11861 = lut_tile_10_3_chanxy_out[35];
    assign wire_11863 = lut_tile_10_3_chanxy_out[36];
    assign wire_11865 = lut_tile_10_3_chanxy_out[37];
    assign wire_11867 = lut_tile_10_3_chanxy_out[38];
    assign wire_11869 = lut_tile_10_3_chanxy_out[39];
    assign wire_11871 = lut_tile_10_3_chanxy_out[40];
    assign wire_11873 = lut_tile_10_3_chanxy_out[41];
    assign wire_11875 = lut_tile_10_3_chanxy_out[42];
    assign wire_11877 = lut_tile_10_3_chanxy_out[43];
    assign wire_11879 = lut_tile_10_3_chanxy_out[44];
    assign wire_11881 = lut_tile_10_3_chanxy_out[45];
    assign wire_11883 = lut_tile_10_3_chanxy_out[46];
    assign wire_11885 = lut_tile_10_3_chanxy_out[47];
    assign wire_11887 = lut_tile_10_3_chanxy_out[48];
    assign wire_11889 = lut_tile_10_3_chanxy_out[49];
    assign wire_11891 = lut_tile_10_3_chanxy_out[50];
    assign wire_11893 = lut_tile_10_3_chanxy_out[51];
    assign wire_11895 = lut_tile_10_3_chanxy_out[52];
    assign wire_11897 = lut_tile_10_3_chanxy_out[53];
    assign wire_11899 = lut_tile_10_3_chanxy_out[54];
    assign wire_11901 = lut_tile_10_3_chanxy_out[55];
    assign wire_11903 = lut_tile_10_3_chanxy_out[56];
    assign wire_11905 = lut_tile_10_3_chanxy_out[57];
    assign wire_11907 = lut_tile_10_3_chanxy_out[58];
    assign wire_11909 = lut_tile_10_3_chanxy_out[59];
    assign wire_11911 = lut_tile_10_3_chanxy_out[60];
    assign wire_11913 = lut_tile_10_3_chanxy_out[61];
    assign wire_11915 = lut_tile_10_3_chanxy_out[62];
    assign wire_11917 = lut_tile_10_3_chanxy_out[63];
    assign wire_11919 = lut_tile_10_3_chanxy_out[64];
    assign wire_11921 = lut_tile_10_3_chanxy_out[65];
    assign wire_11923 = lut_tile_10_3_chanxy_out[66];
    assign wire_11925 = lut_tile_10_3_chanxy_out[67];
    assign wire_11927 = lut_tile_10_3_chanxy_out[68];
    assign wire_11929 = lut_tile_10_3_chanxy_out[69];
    assign wire_11931 = lut_tile_10_3_chanxy_out[70];
    assign wire_11933 = lut_tile_10_3_chanxy_out[71];
    assign wire_11935 = lut_tile_10_3_chanxy_out[72];
    assign wire_11937 = lut_tile_10_3_chanxy_out[73];
    assign wire_11939 = lut_tile_10_3_chanxy_out[74];
    assign wire_11940 = lut_tile_10_3_chanxy_out[75];
    assign wire_11941 = lut_tile_10_3_chanxy_out[76];
    assign wire_11942 = lut_tile_10_3_chanxy_out[77];
    assign wire_11943 = lut_tile_10_3_chanxy_out[78];
    assign wire_11944 = lut_tile_10_3_chanxy_out[79];
    assign wire_11945 = lut_tile_10_3_chanxy_out[80];
    assign wire_11946 = lut_tile_10_3_chanxy_out[81];
    assign wire_11947 = lut_tile_10_3_chanxy_out[82];
    assign wire_11948 = lut_tile_10_3_chanxy_out[83];
    assign wire_11949 = lut_tile_10_3_chanxy_out[84];
    assign wire_11950 = lut_tile_10_3_chanxy_out[85];
    assign wire_11951 = lut_tile_10_3_chanxy_out[86];
    assign wire_11952 = lut_tile_10_3_chanxy_out[87];
    assign wire_11953 = lut_tile_10_3_chanxy_out[88];
    assign wire_11954 = lut_tile_10_3_chanxy_out[89];
    assign wire_11955 = lut_tile_10_3_chanxy_out[90];
    assign wire_11956 = lut_tile_10_3_chanxy_out[91];
    assign wire_11957 = lut_tile_10_3_chanxy_out[92];
    assign wire_11958 = lut_tile_10_3_chanxy_out[93];
    assign wire_11959 = lut_tile_10_3_chanxy_out[94];
    assign wire_11960 = lut_tile_10_3_chanxy_out[95];
    assign wire_11961 = lut_tile_10_3_chanxy_out[96];
    assign wire_11962 = lut_tile_10_3_chanxy_out[97];
    assign wire_11963 = lut_tile_10_3_chanxy_out[98];
    assign wire_11964 = lut_tile_10_3_chanxy_out[99];
    assign wire_11965 = lut_tile_10_3_chanxy_out[100];
    assign wire_11966 = lut_tile_10_3_chanxy_out[101];
    assign wire_11967 = lut_tile_10_3_chanxy_out[102];
    assign wire_11968 = lut_tile_10_3_chanxy_out[103];
    assign wire_11969 = lut_tile_10_3_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_4_chanxy_in = {wire_10153, wire_10152, wire_12238, wire_9841, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9640, wire_3003, wire_10167, wire_10166, wire_12236, wire_9869, wire_9779, wire_9778, wire_9769, wire_9768, wire_9759, wire_9758, wire_9648, wire_3003, wire_10197, wire_10196, wire_12234, wire_9867, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9656, wire_3003, wire_10165, wire_10164, wire_12232, wire_9865, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9664, wire_2493, wire_10149, wire_10148, wire_12230, wire_9863, wire_9777, wire_9776, wire_9767, wire_9766, wire_9757, wire_9756, wire_9672, wire_2493, wire_10179, wire_10178, wire_12228, wire_9861, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9680, wire_2493, wire_10147, wire_10146, wire_12226, wire_9859, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9688, wire_3007, wire_2493, wire_10161, wire_10160, wire_12224, wire_9857, wire_9775, wire_9774, wire_9765, wire_9764, wire_9755, wire_9754, wire_9696, wire_3007, wire_2493, wire_10191, wire_10190, wire_12222, wire_9855, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9704, wire_3007, wire_2493, wire_10159, wire_10158, wire_3007, wire_12220, wire_9853, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9712, wire_3007, wire_2489, wire_10143, wire_10142, wire_3003, wire_12218, wire_9851, wire_9773, wire_9772, wire_9763, wire_9762, wire_9753, wire_9752, wire_9720, wire_3007, wire_2489, wire_10173, wire_10172, wire_3003, wire_12216, wire_9849, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9728, wire_3007, wire_2489, wire_10141, wire_10140, wire_2493, wire_12214, wire_9847, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9736, wire_3003, wire_2489, wire_10155, wire_10154, wire_2489, wire_12212, wire_9845, wire_9771, wire_9770, wire_9761, wire_9760, wire_9751, wire_9750, wire_9744, wire_3003, wire_2489, wire_10185, wire_10184, wire_2489, wire_12210, wire_9843, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9632, wire_3003, wire_2489, wire_10229, wire_10228, wire_10257, wire_10128, wire_10183, wire_10182, wire_10211, wire_10210, wire_10239, wire_10056, wire_10195, wire_10194, wire_10223, wire_10222, wire_10251, wire_10104, wire_10177, wire_10176, wire_10205, wire_10204, wire_3007, wire_10233, wire_10032, wire_3003, wire_10189, wire_10188, wire_3003, wire_10217, wire_10216, wire_2493, wire_10245, wire_10080, wire_2489, wire_10171, wire_10170, wire_2489, wire_10169, wire_10168, wire_10199, wire_10198, wire_10213, wire_10212, wire_10151, wire_10150, wire_10181, wire_10180, wire_10225, wire_10224, wire_10163, wire_10162, wire_10193, wire_10192, wire_10207, wire_10206, wire_10145, wire_10144, wire_3007, wire_10175, wire_10174, wire_3007, wire_10219, wire_10218, wire_3003, wire_10157, wire_10156, wire_2493, wire_10187, wire_10186, wire_2493, wire_10201, wire_10200, wire_2489, wire_10259, wire_10136, wire_10243, wire_10072, wire_10227, wire_10226, wire_10241, wire_10064, wire_10255, wire_10120, wire_10209, wire_10208, wire_10253, wire_10112, wire_10237, wire_10048, wire_10221, wire_10220, wire_10235, wire_10040, wire_3007, wire_10249, wire_10096, wire_3007, wire_10203, wire_10202, wire_3003, wire_10247, wire_10088, wire_2493, wire_10231, wire_10024, wire_2493, wire_10215, wire_10214, wire_2489, wire_11962, wire_11938, wire_11886, wire_11864, wire_10134, wire_2542, wire_2536, wire_2527, wire_2521, wire_11954, wire_11930, wire_11908, wire_11856, wire_10126, wire_2542, wire_2536, wire_2527, wire_2521, wire_11946, wire_11922, wire_11900, wire_11878, wire_10118, wire_2542, wire_2536, wire_2527, wire_2521, wire_11968, wire_11914, wire_11892, wire_11870, wire_10110, wire_2542, wire_2533, wire_2527, wire_2492, wire_11960, wire_11936, wire_11884, wire_11862, wire_10102, wire_2542, wire_2533, wire_2527, wire_2492, wire_11952, wire_11928, wire_11906, wire_11854, wire_10094, wire_2542, wire_2533, wire_2527, wire_2492, wire_11944, wire_11920, wire_11898, wire_11876, wire_10086, wire_2539, wire_2533, wire_2524, wire_2492, wire_11966, wire_11912, wire_11890, wire_11868, wire_10078, wire_2539, wire_2533, wire_2524, wire_2492, wire_11958, wire_11934, wire_11882, wire_11860, wire_10070, wire_2539, wire_2533, wire_2524, wire_2492, wire_11950, wire_11926, wire_11904, wire_11852, wire_10062, wire_2539, wire_2530, wire_2524, wire_2488, wire_11942, wire_11918, wire_11896, wire_11874, wire_10054, wire_2539, wire_2530, wire_2524, wire_2488, wire_11964, wire_11910, wire_11888, wire_11866, wire_10046, wire_2539, wire_2530, wire_2524, wire_2488, wire_11956, wire_11932, wire_11880, wire_11858, wire_10038, wire_2536, wire_2530, wire_2521, wire_2488, wire_11948, wire_11924, wire_11902, wire_11850, wire_10030, wire_2536, wire_2530, wire_2521, wire_2488, wire_11940, wire_11916, wire_11894, wire_11872, wire_10022, wire_2536, wire_2530, wire_2521, wire_2488, wire_12344, wire_12322, wire_12298, wire_12246, wire_10259, wire_2542, wire_2536, wire_2527, wire_2521, wire_12336, wire_12314, wire_12290, wire_12268, wire_10257, wire_2542, wire_2536, wire_2527, wire_2521, wire_12358, wire_12306, wire_12282, wire_12260, wire_10255, wire_2542, wire_2536, wire_2527, wire_2521, wire_12350, wire_12328, wire_12274, wire_12252, wire_10253, wire_2542, wire_2533, wire_2527, wire_2492, wire_12342, wire_12320, wire_12296, wire_12244, wire_10251, wire_2542, wire_2533, wire_2527, wire_2492, wire_12334, wire_12312, wire_12288, wire_12266, wire_10249, wire_2542, wire_2533, wire_2527, wire_2492, wire_12356, wire_12304, wire_12280, wire_12258, wire_10247, wire_2539, wire_2533, wire_2524, wire_2492, wire_12348, wire_12326, wire_12272, wire_12250, wire_10245, wire_2539, wire_2533, wire_2524, wire_2492, wire_12340, wire_12318, wire_12294, wire_12242, wire_10243, wire_2539, wire_2533, wire_2524, wire_2492, wire_12332, wire_12310, wire_12286, wire_12264, wire_10241, wire_2539, wire_2530, wire_2524, wire_2488, wire_12354, wire_12302, wire_12278, wire_12256, wire_10239, wire_2539, wire_2530, wire_2524, wire_2488, wire_12346, wire_12324, wire_12270, wire_12248, wire_10237, wire_2539, wire_2530, wire_2524, wire_2488, wire_12338, wire_12316, wire_12292, wire_12240, wire_10235, wire_2536, wire_2530, wire_2521, wire_2488, wire_12330, wire_12308, wire_12284, wire_12262, wire_10233, wire_2536, wire_2530, wire_2521, wire_2488, wire_12352, wire_12300, wire_12276, wire_12254, wire_10231, wire_2536, wire_2530, wire_2521, wire_2488};
    // CHNAXY TOTAL: 573
    assign wire_10025 = lut_tile_10_4_chanxy_out[0];
    assign wire_10033 = lut_tile_10_4_chanxy_out[1];
    assign wire_10041 = lut_tile_10_4_chanxy_out[2];
    assign wire_10049 = lut_tile_10_4_chanxy_out[3];
    assign wire_10057 = lut_tile_10_4_chanxy_out[4];
    assign wire_10065 = lut_tile_10_4_chanxy_out[5];
    assign wire_10073 = lut_tile_10_4_chanxy_out[6];
    assign wire_10081 = lut_tile_10_4_chanxy_out[7];
    assign wire_10089 = lut_tile_10_4_chanxy_out[8];
    assign wire_10097 = lut_tile_10_4_chanxy_out[9];
    assign wire_10105 = lut_tile_10_4_chanxy_out[10];
    assign wire_10113 = lut_tile_10_4_chanxy_out[11];
    assign wire_10121 = lut_tile_10_4_chanxy_out[12];
    assign wire_10129 = lut_tile_10_4_chanxy_out[13];
    assign wire_10137 = lut_tile_10_4_chanxy_out[14];
    assign wire_10200 = lut_tile_10_4_chanxy_out[15];
    assign wire_10202 = lut_tile_10_4_chanxy_out[16];
    assign wire_10204 = lut_tile_10_4_chanxy_out[17];
    assign wire_10206 = lut_tile_10_4_chanxy_out[18];
    assign wire_10208 = lut_tile_10_4_chanxy_out[19];
    assign wire_10210 = lut_tile_10_4_chanxy_out[20];
    assign wire_10212 = lut_tile_10_4_chanxy_out[21];
    assign wire_10214 = lut_tile_10_4_chanxy_out[22];
    assign wire_10216 = lut_tile_10_4_chanxy_out[23];
    assign wire_10218 = lut_tile_10_4_chanxy_out[24];
    assign wire_10220 = lut_tile_10_4_chanxy_out[25];
    assign wire_10222 = lut_tile_10_4_chanxy_out[26];
    assign wire_10224 = lut_tile_10_4_chanxy_out[27];
    assign wire_10226 = lut_tile_10_4_chanxy_out[28];
    assign wire_10228 = lut_tile_10_4_chanxy_out[29];
    assign wire_12241 = lut_tile_10_4_chanxy_out[30];
    assign wire_12243 = lut_tile_10_4_chanxy_out[31];
    assign wire_12245 = lut_tile_10_4_chanxy_out[32];
    assign wire_12247 = lut_tile_10_4_chanxy_out[33];
    assign wire_12249 = lut_tile_10_4_chanxy_out[34];
    assign wire_12251 = lut_tile_10_4_chanxy_out[35];
    assign wire_12253 = lut_tile_10_4_chanxy_out[36];
    assign wire_12255 = lut_tile_10_4_chanxy_out[37];
    assign wire_12257 = lut_tile_10_4_chanxy_out[38];
    assign wire_12259 = lut_tile_10_4_chanxy_out[39];
    assign wire_12261 = lut_tile_10_4_chanxy_out[40];
    assign wire_12263 = lut_tile_10_4_chanxy_out[41];
    assign wire_12265 = lut_tile_10_4_chanxy_out[42];
    assign wire_12267 = lut_tile_10_4_chanxy_out[43];
    assign wire_12269 = lut_tile_10_4_chanxy_out[44];
    assign wire_12271 = lut_tile_10_4_chanxy_out[45];
    assign wire_12273 = lut_tile_10_4_chanxy_out[46];
    assign wire_12275 = lut_tile_10_4_chanxy_out[47];
    assign wire_12277 = lut_tile_10_4_chanxy_out[48];
    assign wire_12279 = lut_tile_10_4_chanxy_out[49];
    assign wire_12281 = lut_tile_10_4_chanxy_out[50];
    assign wire_12283 = lut_tile_10_4_chanxy_out[51];
    assign wire_12285 = lut_tile_10_4_chanxy_out[52];
    assign wire_12287 = lut_tile_10_4_chanxy_out[53];
    assign wire_12289 = lut_tile_10_4_chanxy_out[54];
    assign wire_12291 = lut_tile_10_4_chanxy_out[55];
    assign wire_12293 = lut_tile_10_4_chanxy_out[56];
    assign wire_12295 = lut_tile_10_4_chanxy_out[57];
    assign wire_12297 = lut_tile_10_4_chanxy_out[58];
    assign wire_12299 = lut_tile_10_4_chanxy_out[59];
    assign wire_12301 = lut_tile_10_4_chanxy_out[60];
    assign wire_12303 = lut_tile_10_4_chanxy_out[61];
    assign wire_12305 = lut_tile_10_4_chanxy_out[62];
    assign wire_12307 = lut_tile_10_4_chanxy_out[63];
    assign wire_12309 = lut_tile_10_4_chanxy_out[64];
    assign wire_12311 = lut_tile_10_4_chanxy_out[65];
    assign wire_12313 = lut_tile_10_4_chanxy_out[66];
    assign wire_12315 = lut_tile_10_4_chanxy_out[67];
    assign wire_12317 = lut_tile_10_4_chanxy_out[68];
    assign wire_12319 = lut_tile_10_4_chanxy_out[69];
    assign wire_12321 = lut_tile_10_4_chanxy_out[70];
    assign wire_12323 = lut_tile_10_4_chanxy_out[71];
    assign wire_12325 = lut_tile_10_4_chanxy_out[72];
    assign wire_12327 = lut_tile_10_4_chanxy_out[73];
    assign wire_12329 = lut_tile_10_4_chanxy_out[74];
    assign wire_12330 = lut_tile_10_4_chanxy_out[75];
    assign wire_12331 = lut_tile_10_4_chanxy_out[76];
    assign wire_12332 = lut_tile_10_4_chanxy_out[77];
    assign wire_12333 = lut_tile_10_4_chanxy_out[78];
    assign wire_12334 = lut_tile_10_4_chanxy_out[79];
    assign wire_12335 = lut_tile_10_4_chanxy_out[80];
    assign wire_12336 = lut_tile_10_4_chanxy_out[81];
    assign wire_12337 = lut_tile_10_4_chanxy_out[82];
    assign wire_12338 = lut_tile_10_4_chanxy_out[83];
    assign wire_12339 = lut_tile_10_4_chanxy_out[84];
    assign wire_12340 = lut_tile_10_4_chanxy_out[85];
    assign wire_12341 = lut_tile_10_4_chanxy_out[86];
    assign wire_12342 = lut_tile_10_4_chanxy_out[87];
    assign wire_12343 = lut_tile_10_4_chanxy_out[88];
    assign wire_12344 = lut_tile_10_4_chanxy_out[89];
    assign wire_12345 = lut_tile_10_4_chanxy_out[90];
    assign wire_12346 = lut_tile_10_4_chanxy_out[91];
    assign wire_12347 = lut_tile_10_4_chanxy_out[92];
    assign wire_12348 = lut_tile_10_4_chanxy_out[93];
    assign wire_12349 = lut_tile_10_4_chanxy_out[94];
    assign wire_12350 = lut_tile_10_4_chanxy_out[95];
    assign wire_12351 = lut_tile_10_4_chanxy_out[96];
    assign wire_12352 = lut_tile_10_4_chanxy_out[97];
    assign wire_12353 = lut_tile_10_4_chanxy_out[98];
    assign wire_12354 = lut_tile_10_4_chanxy_out[99];
    assign wire_12355 = lut_tile_10_4_chanxy_out[100];
    assign wire_12356 = lut_tile_10_4_chanxy_out[101];
    assign wire_12357 = lut_tile_10_4_chanxy_out[102];
    assign wire_12358 = lut_tile_10_4_chanxy_out[103];
    assign wire_12359 = lut_tile_10_4_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_5_chanxy_in = {wire_10259, wire_10258, wire_12628, wire_9871, wire_9809, wire_9808, wire_9799, wire_9798, wire_9789, wire_9788, wire_9752, wire_3519, wire_10243, wire_10242, wire_12626, wire_9899, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9754, wire_3519, wire_10227, wire_10226, wire_12624, wire_9897, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9756, wire_3519, wire_10241, wire_10240, wire_12622, wire_9895, wire_9807, wire_9806, wire_9797, wire_9796, wire_9787, wire_9786, wire_9758, wire_3009, wire_10255, wire_10254, wire_12620, wire_9893, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9760, wire_3009, wire_10209, wire_10208, wire_12618, wire_9891, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9762, wire_3009, wire_10253, wire_10252, wire_12616, wire_9889, wire_9805, wire_9804, wire_9795, wire_9794, wire_9785, wire_9784, wire_9764, wire_3523, wire_3009, wire_10237, wire_10236, wire_12614, wire_9887, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9766, wire_3523, wire_3009, wire_10221, wire_10220, wire_12612, wire_9885, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9768, wire_3523, wire_3009, wire_10235, wire_10234, wire_3523, wire_12610, wire_9883, wire_9803, wire_9802, wire_9793, wire_9792, wire_9783, wire_9782, wire_9770, wire_3523, wire_3005, wire_10249, wire_10248, wire_3523, wire_12608, wire_9881, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9772, wire_3523, wire_3005, wire_10203, wire_10202, wire_3519, wire_12606, wire_9879, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9774, wire_3523, wire_3005, wire_10247, wire_10246, wire_3009, wire_12604, wire_9877, wire_9801, wire_9800, wire_9791, wire_9790, wire_9781, wire_9780, wire_9776, wire_3519, wire_3005, wire_10231, wire_10230, wire_3009, wire_12602, wire_9875, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9778, wire_3519, wire_3005, wire_10215, wire_10214, wire_3005, wire_12600, wire_9873, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9750, wire_3519, wire_3005, wire_10273, wire_10152, wire_10287, wire_10166, wire_10197, wire_10196, wire_10285, wire_10164, wire_10269, wire_10148, wire_10179, wire_10178, wire_10267, wire_10146, wire_10281, wire_10160, wire_10191, wire_10190, wire_10279, wire_10158, wire_3523, wire_10263, wire_10142, wire_3519, wire_10173, wire_10172, wire_3519, wire_10261, wire_10140, wire_3009, wire_10275, wire_10154, wire_3005, wire_10185, wire_10184, wire_3005, wire_10229, wire_10228, wire_10257, wire_10256, wire_10183, wire_10182, wire_10211, wire_10210, wire_10239, wire_10238, wire_10195, wire_10194, wire_10223, wire_10222, wire_10251, wire_10250, wire_10177, wire_10176, wire_10205, wire_10204, wire_3523, wire_10233, wire_10232, wire_3519, wire_10189, wire_10188, wire_3519, wire_10217, wire_10216, wire_3009, wire_10245, wire_10244, wire_3005, wire_10171, wire_10170, wire_3005, wire_10289, wire_10168, wire_10199, wire_10198, wire_10213, wire_10212, wire_10271, wire_10150, wire_10181, wire_10180, wire_10225, wire_10224, wire_10283, wire_10162, wire_10193, wire_10192, wire_10207, wire_10206, wire_10265, wire_10144, wire_3523, wire_10175, wire_10174, wire_3523, wire_10219, wire_10218, wire_3519, wire_10277, wire_10156, wire_3009, wire_10187, wire_10186, wire_3009, wire_10201, wire_10200, wire_3005, wire_12344, wire_12322, wire_12298, wire_12246, wire_10136, wire_3058, wire_3052, wire_3043, wire_3037, wire_12336, wire_12314, wire_12290, wire_12268, wire_10128, wire_3058, wire_3052, wire_3043, wire_3037, wire_12358, wire_12306, wire_12282, wire_12260, wire_10120, wire_3058, wire_3052, wire_3043, wire_3037, wire_12350, wire_12328, wire_12274, wire_12252, wire_10112, wire_3058, wire_3049, wire_3043, wire_3008, wire_12342, wire_12320, wire_12296, wire_12244, wire_10104, wire_3058, wire_3049, wire_3043, wire_3008, wire_12334, wire_12312, wire_12288, wire_12266, wire_10096, wire_3058, wire_3049, wire_3043, wire_3008, wire_12356, wire_12304, wire_12280, wire_12258, wire_10088, wire_3055, wire_3049, wire_3040, wire_3008, wire_12348, wire_12326, wire_12272, wire_12250, wire_10080, wire_3055, wire_3049, wire_3040, wire_3008, wire_12340, wire_12318, wire_12294, wire_12242, wire_10072, wire_3055, wire_3049, wire_3040, wire_3008, wire_12332, wire_12310, wire_12286, wire_12264, wire_10064, wire_3055, wire_3046, wire_3040, wire_3004, wire_12354, wire_12302, wire_12278, wire_12256, wire_10056, wire_3055, wire_3046, wire_3040, wire_3004, wire_12346, wire_12324, wire_12270, wire_12248, wire_10048, wire_3055, wire_3046, wire_3040, wire_3004, wire_12338, wire_12316, wire_12292, wire_12240, wire_10040, wire_3052, wire_3046, wire_3037, wire_3004, wire_12330, wire_12308, wire_12284, wire_12262, wire_10032, wire_3052, wire_3046, wire_3037, wire_3004, wire_12352, wire_12300, wire_12276, wire_12254, wire_10024, wire_3052, wire_3046, wire_3037, wire_3004, wire_12726, wire_12704, wire_12682, wire_12658, wire_10289, wire_3058, wire_3052, wire_3043, wire_3037, wire_12748, wire_12696, wire_12674, wire_12650, wire_10287, wire_3058, wire_3052, wire_3043, wire_3037, wire_12740, wire_12718, wire_12666, wire_12642, wire_10285, wire_3058, wire_3052, wire_3043, wire_3037, wire_12732, wire_12710, wire_12688, wire_12634, wire_10283, wire_3058, wire_3049, wire_3043, wire_3008, wire_12724, wire_12702, wire_12680, wire_12656, wire_10281, wire_3058, wire_3049, wire_3043, wire_3008, wire_12746, wire_12694, wire_12672, wire_12648, wire_10279, wire_3058, wire_3049, wire_3043, wire_3008, wire_12738, wire_12716, wire_12664, wire_12640, wire_10277, wire_3055, wire_3049, wire_3040, wire_3008, wire_12730, wire_12708, wire_12686, wire_12632, wire_10275, wire_3055, wire_3049, wire_3040, wire_3008, wire_12722, wire_12700, wire_12678, wire_12654, wire_10273, wire_3055, wire_3049, wire_3040, wire_3008, wire_12744, wire_12692, wire_12670, wire_12646, wire_10271, wire_3055, wire_3046, wire_3040, wire_3004, wire_12736, wire_12714, wire_12662, wire_12638, wire_10269, wire_3055, wire_3046, wire_3040, wire_3004, wire_12728, wire_12706, wire_12684, wire_12630, wire_10267, wire_3055, wire_3046, wire_3040, wire_3004, wire_12720, wire_12698, wire_12676, wire_12652, wire_10265, wire_3052, wire_3046, wire_3037, wire_3004, wire_12742, wire_12690, wire_12668, wire_12644, wire_10263, wire_3052, wire_3046, wire_3037, wire_3004, wire_12734, wire_12712, wire_12660, wire_12636, wire_10261, wire_3052, wire_3046, wire_3037, wire_3004};
    // CHNAXY TOTAL: 573
    assign wire_10141 = lut_tile_10_5_chanxy_out[0];
    assign wire_10143 = lut_tile_10_5_chanxy_out[1];
    assign wire_10145 = lut_tile_10_5_chanxy_out[2];
    assign wire_10147 = lut_tile_10_5_chanxy_out[3];
    assign wire_10149 = lut_tile_10_5_chanxy_out[4];
    assign wire_10151 = lut_tile_10_5_chanxy_out[5];
    assign wire_10153 = lut_tile_10_5_chanxy_out[6];
    assign wire_10155 = lut_tile_10_5_chanxy_out[7];
    assign wire_10157 = lut_tile_10_5_chanxy_out[8];
    assign wire_10159 = lut_tile_10_5_chanxy_out[9];
    assign wire_10161 = lut_tile_10_5_chanxy_out[10];
    assign wire_10163 = lut_tile_10_5_chanxy_out[11];
    assign wire_10165 = lut_tile_10_5_chanxy_out[12];
    assign wire_10167 = lut_tile_10_5_chanxy_out[13];
    assign wire_10169 = lut_tile_10_5_chanxy_out[14];
    assign wire_10230 = lut_tile_10_5_chanxy_out[15];
    assign wire_10232 = lut_tile_10_5_chanxy_out[16];
    assign wire_10234 = lut_tile_10_5_chanxy_out[17];
    assign wire_10236 = lut_tile_10_5_chanxy_out[18];
    assign wire_10238 = lut_tile_10_5_chanxy_out[19];
    assign wire_10240 = lut_tile_10_5_chanxy_out[20];
    assign wire_10242 = lut_tile_10_5_chanxy_out[21];
    assign wire_10244 = lut_tile_10_5_chanxy_out[22];
    assign wire_10246 = lut_tile_10_5_chanxy_out[23];
    assign wire_10248 = lut_tile_10_5_chanxy_out[24];
    assign wire_10250 = lut_tile_10_5_chanxy_out[25];
    assign wire_10252 = lut_tile_10_5_chanxy_out[26];
    assign wire_10254 = lut_tile_10_5_chanxy_out[27];
    assign wire_10256 = lut_tile_10_5_chanxy_out[28];
    assign wire_10258 = lut_tile_10_5_chanxy_out[29];
    assign wire_12631 = lut_tile_10_5_chanxy_out[30];
    assign wire_12633 = lut_tile_10_5_chanxy_out[31];
    assign wire_12635 = lut_tile_10_5_chanxy_out[32];
    assign wire_12637 = lut_tile_10_5_chanxy_out[33];
    assign wire_12639 = lut_tile_10_5_chanxy_out[34];
    assign wire_12641 = lut_tile_10_5_chanxy_out[35];
    assign wire_12643 = lut_tile_10_5_chanxy_out[36];
    assign wire_12645 = lut_tile_10_5_chanxy_out[37];
    assign wire_12647 = lut_tile_10_5_chanxy_out[38];
    assign wire_12649 = lut_tile_10_5_chanxy_out[39];
    assign wire_12651 = lut_tile_10_5_chanxy_out[40];
    assign wire_12653 = lut_tile_10_5_chanxy_out[41];
    assign wire_12655 = lut_tile_10_5_chanxy_out[42];
    assign wire_12657 = lut_tile_10_5_chanxy_out[43];
    assign wire_12659 = lut_tile_10_5_chanxy_out[44];
    assign wire_12661 = lut_tile_10_5_chanxy_out[45];
    assign wire_12663 = lut_tile_10_5_chanxy_out[46];
    assign wire_12665 = lut_tile_10_5_chanxy_out[47];
    assign wire_12667 = lut_tile_10_5_chanxy_out[48];
    assign wire_12669 = lut_tile_10_5_chanxy_out[49];
    assign wire_12671 = lut_tile_10_5_chanxy_out[50];
    assign wire_12673 = lut_tile_10_5_chanxy_out[51];
    assign wire_12675 = lut_tile_10_5_chanxy_out[52];
    assign wire_12677 = lut_tile_10_5_chanxy_out[53];
    assign wire_12679 = lut_tile_10_5_chanxy_out[54];
    assign wire_12681 = lut_tile_10_5_chanxy_out[55];
    assign wire_12683 = lut_tile_10_5_chanxy_out[56];
    assign wire_12685 = lut_tile_10_5_chanxy_out[57];
    assign wire_12687 = lut_tile_10_5_chanxy_out[58];
    assign wire_12689 = lut_tile_10_5_chanxy_out[59];
    assign wire_12691 = lut_tile_10_5_chanxy_out[60];
    assign wire_12693 = lut_tile_10_5_chanxy_out[61];
    assign wire_12695 = lut_tile_10_5_chanxy_out[62];
    assign wire_12697 = lut_tile_10_5_chanxy_out[63];
    assign wire_12699 = lut_tile_10_5_chanxy_out[64];
    assign wire_12701 = lut_tile_10_5_chanxy_out[65];
    assign wire_12703 = lut_tile_10_5_chanxy_out[66];
    assign wire_12705 = lut_tile_10_5_chanxy_out[67];
    assign wire_12707 = lut_tile_10_5_chanxy_out[68];
    assign wire_12709 = lut_tile_10_5_chanxy_out[69];
    assign wire_12711 = lut_tile_10_5_chanxy_out[70];
    assign wire_12713 = lut_tile_10_5_chanxy_out[71];
    assign wire_12715 = lut_tile_10_5_chanxy_out[72];
    assign wire_12717 = lut_tile_10_5_chanxy_out[73];
    assign wire_12719 = lut_tile_10_5_chanxy_out[74];
    assign wire_12720 = lut_tile_10_5_chanxy_out[75];
    assign wire_12721 = lut_tile_10_5_chanxy_out[76];
    assign wire_12722 = lut_tile_10_5_chanxy_out[77];
    assign wire_12723 = lut_tile_10_5_chanxy_out[78];
    assign wire_12724 = lut_tile_10_5_chanxy_out[79];
    assign wire_12725 = lut_tile_10_5_chanxy_out[80];
    assign wire_12726 = lut_tile_10_5_chanxy_out[81];
    assign wire_12727 = lut_tile_10_5_chanxy_out[82];
    assign wire_12728 = lut_tile_10_5_chanxy_out[83];
    assign wire_12729 = lut_tile_10_5_chanxy_out[84];
    assign wire_12730 = lut_tile_10_5_chanxy_out[85];
    assign wire_12731 = lut_tile_10_5_chanxy_out[86];
    assign wire_12732 = lut_tile_10_5_chanxy_out[87];
    assign wire_12733 = lut_tile_10_5_chanxy_out[88];
    assign wire_12734 = lut_tile_10_5_chanxy_out[89];
    assign wire_12735 = lut_tile_10_5_chanxy_out[90];
    assign wire_12736 = lut_tile_10_5_chanxy_out[91];
    assign wire_12737 = lut_tile_10_5_chanxy_out[92];
    assign wire_12738 = lut_tile_10_5_chanxy_out[93];
    assign wire_12739 = lut_tile_10_5_chanxy_out[94];
    assign wire_12740 = lut_tile_10_5_chanxy_out[95];
    assign wire_12741 = lut_tile_10_5_chanxy_out[96];
    assign wire_12742 = lut_tile_10_5_chanxy_out[97];
    assign wire_12743 = lut_tile_10_5_chanxy_out[98];
    assign wire_12744 = lut_tile_10_5_chanxy_out[99];
    assign wire_12745 = lut_tile_10_5_chanxy_out[100];
    assign wire_12746 = lut_tile_10_5_chanxy_out[101];
    assign wire_12747 = lut_tile_10_5_chanxy_out[102];
    assign wire_12748 = lut_tile_10_5_chanxy_out[103];
    assign wire_12749 = lut_tile_10_5_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_6_chanxy_in = {wire_10289, wire_10288, wire_13018, wire_9901, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9782, wire_4035, wire_10319, wire_10198, wire_13016, wire_9929, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9784, wire_4035, wire_10213, wire_10212, wire_13014, wire_9927, wire_9839, wire_9838, wire_9829, wire_9828, wire_9819, wire_9818, wire_9786, wire_4035, wire_10271, wire_10270, wire_13012, wire_9925, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9788, wire_3525, wire_10301, wire_10180, wire_13010, wire_9923, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9790, wire_3525, wire_10225, wire_10224, wire_13008, wire_9921, wire_9837, wire_9836, wire_9827, wire_9826, wire_9817, wire_9816, wire_9792, wire_3525, wire_10283, wire_10282, wire_13006, wire_9919, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9794, wire_4039, wire_3525, wire_10313, wire_10192, wire_13004, wire_9917, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9796, wire_4039, wire_3525, wire_10207, wire_10206, wire_13002, wire_9915, wire_9835, wire_9834, wire_9825, wire_9824, wire_9815, wire_9814, wire_9798, wire_4039, wire_3525, wire_10265, wire_10264, wire_4039, wire_13000, wire_9913, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9800, wire_4039, wire_3521, wire_10295, wire_10174, wire_4039, wire_12998, wire_9911, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9802, wire_4039, wire_3521, wire_10219, wire_10218, wire_4035, wire_12996, wire_9909, wire_9833, wire_9832, wire_9823, wire_9822, wire_9813, wire_9812, wire_9804, wire_4039, wire_3521, wire_10277, wire_10276, wire_3525, wire_12994, wire_9907, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9806, wire_4035, wire_3521, wire_10307, wire_10186, wire_3525, wire_12992, wire_9905, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9808, wire_4035, wire_3521, wire_10201, wire_10200, wire_3521, wire_12990, wire_9903, wire_9831, wire_9830, wire_9821, wire_9820, wire_9811, wire_9810, wire_9780, wire_4035, wire_3521, wire_10259, wire_10258, wire_10243, wire_10242, wire_10227, wire_10226, wire_10241, wire_10240, wire_10255, wire_10254, wire_10209, wire_10208, wire_10253, wire_10252, wire_10237, wire_10236, wire_10221, wire_10220, wire_10235, wire_10234, wire_4039, wire_10249, wire_10248, wire_4039, wire_10203, wire_10202, wire_4035, wire_10247, wire_10246, wire_3525, wire_10231, wire_10230, wire_3525, wire_10215, wire_10214, wire_3521, wire_10273, wire_10272, wire_10287, wire_10286, wire_10317, wire_10196, wire_10285, wire_10284, wire_10269, wire_10268, wire_10299, wire_10178, wire_10267, wire_10266, wire_10281, wire_10280, wire_10311, wire_10190, wire_10279, wire_10278, wire_4039, wire_10263, wire_10262, wire_4035, wire_10293, wire_10172, wire_4035, wire_10261, wire_10260, wire_3525, wire_10275, wire_10274, wire_3521, wire_10305, wire_10184, wire_3521, wire_10229, wire_10228, wire_10257, wire_10256, wire_10303, wire_10182, wire_10211, wire_10210, wire_10239, wire_10238, wire_10315, wire_10194, wire_10223, wire_10222, wire_10251, wire_10250, wire_10297, wire_10176, wire_10205, wire_10204, wire_4039, wire_10233, wire_10232, wire_4035, wire_10309, wire_10188, wire_4035, wire_10217, wire_10216, wire_3525, wire_10245, wire_10244, wire_3521, wire_10291, wire_10170, wire_3521, wire_12726, wire_12704, wire_12682, wire_12658, wire_10168, wire_3574, wire_3568, wire_3559, wire_3553, wire_12748, wire_12696, wire_12674, wire_12650, wire_10166, wire_3574, wire_3568, wire_3559, wire_3553, wire_12740, wire_12718, wire_12666, wire_12642, wire_10164, wire_3574, wire_3568, wire_3559, wire_3553, wire_12732, wire_12710, wire_12688, wire_12634, wire_10162, wire_3574, wire_3565, wire_3559, wire_3524, wire_12724, wire_12702, wire_12680, wire_12656, wire_10160, wire_3574, wire_3565, wire_3559, wire_3524, wire_12746, wire_12694, wire_12672, wire_12648, wire_10158, wire_3574, wire_3565, wire_3559, wire_3524, wire_12738, wire_12716, wire_12664, wire_12640, wire_10156, wire_3571, wire_3565, wire_3556, wire_3524, wire_12730, wire_12708, wire_12686, wire_12632, wire_10154, wire_3571, wire_3565, wire_3556, wire_3524, wire_12722, wire_12700, wire_12678, wire_12654, wire_10152, wire_3571, wire_3565, wire_3556, wire_3524, wire_12744, wire_12692, wire_12670, wire_12646, wire_10150, wire_3571, wire_3562, wire_3556, wire_3520, wire_12736, wire_12714, wire_12662, wire_12638, wire_10148, wire_3571, wire_3562, wire_3556, wire_3520, wire_12728, wire_12706, wire_12684, wire_12630, wire_10146, wire_3571, wire_3562, wire_3556, wire_3520, wire_12720, wire_12698, wire_12676, wire_12652, wire_10144, wire_3568, wire_3562, wire_3553, wire_3520, wire_12742, wire_12690, wire_12668, wire_12644, wire_10142, wire_3568, wire_3562, wire_3553, wire_3520, wire_12734, wire_12712, wire_12660, wire_12636, wire_10140, wire_3568, wire_3562, wire_3553, wire_3520, wire_13138, wire_13086, wire_13064, wire_13042, wire_10319, wire_3574, wire_3568, wire_3559, wire_3553, wire_13130, wire_13108, wire_13056, wire_13034, wire_10317, wire_3574, wire_3568, wire_3559, wire_3553, wire_13122, wire_13100, wire_13078, wire_13026, wire_10315, wire_3574, wire_3568, wire_3559, wire_3553, wire_13114, wire_13092, wire_13070, wire_13048, wire_10313, wire_3574, wire_3565, wire_3559, wire_3524, wire_13136, wire_13084, wire_13062, wire_13040, wire_10311, wire_3574, wire_3565, wire_3559, wire_3524, wire_13128, wire_13106, wire_13054, wire_13032, wire_10309, wire_3574, wire_3565, wire_3559, wire_3524, wire_13120, wire_13098, wire_13076, wire_13024, wire_10307, wire_3571, wire_3565, wire_3556, wire_3524, wire_13112, wire_13090, wire_13068, wire_13046, wire_10305, wire_3571, wire_3565, wire_3556, wire_3524, wire_13134, wire_13082, wire_13060, wire_13038, wire_10303, wire_3571, wire_3565, wire_3556, wire_3524, wire_13126, wire_13104, wire_13052, wire_13030, wire_10301, wire_3571, wire_3562, wire_3556, wire_3520, wire_13118, wire_13096, wire_13074, wire_13022, wire_10299, wire_3571, wire_3562, wire_3556, wire_3520, wire_13110, wire_13088, wire_13066, wire_13044, wire_10297, wire_3571, wire_3562, wire_3556, wire_3520, wire_13132, wire_13080, wire_13058, wire_13036, wire_10295, wire_3568, wire_3562, wire_3553, wire_3520, wire_13124, wire_13102, wire_13050, wire_13028, wire_10293, wire_3568, wire_3562, wire_3553, wire_3520, wire_13116, wire_13094, wire_13072, wire_13020, wire_10291, wire_3568, wire_3562, wire_3553, wire_3520};
    // CHNAXY TOTAL: 573
    assign wire_10171 = lut_tile_10_6_chanxy_out[0];
    assign wire_10173 = lut_tile_10_6_chanxy_out[1];
    assign wire_10175 = lut_tile_10_6_chanxy_out[2];
    assign wire_10177 = lut_tile_10_6_chanxy_out[3];
    assign wire_10179 = lut_tile_10_6_chanxy_out[4];
    assign wire_10181 = lut_tile_10_6_chanxy_out[5];
    assign wire_10183 = lut_tile_10_6_chanxy_out[6];
    assign wire_10185 = lut_tile_10_6_chanxy_out[7];
    assign wire_10187 = lut_tile_10_6_chanxy_out[8];
    assign wire_10189 = lut_tile_10_6_chanxy_out[9];
    assign wire_10191 = lut_tile_10_6_chanxy_out[10];
    assign wire_10193 = lut_tile_10_6_chanxy_out[11];
    assign wire_10195 = lut_tile_10_6_chanxy_out[12];
    assign wire_10197 = lut_tile_10_6_chanxy_out[13];
    assign wire_10199 = lut_tile_10_6_chanxy_out[14];
    assign wire_10260 = lut_tile_10_6_chanxy_out[15];
    assign wire_10262 = lut_tile_10_6_chanxy_out[16];
    assign wire_10264 = lut_tile_10_6_chanxy_out[17];
    assign wire_10266 = lut_tile_10_6_chanxy_out[18];
    assign wire_10268 = lut_tile_10_6_chanxy_out[19];
    assign wire_10270 = lut_tile_10_6_chanxy_out[20];
    assign wire_10272 = lut_tile_10_6_chanxy_out[21];
    assign wire_10274 = lut_tile_10_6_chanxy_out[22];
    assign wire_10276 = lut_tile_10_6_chanxy_out[23];
    assign wire_10278 = lut_tile_10_6_chanxy_out[24];
    assign wire_10280 = lut_tile_10_6_chanxy_out[25];
    assign wire_10282 = lut_tile_10_6_chanxy_out[26];
    assign wire_10284 = lut_tile_10_6_chanxy_out[27];
    assign wire_10286 = lut_tile_10_6_chanxy_out[28];
    assign wire_10288 = lut_tile_10_6_chanxy_out[29];
    assign wire_13021 = lut_tile_10_6_chanxy_out[30];
    assign wire_13023 = lut_tile_10_6_chanxy_out[31];
    assign wire_13025 = lut_tile_10_6_chanxy_out[32];
    assign wire_13027 = lut_tile_10_6_chanxy_out[33];
    assign wire_13029 = lut_tile_10_6_chanxy_out[34];
    assign wire_13031 = lut_tile_10_6_chanxy_out[35];
    assign wire_13033 = lut_tile_10_6_chanxy_out[36];
    assign wire_13035 = lut_tile_10_6_chanxy_out[37];
    assign wire_13037 = lut_tile_10_6_chanxy_out[38];
    assign wire_13039 = lut_tile_10_6_chanxy_out[39];
    assign wire_13041 = lut_tile_10_6_chanxy_out[40];
    assign wire_13043 = lut_tile_10_6_chanxy_out[41];
    assign wire_13045 = lut_tile_10_6_chanxy_out[42];
    assign wire_13047 = lut_tile_10_6_chanxy_out[43];
    assign wire_13049 = lut_tile_10_6_chanxy_out[44];
    assign wire_13051 = lut_tile_10_6_chanxy_out[45];
    assign wire_13053 = lut_tile_10_6_chanxy_out[46];
    assign wire_13055 = lut_tile_10_6_chanxy_out[47];
    assign wire_13057 = lut_tile_10_6_chanxy_out[48];
    assign wire_13059 = lut_tile_10_6_chanxy_out[49];
    assign wire_13061 = lut_tile_10_6_chanxy_out[50];
    assign wire_13063 = lut_tile_10_6_chanxy_out[51];
    assign wire_13065 = lut_tile_10_6_chanxy_out[52];
    assign wire_13067 = lut_tile_10_6_chanxy_out[53];
    assign wire_13069 = lut_tile_10_6_chanxy_out[54];
    assign wire_13071 = lut_tile_10_6_chanxy_out[55];
    assign wire_13073 = lut_tile_10_6_chanxy_out[56];
    assign wire_13075 = lut_tile_10_6_chanxy_out[57];
    assign wire_13077 = lut_tile_10_6_chanxy_out[58];
    assign wire_13079 = lut_tile_10_6_chanxy_out[59];
    assign wire_13081 = lut_tile_10_6_chanxy_out[60];
    assign wire_13083 = lut_tile_10_6_chanxy_out[61];
    assign wire_13085 = lut_tile_10_6_chanxy_out[62];
    assign wire_13087 = lut_tile_10_6_chanxy_out[63];
    assign wire_13089 = lut_tile_10_6_chanxy_out[64];
    assign wire_13091 = lut_tile_10_6_chanxy_out[65];
    assign wire_13093 = lut_tile_10_6_chanxy_out[66];
    assign wire_13095 = lut_tile_10_6_chanxy_out[67];
    assign wire_13097 = lut_tile_10_6_chanxy_out[68];
    assign wire_13099 = lut_tile_10_6_chanxy_out[69];
    assign wire_13101 = lut_tile_10_6_chanxy_out[70];
    assign wire_13103 = lut_tile_10_6_chanxy_out[71];
    assign wire_13105 = lut_tile_10_6_chanxy_out[72];
    assign wire_13107 = lut_tile_10_6_chanxy_out[73];
    assign wire_13109 = lut_tile_10_6_chanxy_out[74];
    assign wire_13110 = lut_tile_10_6_chanxy_out[75];
    assign wire_13111 = lut_tile_10_6_chanxy_out[76];
    assign wire_13112 = lut_tile_10_6_chanxy_out[77];
    assign wire_13113 = lut_tile_10_6_chanxy_out[78];
    assign wire_13114 = lut_tile_10_6_chanxy_out[79];
    assign wire_13115 = lut_tile_10_6_chanxy_out[80];
    assign wire_13116 = lut_tile_10_6_chanxy_out[81];
    assign wire_13117 = lut_tile_10_6_chanxy_out[82];
    assign wire_13118 = lut_tile_10_6_chanxy_out[83];
    assign wire_13119 = lut_tile_10_6_chanxy_out[84];
    assign wire_13120 = lut_tile_10_6_chanxy_out[85];
    assign wire_13121 = lut_tile_10_6_chanxy_out[86];
    assign wire_13122 = lut_tile_10_6_chanxy_out[87];
    assign wire_13123 = lut_tile_10_6_chanxy_out[88];
    assign wire_13124 = lut_tile_10_6_chanxy_out[89];
    assign wire_13125 = lut_tile_10_6_chanxy_out[90];
    assign wire_13126 = lut_tile_10_6_chanxy_out[91];
    assign wire_13127 = lut_tile_10_6_chanxy_out[92];
    assign wire_13128 = lut_tile_10_6_chanxy_out[93];
    assign wire_13129 = lut_tile_10_6_chanxy_out[94];
    assign wire_13130 = lut_tile_10_6_chanxy_out[95];
    assign wire_13131 = lut_tile_10_6_chanxy_out[96];
    assign wire_13132 = lut_tile_10_6_chanxy_out[97];
    assign wire_13133 = lut_tile_10_6_chanxy_out[98];
    assign wire_13134 = lut_tile_10_6_chanxy_out[99];
    assign wire_13135 = lut_tile_10_6_chanxy_out[100];
    assign wire_13136 = lut_tile_10_6_chanxy_out[101];
    assign wire_13137 = lut_tile_10_6_chanxy_out[102];
    assign wire_13138 = lut_tile_10_6_chanxy_out[103];
    assign wire_13139 = lut_tile_10_6_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_7_chanxy_in = {wire_10349, wire_10228, wire_13408, wire_9931, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9812, wire_4551, wire_10257, wire_10256, wire_13406, wire_9959, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9814, wire_4551, wire_10303, wire_10302, wire_13404, wire_9957, wire_9869, wire_9868, wire_9859, wire_9858, wire_9849, wire_9848, wire_9816, wire_4551, wire_10331, wire_10210, wire_13402, wire_9955, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9818, wire_4041, wire_10239, wire_10238, wire_13400, wire_9953, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9820, wire_4041, wire_10315, wire_10314, wire_13398, wire_9951, wire_9867, wire_9866, wire_9857, wire_9856, wire_9847, wire_9846, wire_9822, wire_4041, wire_10343, wire_10222, wire_13396, wire_9949, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9824, wire_4555, wire_4041, wire_10251, wire_10250, wire_13394, wire_9947, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9826, wire_4555, wire_4041, wire_10297, wire_10296, wire_13392, wire_9945, wire_9865, wire_9864, wire_9855, wire_9854, wire_9845, wire_9844, wire_9828, wire_4555, wire_4041, wire_10325, wire_10204, wire_4555, wire_13390, wire_9943, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9830, wire_4555, wire_4037, wire_10233, wire_10232, wire_4551, wire_13388, wire_9941, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9832, wire_4555, wire_4037, wire_10309, wire_10308, wire_4551, wire_13386, wire_9939, wire_9863, wire_9862, wire_9853, wire_9852, wire_9843, wire_9842, wire_9834, wire_4555, wire_4037, wire_10337, wire_10216, wire_4041, wire_13384, wire_9937, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9836, wire_4551, wire_4037, wire_10245, wire_10244, wire_4037, wire_13382, wire_9935, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9838, wire_4551, wire_4037, wire_10291, wire_10290, wire_4037, wire_13380, wire_9933, wire_9861, wire_9860, wire_9851, wire_9850, wire_9841, wire_9840, wire_9810, wire_4551, wire_4037, wire_10289, wire_10288, wire_10319, wire_10318, wire_10333, wire_10212, wire_10271, wire_10270, wire_10301, wire_10300, wire_10345, wire_10224, wire_10283, wire_10282, wire_10313, wire_10312, wire_10327, wire_10206, wire_10265, wire_10264, wire_4555, wire_10295, wire_10294, wire_4555, wire_10339, wire_10218, wire_4551, wire_10277, wire_10276, wire_4041, wire_10307, wire_10306, wire_4041, wire_10321, wire_10200, wire_4037, wire_10259, wire_10258, wire_10243, wire_10242, wire_10347, wire_10226, wire_10241, wire_10240, wire_10255, wire_10254, wire_10329, wire_10208, wire_10253, wire_10252, wire_10237, wire_10236, wire_10341, wire_10220, wire_10235, wire_10234, wire_4555, wire_10249, wire_10248, wire_4555, wire_10323, wire_10202, wire_4551, wire_10247, wire_10246, wire_4041, wire_10231, wire_10230, wire_4041, wire_10335, wire_10214, wire_4037, wire_10273, wire_10272, wire_10287, wire_10286, wire_10317, wire_10316, wire_10285, wire_10284, wire_10269, wire_10268, wire_10299, wire_10298, wire_10267, wire_10266, wire_10281, wire_10280, wire_10311, wire_10310, wire_10279, wire_10278, wire_4555, wire_10263, wire_10262, wire_4551, wire_10293, wire_10292, wire_4551, wire_10261, wire_10260, wire_4041, wire_10275, wire_10274, wire_4037, wire_10305, wire_10304, wire_4037, wire_13138, wire_13086, wire_13064, wire_13042, wire_10198, wire_4090, wire_4084, wire_4075, wire_4069, wire_13130, wire_13108, wire_13056, wire_13034, wire_10196, wire_4090, wire_4084, wire_4075, wire_4069, wire_13122, wire_13100, wire_13078, wire_13026, wire_10194, wire_4090, wire_4084, wire_4075, wire_4069, wire_13114, wire_13092, wire_13070, wire_13048, wire_10192, wire_4090, wire_4081, wire_4075, wire_4040, wire_13136, wire_13084, wire_13062, wire_13040, wire_10190, wire_4090, wire_4081, wire_4075, wire_4040, wire_13128, wire_13106, wire_13054, wire_13032, wire_10188, wire_4090, wire_4081, wire_4075, wire_4040, wire_13120, wire_13098, wire_13076, wire_13024, wire_10186, wire_4087, wire_4081, wire_4072, wire_4040, wire_13112, wire_13090, wire_13068, wire_13046, wire_10184, wire_4087, wire_4081, wire_4072, wire_4040, wire_13134, wire_13082, wire_13060, wire_13038, wire_10182, wire_4087, wire_4081, wire_4072, wire_4040, wire_13126, wire_13104, wire_13052, wire_13030, wire_10180, wire_4087, wire_4078, wire_4072, wire_4036, wire_13118, wire_13096, wire_13074, wire_13022, wire_10178, wire_4087, wire_4078, wire_4072, wire_4036, wire_13110, wire_13088, wire_13066, wire_13044, wire_10176, wire_4087, wire_4078, wire_4072, wire_4036, wire_13132, wire_13080, wire_13058, wire_13036, wire_10174, wire_4084, wire_4078, wire_4069, wire_4036, wire_13124, wire_13102, wire_13050, wire_13028, wire_10172, wire_4084, wire_4078, wire_4069, wire_4036, wire_13116, wire_13094, wire_13072, wire_13020, wire_10170, wire_4084, wire_4078, wire_4069, wire_4036, wire_13522, wire_13498, wire_13446, wire_13424, wire_10349, wire_4090, wire_4084, wire_4075, wire_4069, wire_13514, wire_13490, wire_13468, wire_13416, wire_10347, wire_4090, wire_4084, wire_4075, wire_4069, wire_13506, wire_13482, wire_13460, wire_13438, wire_10345, wire_4090, wire_4084, wire_4075, wire_4069, wire_13528, wire_13474, wire_13452, wire_13430, wire_10343, wire_4090, wire_4081, wire_4075, wire_4040, wire_13520, wire_13496, wire_13444, wire_13422, wire_10341, wire_4090, wire_4081, wire_4075, wire_4040, wire_13512, wire_13488, wire_13466, wire_13414, wire_10339, wire_4090, wire_4081, wire_4075, wire_4040, wire_13504, wire_13480, wire_13458, wire_13436, wire_10337, wire_4087, wire_4081, wire_4072, wire_4040, wire_13526, wire_13472, wire_13450, wire_13428, wire_10335, wire_4087, wire_4081, wire_4072, wire_4040, wire_13518, wire_13494, wire_13442, wire_13420, wire_10333, wire_4087, wire_4081, wire_4072, wire_4040, wire_13510, wire_13486, wire_13464, wire_13412, wire_10331, wire_4087, wire_4078, wire_4072, wire_4036, wire_13502, wire_13478, wire_13456, wire_13434, wire_10329, wire_4087, wire_4078, wire_4072, wire_4036, wire_13524, wire_13470, wire_13448, wire_13426, wire_10327, wire_4087, wire_4078, wire_4072, wire_4036, wire_13516, wire_13492, wire_13440, wire_13418, wire_10325, wire_4084, wire_4078, wire_4069, wire_4036, wire_13508, wire_13484, wire_13462, wire_13410, wire_10323, wire_4084, wire_4078, wire_4069, wire_4036, wire_13500, wire_13476, wire_13454, wire_13432, wire_10321, wire_4084, wire_4078, wire_4069, wire_4036};
    // CHNAXY TOTAL: 573
    assign wire_10201 = lut_tile_10_7_chanxy_out[0];
    assign wire_10203 = lut_tile_10_7_chanxy_out[1];
    assign wire_10205 = lut_tile_10_7_chanxy_out[2];
    assign wire_10207 = lut_tile_10_7_chanxy_out[3];
    assign wire_10209 = lut_tile_10_7_chanxy_out[4];
    assign wire_10211 = lut_tile_10_7_chanxy_out[5];
    assign wire_10213 = lut_tile_10_7_chanxy_out[6];
    assign wire_10215 = lut_tile_10_7_chanxy_out[7];
    assign wire_10217 = lut_tile_10_7_chanxy_out[8];
    assign wire_10219 = lut_tile_10_7_chanxy_out[9];
    assign wire_10221 = lut_tile_10_7_chanxy_out[10];
    assign wire_10223 = lut_tile_10_7_chanxy_out[11];
    assign wire_10225 = lut_tile_10_7_chanxy_out[12];
    assign wire_10227 = lut_tile_10_7_chanxy_out[13];
    assign wire_10229 = lut_tile_10_7_chanxy_out[14];
    assign wire_10290 = lut_tile_10_7_chanxy_out[15];
    assign wire_10292 = lut_tile_10_7_chanxy_out[16];
    assign wire_10294 = lut_tile_10_7_chanxy_out[17];
    assign wire_10296 = lut_tile_10_7_chanxy_out[18];
    assign wire_10298 = lut_tile_10_7_chanxy_out[19];
    assign wire_10300 = lut_tile_10_7_chanxy_out[20];
    assign wire_10302 = lut_tile_10_7_chanxy_out[21];
    assign wire_10304 = lut_tile_10_7_chanxy_out[22];
    assign wire_10306 = lut_tile_10_7_chanxy_out[23];
    assign wire_10308 = lut_tile_10_7_chanxy_out[24];
    assign wire_10310 = lut_tile_10_7_chanxy_out[25];
    assign wire_10312 = lut_tile_10_7_chanxy_out[26];
    assign wire_10314 = lut_tile_10_7_chanxy_out[27];
    assign wire_10316 = lut_tile_10_7_chanxy_out[28];
    assign wire_10318 = lut_tile_10_7_chanxy_out[29];
    assign wire_13411 = lut_tile_10_7_chanxy_out[30];
    assign wire_13413 = lut_tile_10_7_chanxy_out[31];
    assign wire_13415 = lut_tile_10_7_chanxy_out[32];
    assign wire_13417 = lut_tile_10_7_chanxy_out[33];
    assign wire_13419 = lut_tile_10_7_chanxy_out[34];
    assign wire_13421 = lut_tile_10_7_chanxy_out[35];
    assign wire_13423 = lut_tile_10_7_chanxy_out[36];
    assign wire_13425 = lut_tile_10_7_chanxy_out[37];
    assign wire_13427 = lut_tile_10_7_chanxy_out[38];
    assign wire_13429 = lut_tile_10_7_chanxy_out[39];
    assign wire_13431 = lut_tile_10_7_chanxy_out[40];
    assign wire_13433 = lut_tile_10_7_chanxy_out[41];
    assign wire_13435 = lut_tile_10_7_chanxy_out[42];
    assign wire_13437 = lut_tile_10_7_chanxy_out[43];
    assign wire_13439 = lut_tile_10_7_chanxy_out[44];
    assign wire_13441 = lut_tile_10_7_chanxy_out[45];
    assign wire_13443 = lut_tile_10_7_chanxy_out[46];
    assign wire_13445 = lut_tile_10_7_chanxy_out[47];
    assign wire_13447 = lut_tile_10_7_chanxy_out[48];
    assign wire_13449 = lut_tile_10_7_chanxy_out[49];
    assign wire_13451 = lut_tile_10_7_chanxy_out[50];
    assign wire_13453 = lut_tile_10_7_chanxy_out[51];
    assign wire_13455 = lut_tile_10_7_chanxy_out[52];
    assign wire_13457 = lut_tile_10_7_chanxy_out[53];
    assign wire_13459 = lut_tile_10_7_chanxy_out[54];
    assign wire_13461 = lut_tile_10_7_chanxy_out[55];
    assign wire_13463 = lut_tile_10_7_chanxy_out[56];
    assign wire_13465 = lut_tile_10_7_chanxy_out[57];
    assign wire_13467 = lut_tile_10_7_chanxy_out[58];
    assign wire_13469 = lut_tile_10_7_chanxy_out[59];
    assign wire_13471 = lut_tile_10_7_chanxy_out[60];
    assign wire_13473 = lut_tile_10_7_chanxy_out[61];
    assign wire_13475 = lut_tile_10_7_chanxy_out[62];
    assign wire_13477 = lut_tile_10_7_chanxy_out[63];
    assign wire_13479 = lut_tile_10_7_chanxy_out[64];
    assign wire_13481 = lut_tile_10_7_chanxy_out[65];
    assign wire_13483 = lut_tile_10_7_chanxy_out[66];
    assign wire_13485 = lut_tile_10_7_chanxy_out[67];
    assign wire_13487 = lut_tile_10_7_chanxy_out[68];
    assign wire_13489 = lut_tile_10_7_chanxy_out[69];
    assign wire_13491 = lut_tile_10_7_chanxy_out[70];
    assign wire_13493 = lut_tile_10_7_chanxy_out[71];
    assign wire_13495 = lut_tile_10_7_chanxy_out[72];
    assign wire_13497 = lut_tile_10_7_chanxy_out[73];
    assign wire_13499 = lut_tile_10_7_chanxy_out[74];
    assign wire_13500 = lut_tile_10_7_chanxy_out[75];
    assign wire_13501 = lut_tile_10_7_chanxy_out[76];
    assign wire_13502 = lut_tile_10_7_chanxy_out[77];
    assign wire_13503 = lut_tile_10_7_chanxy_out[78];
    assign wire_13504 = lut_tile_10_7_chanxy_out[79];
    assign wire_13505 = lut_tile_10_7_chanxy_out[80];
    assign wire_13506 = lut_tile_10_7_chanxy_out[81];
    assign wire_13507 = lut_tile_10_7_chanxy_out[82];
    assign wire_13508 = lut_tile_10_7_chanxy_out[83];
    assign wire_13509 = lut_tile_10_7_chanxy_out[84];
    assign wire_13510 = lut_tile_10_7_chanxy_out[85];
    assign wire_13511 = lut_tile_10_7_chanxy_out[86];
    assign wire_13512 = lut_tile_10_7_chanxy_out[87];
    assign wire_13513 = lut_tile_10_7_chanxy_out[88];
    assign wire_13514 = lut_tile_10_7_chanxy_out[89];
    assign wire_13515 = lut_tile_10_7_chanxy_out[90];
    assign wire_13516 = lut_tile_10_7_chanxy_out[91];
    assign wire_13517 = lut_tile_10_7_chanxy_out[92];
    assign wire_13518 = lut_tile_10_7_chanxy_out[93];
    assign wire_13519 = lut_tile_10_7_chanxy_out[94];
    assign wire_13520 = lut_tile_10_7_chanxy_out[95];
    assign wire_13521 = lut_tile_10_7_chanxy_out[96];
    assign wire_13522 = lut_tile_10_7_chanxy_out[97];
    assign wire_13523 = lut_tile_10_7_chanxy_out[98];
    assign wire_13524 = lut_tile_10_7_chanxy_out[99];
    assign wire_13525 = lut_tile_10_7_chanxy_out[100];
    assign wire_13526 = lut_tile_10_7_chanxy_out[101];
    assign wire_13527 = lut_tile_10_7_chanxy_out[102];
    assign wire_13528 = lut_tile_10_7_chanxy_out[103];
    assign wire_13529 = lut_tile_10_7_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_8_chanxy_in = {wire_10273, wire_10272, wire_13798, wire_9961, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9842, wire_5067, wire_10287, wire_10286, wire_13796, wire_9989, wire_9899, wire_9898, wire_9889, wire_9888, wire_9879, wire_9878, wire_9844, wire_5067, wire_10317, wire_10316, wire_13794, wire_9987, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9846, wire_5067, wire_10285, wire_10284, wire_13792, wire_9985, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9848, wire_4557, wire_10269, wire_10268, wire_13790, wire_9983, wire_9897, wire_9896, wire_9887, wire_9886, wire_9877, wire_9876, wire_9850, wire_4557, wire_10299, wire_10298, wire_13788, wire_9981, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9852, wire_4557, wire_10267, wire_10266, wire_13786, wire_9979, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9854, wire_5071, wire_4557, wire_10281, wire_10280, wire_13784, wire_9977, wire_9895, wire_9894, wire_9885, wire_9884, wire_9875, wire_9874, wire_9856, wire_5071, wire_4557, wire_10311, wire_10310, wire_13782, wire_9975, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9858, wire_5071, wire_4557, wire_10279, wire_10278, wire_5071, wire_13780, wire_9973, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9860, wire_5071, wire_4553, wire_10263, wire_10262, wire_5067, wire_13778, wire_9971, wire_9893, wire_9892, wire_9883, wire_9882, wire_9873, wire_9872, wire_9862, wire_5071, wire_4553, wire_10293, wire_10292, wire_5067, wire_13776, wire_9969, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9864, wire_5071, wire_4553, wire_10261, wire_10260, wire_4557, wire_13774, wire_9967, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9866, wire_5067, wire_4553, wire_10275, wire_10274, wire_4553, wire_13772, wire_9965, wire_9891, wire_9890, wire_9881, wire_9880, wire_9871, wire_9870, wire_9868, wire_5067, wire_4553, wire_10305, wire_10304, wire_4553, wire_13770, wire_9963, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9840, wire_5067, wire_4553, wire_10349, wire_10348, wire_10377, wire_10256, wire_10303, wire_10302, wire_10331, wire_10330, wire_10359, wire_10238, wire_10315, wire_10314, wire_10343, wire_10342, wire_10371, wire_10250, wire_10297, wire_10296, wire_10325, wire_10324, wire_5071, wire_10353, wire_10232, wire_5067, wire_10309, wire_10308, wire_5067, wire_10337, wire_10336, wire_4557, wire_10365, wire_10244, wire_4553, wire_10291, wire_10290, wire_4553, wire_10289, wire_10288, wire_10319, wire_10318, wire_10333, wire_10332, wire_10271, wire_10270, wire_10301, wire_10300, wire_10345, wire_10344, wire_10283, wire_10282, wire_10313, wire_10312, wire_10327, wire_10326, wire_10265, wire_10264, wire_5071, wire_10295, wire_10294, wire_5071, wire_10339, wire_10338, wire_5067, wire_10277, wire_10276, wire_4557, wire_10307, wire_10306, wire_4557, wire_10321, wire_10320, wire_4553, wire_10379, wire_10258, wire_10363, wire_10242, wire_10347, wire_10346, wire_10361, wire_10240, wire_10375, wire_10254, wire_10329, wire_10328, wire_10373, wire_10252, wire_10357, wire_10236, wire_10341, wire_10340, wire_10355, wire_10234, wire_5071, wire_10369, wire_10248, wire_5071, wire_10323, wire_10322, wire_5067, wire_10367, wire_10246, wire_4557, wire_10351, wire_10230, wire_4557, wire_10335, wire_10334, wire_4553, wire_13522, wire_13498, wire_13446, wire_13424, wire_10228, wire_4606, wire_4600, wire_4591, wire_4585, wire_13514, wire_13490, wire_13468, wire_13416, wire_10226, wire_4606, wire_4600, wire_4591, wire_4585, wire_13506, wire_13482, wire_13460, wire_13438, wire_10224, wire_4606, wire_4600, wire_4591, wire_4585, wire_13528, wire_13474, wire_13452, wire_13430, wire_10222, wire_4606, wire_4597, wire_4591, wire_4556, wire_13520, wire_13496, wire_13444, wire_13422, wire_10220, wire_4606, wire_4597, wire_4591, wire_4556, wire_13512, wire_13488, wire_13466, wire_13414, wire_10218, wire_4606, wire_4597, wire_4591, wire_4556, wire_13504, wire_13480, wire_13458, wire_13436, wire_10216, wire_4603, wire_4597, wire_4588, wire_4556, wire_13526, wire_13472, wire_13450, wire_13428, wire_10214, wire_4603, wire_4597, wire_4588, wire_4556, wire_13518, wire_13494, wire_13442, wire_13420, wire_10212, wire_4603, wire_4597, wire_4588, wire_4556, wire_13510, wire_13486, wire_13464, wire_13412, wire_10210, wire_4603, wire_4594, wire_4588, wire_4552, wire_13502, wire_13478, wire_13456, wire_13434, wire_10208, wire_4603, wire_4594, wire_4588, wire_4552, wire_13524, wire_13470, wire_13448, wire_13426, wire_10206, wire_4603, wire_4594, wire_4588, wire_4552, wire_13516, wire_13492, wire_13440, wire_13418, wire_10204, wire_4600, wire_4594, wire_4585, wire_4552, wire_13508, wire_13484, wire_13462, wire_13410, wire_10202, wire_4600, wire_4594, wire_4585, wire_4552, wire_13500, wire_13476, wire_13454, wire_13432, wire_10200, wire_4600, wire_4594, wire_4585, wire_4552, wire_13904, wire_13882, wire_13858, wire_13806, wire_10379, wire_4606, wire_4600, wire_4591, wire_4585, wire_13896, wire_13874, wire_13850, wire_13828, wire_10377, wire_4606, wire_4600, wire_4591, wire_4585, wire_13918, wire_13866, wire_13842, wire_13820, wire_10375, wire_4606, wire_4600, wire_4591, wire_4585, wire_13910, wire_13888, wire_13834, wire_13812, wire_10373, wire_4606, wire_4597, wire_4591, wire_4556, wire_13902, wire_13880, wire_13856, wire_13804, wire_10371, wire_4606, wire_4597, wire_4591, wire_4556, wire_13894, wire_13872, wire_13848, wire_13826, wire_10369, wire_4606, wire_4597, wire_4591, wire_4556, wire_13916, wire_13864, wire_13840, wire_13818, wire_10367, wire_4603, wire_4597, wire_4588, wire_4556, wire_13908, wire_13886, wire_13832, wire_13810, wire_10365, wire_4603, wire_4597, wire_4588, wire_4556, wire_13900, wire_13878, wire_13854, wire_13802, wire_10363, wire_4603, wire_4597, wire_4588, wire_4556, wire_13892, wire_13870, wire_13846, wire_13824, wire_10361, wire_4603, wire_4594, wire_4588, wire_4552, wire_13914, wire_13862, wire_13838, wire_13816, wire_10359, wire_4603, wire_4594, wire_4588, wire_4552, wire_13906, wire_13884, wire_13830, wire_13808, wire_10357, wire_4603, wire_4594, wire_4588, wire_4552, wire_13898, wire_13876, wire_13852, wire_13800, wire_10355, wire_4600, wire_4594, wire_4585, wire_4552, wire_13890, wire_13868, wire_13844, wire_13822, wire_10353, wire_4600, wire_4594, wire_4585, wire_4552, wire_13912, wire_13860, wire_13836, wire_13814, wire_10351, wire_4600, wire_4594, wire_4585, wire_4552};
    // CHNAXY TOTAL: 573
    assign wire_10231 = lut_tile_10_8_chanxy_out[0];
    assign wire_10233 = lut_tile_10_8_chanxy_out[1];
    assign wire_10235 = lut_tile_10_8_chanxy_out[2];
    assign wire_10237 = lut_tile_10_8_chanxy_out[3];
    assign wire_10239 = lut_tile_10_8_chanxy_out[4];
    assign wire_10241 = lut_tile_10_8_chanxy_out[5];
    assign wire_10243 = lut_tile_10_8_chanxy_out[6];
    assign wire_10245 = lut_tile_10_8_chanxy_out[7];
    assign wire_10247 = lut_tile_10_8_chanxy_out[8];
    assign wire_10249 = lut_tile_10_8_chanxy_out[9];
    assign wire_10251 = lut_tile_10_8_chanxy_out[10];
    assign wire_10253 = lut_tile_10_8_chanxy_out[11];
    assign wire_10255 = lut_tile_10_8_chanxy_out[12];
    assign wire_10257 = lut_tile_10_8_chanxy_out[13];
    assign wire_10259 = lut_tile_10_8_chanxy_out[14];
    assign wire_10320 = lut_tile_10_8_chanxy_out[15];
    assign wire_10322 = lut_tile_10_8_chanxy_out[16];
    assign wire_10324 = lut_tile_10_8_chanxy_out[17];
    assign wire_10326 = lut_tile_10_8_chanxy_out[18];
    assign wire_10328 = lut_tile_10_8_chanxy_out[19];
    assign wire_10330 = lut_tile_10_8_chanxy_out[20];
    assign wire_10332 = lut_tile_10_8_chanxy_out[21];
    assign wire_10334 = lut_tile_10_8_chanxy_out[22];
    assign wire_10336 = lut_tile_10_8_chanxy_out[23];
    assign wire_10338 = lut_tile_10_8_chanxy_out[24];
    assign wire_10340 = lut_tile_10_8_chanxy_out[25];
    assign wire_10342 = lut_tile_10_8_chanxy_out[26];
    assign wire_10344 = lut_tile_10_8_chanxy_out[27];
    assign wire_10346 = lut_tile_10_8_chanxy_out[28];
    assign wire_10348 = lut_tile_10_8_chanxy_out[29];
    assign wire_13801 = lut_tile_10_8_chanxy_out[30];
    assign wire_13803 = lut_tile_10_8_chanxy_out[31];
    assign wire_13805 = lut_tile_10_8_chanxy_out[32];
    assign wire_13807 = lut_tile_10_8_chanxy_out[33];
    assign wire_13809 = lut_tile_10_8_chanxy_out[34];
    assign wire_13811 = lut_tile_10_8_chanxy_out[35];
    assign wire_13813 = lut_tile_10_8_chanxy_out[36];
    assign wire_13815 = lut_tile_10_8_chanxy_out[37];
    assign wire_13817 = lut_tile_10_8_chanxy_out[38];
    assign wire_13819 = lut_tile_10_8_chanxy_out[39];
    assign wire_13821 = lut_tile_10_8_chanxy_out[40];
    assign wire_13823 = lut_tile_10_8_chanxy_out[41];
    assign wire_13825 = lut_tile_10_8_chanxy_out[42];
    assign wire_13827 = lut_tile_10_8_chanxy_out[43];
    assign wire_13829 = lut_tile_10_8_chanxy_out[44];
    assign wire_13831 = lut_tile_10_8_chanxy_out[45];
    assign wire_13833 = lut_tile_10_8_chanxy_out[46];
    assign wire_13835 = lut_tile_10_8_chanxy_out[47];
    assign wire_13837 = lut_tile_10_8_chanxy_out[48];
    assign wire_13839 = lut_tile_10_8_chanxy_out[49];
    assign wire_13841 = lut_tile_10_8_chanxy_out[50];
    assign wire_13843 = lut_tile_10_8_chanxy_out[51];
    assign wire_13845 = lut_tile_10_8_chanxy_out[52];
    assign wire_13847 = lut_tile_10_8_chanxy_out[53];
    assign wire_13849 = lut_tile_10_8_chanxy_out[54];
    assign wire_13851 = lut_tile_10_8_chanxy_out[55];
    assign wire_13853 = lut_tile_10_8_chanxy_out[56];
    assign wire_13855 = lut_tile_10_8_chanxy_out[57];
    assign wire_13857 = lut_tile_10_8_chanxy_out[58];
    assign wire_13859 = lut_tile_10_8_chanxy_out[59];
    assign wire_13861 = lut_tile_10_8_chanxy_out[60];
    assign wire_13863 = lut_tile_10_8_chanxy_out[61];
    assign wire_13865 = lut_tile_10_8_chanxy_out[62];
    assign wire_13867 = lut_tile_10_8_chanxy_out[63];
    assign wire_13869 = lut_tile_10_8_chanxy_out[64];
    assign wire_13871 = lut_tile_10_8_chanxy_out[65];
    assign wire_13873 = lut_tile_10_8_chanxy_out[66];
    assign wire_13875 = lut_tile_10_8_chanxy_out[67];
    assign wire_13877 = lut_tile_10_8_chanxy_out[68];
    assign wire_13879 = lut_tile_10_8_chanxy_out[69];
    assign wire_13881 = lut_tile_10_8_chanxy_out[70];
    assign wire_13883 = lut_tile_10_8_chanxy_out[71];
    assign wire_13885 = lut_tile_10_8_chanxy_out[72];
    assign wire_13887 = lut_tile_10_8_chanxy_out[73];
    assign wire_13889 = lut_tile_10_8_chanxy_out[74];
    assign wire_13890 = lut_tile_10_8_chanxy_out[75];
    assign wire_13891 = lut_tile_10_8_chanxy_out[76];
    assign wire_13892 = lut_tile_10_8_chanxy_out[77];
    assign wire_13893 = lut_tile_10_8_chanxy_out[78];
    assign wire_13894 = lut_tile_10_8_chanxy_out[79];
    assign wire_13895 = lut_tile_10_8_chanxy_out[80];
    assign wire_13896 = lut_tile_10_8_chanxy_out[81];
    assign wire_13897 = lut_tile_10_8_chanxy_out[82];
    assign wire_13898 = lut_tile_10_8_chanxy_out[83];
    assign wire_13899 = lut_tile_10_8_chanxy_out[84];
    assign wire_13900 = lut_tile_10_8_chanxy_out[85];
    assign wire_13901 = lut_tile_10_8_chanxy_out[86];
    assign wire_13902 = lut_tile_10_8_chanxy_out[87];
    assign wire_13903 = lut_tile_10_8_chanxy_out[88];
    assign wire_13904 = lut_tile_10_8_chanxy_out[89];
    assign wire_13905 = lut_tile_10_8_chanxy_out[90];
    assign wire_13906 = lut_tile_10_8_chanxy_out[91];
    assign wire_13907 = lut_tile_10_8_chanxy_out[92];
    assign wire_13908 = lut_tile_10_8_chanxy_out[93];
    assign wire_13909 = lut_tile_10_8_chanxy_out[94];
    assign wire_13910 = lut_tile_10_8_chanxy_out[95];
    assign wire_13911 = lut_tile_10_8_chanxy_out[96];
    assign wire_13912 = lut_tile_10_8_chanxy_out[97];
    assign wire_13913 = lut_tile_10_8_chanxy_out[98];
    assign wire_13914 = lut_tile_10_8_chanxy_out[99];
    assign wire_13915 = lut_tile_10_8_chanxy_out[100];
    assign wire_13916 = lut_tile_10_8_chanxy_out[101];
    assign wire_13917 = lut_tile_10_8_chanxy_out[102];
    assign wire_13918 = lut_tile_10_8_chanxy_out[103];
    assign wire_13919 = lut_tile_10_8_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_9_chanxy_in = {wire_10379, wire_10378, wire_14188, wire_9991, wire_9929, wire_9928, wire_9919, wire_9918, wire_9909, wire_9908, wire_9872, wire_5583, wire_10363, wire_10362, wire_14186, wire_10019, wire_9989, wire_9988, wire_9979, wire_9978, wire_9969, wire_9968, wire_9874, wire_5583, wire_10347, wire_10346, wire_14184, wire_10017, wire_9959, wire_9958, wire_9949, wire_9948, wire_9939, wire_9938, wire_9876, wire_5583, wire_10361, wire_10360, wire_14182, wire_10015, wire_9927, wire_9926, wire_9917, wire_9916, wire_9907, wire_9906, wire_9878, wire_5073, wire_10375, wire_10374, wire_14180, wire_10013, wire_9987, wire_9986, wire_9977, wire_9976, wire_9967, wire_9966, wire_9880, wire_5073, wire_10329, wire_10328, wire_14178, wire_10011, wire_9957, wire_9956, wire_9947, wire_9946, wire_9937, wire_9936, wire_9882, wire_5073, wire_10373, wire_10372, wire_14176, wire_10009, wire_9925, wire_9924, wire_9915, wire_9914, wire_9905, wire_9904, wire_9884, wire_5587, wire_5073, wire_10357, wire_10356, wire_14174, wire_10007, wire_9985, wire_9984, wire_9975, wire_9974, wire_9965, wire_9964, wire_9886, wire_5587, wire_5073, wire_10341, wire_10340, wire_14172, wire_10005, wire_9955, wire_9954, wire_9945, wire_9944, wire_9935, wire_9934, wire_9888, wire_5587, wire_5073, wire_10355, wire_10354, wire_5587, wire_14170, wire_10003, wire_9923, wire_9922, wire_9913, wire_9912, wire_9903, wire_9902, wire_9890, wire_5587, wire_5069, wire_10369, wire_10368, wire_5587, wire_14168, wire_10001, wire_9983, wire_9982, wire_9973, wire_9972, wire_9963, wire_9962, wire_9892, wire_5587, wire_5069, wire_10323, wire_10322, wire_5583, wire_14166, wire_9999, wire_9953, wire_9952, wire_9943, wire_9942, wire_9933, wire_9932, wire_9894, wire_5587, wire_5069, wire_10367, wire_10366, wire_5073, wire_14164, wire_9997, wire_9921, wire_9920, wire_9911, wire_9910, wire_9901, wire_9900, wire_9896, wire_5583, wire_5069, wire_10351, wire_10350, wire_5073, wire_14162, wire_9995, wire_9981, wire_9980, wire_9971, wire_9970, wire_9961, wire_9960, wire_9898, wire_5583, wire_5069, wire_10335, wire_10334, wire_5069, wire_14160, wire_9993, wire_9951, wire_9950, wire_9941, wire_9940, wire_9931, wire_9930, wire_9870, wire_5583, wire_5069, wire_10393, wire_10272, wire_10407, wire_10286, wire_10317, wire_10316, wire_10405, wire_10284, wire_10389, wire_10268, wire_10299, wire_10298, wire_10387, wire_10266, wire_10401, wire_10280, wire_10311, wire_10310, wire_10399, wire_10278, wire_5587, wire_10383, wire_10262, wire_5583, wire_10293, wire_10292, wire_5583, wire_10381, wire_10260, wire_5073, wire_10395, wire_10274, wire_5069, wire_10305, wire_10304, wire_5069, wire_10349, wire_10348, wire_10377, wire_10376, wire_10303, wire_10302, wire_10331, wire_10330, wire_10359, wire_10358, wire_10315, wire_10314, wire_10343, wire_10342, wire_10371, wire_10370, wire_10297, wire_10296, wire_10325, wire_10324, wire_5587, wire_10353, wire_10352, wire_5583, wire_10309, wire_10308, wire_5583, wire_10337, wire_10336, wire_5073, wire_10365, wire_10364, wire_5069, wire_10291, wire_10290, wire_5069, wire_10409, wire_10288, wire_10319, wire_10318, wire_10333, wire_10332, wire_10391, wire_10270, wire_10301, wire_10300, wire_10345, wire_10344, wire_10403, wire_10282, wire_10313, wire_10312, wire_10327, wire_10326, wire_10385, wire_10264, wire_5587, wire_10295, wire_10294, wire_5587, wire_10339, wire_10338, wire_5583, wire_10397, wire_10276, wire_5073, wire_10307, wire_10306, wire_5073, wire_10321, wire_10320, wire_5069, wire_13904, wire_13882, wire_13858, wire_13806, wire_10258, wire_5122, wire_5116, wire_5107, wire_5101, wire_13896, wire_13874, wire_13850, wire_13828, wire_10256, wire_5122, wire_5116, wire_5107, wire_5101, wire_13918, wire_13866, wire_13842, wire_13820, wire_10254, wire_5122, wire_5116, wire_5107, wire_5101, wire_13910, wire_13888, wire_13834, wire_13812, wire_10252, wire_5122, wire_5113, wire_5107, wire_5072, wire_13902, wire_13880, wire_13856, wire_13804, wire_10250, wire_5122, wire_5113, wire_5107, wire_5072, wire_13894, wire_13872, wire_13848, wire_13826, wire_10248, wire_5122, wire_5113, wire_5107, wire_5072, wire_13916, wire_13864, wire_13840, wire_13818, wire_10246, wire_5119, wire_5113, wire_5104, wire_5072, wire_13908, wire_13886, wire_13832, wire_13810, wire_10244, wire_5119, wire_5113, wire_5104, wire_5072, wire_13900, wire_13878, wire_13854, wire_13802, wire_10242, wire_5119, wire_5113, wire_5104, wire_5072, wire_13892, wire_13870, wire_13846, wire_13824, wire_10240, wire_5119, wire_5110, wire_5104, wire_5068, wire_13914, wire_13862, wire_13838, wire_13816, wire_10238, wire_5119, wire_5110, wire_5104, wire_5068, wire_13906, wire_13884, wire_13830, wire_13808, wire_10236, wire_5119, wire_5110, wire_5104, wire_5068, wire_13898, wire_13876, wire_13852, wire_13800, wire_10234, wire_5116, wire_5110, wire_5101, wire_5068, wire_13890, wire_13868, wire_13844, wire_13822, wire_10232, wire_5116, wire_5110, wire_5101, wire_5068, wire_13912, wire_13860, wire_13836, wire_13814, wire_10230, wire_5116, wire_5110, wire_5101, wire_5068, wire_14286, wire_14264, wire_14242, wire_14218, wire_10409, wire_5122, wire_5116, wire_5107, wire_5101, wire_14308, wire_14256, wire_14234, wire_14210, wire_10407, wire_5122, wire_5116, wire_5107, wire_5101, wire_14300, wire_14278, wire_14226, wire_14202, wire_10405, wire_5122, wire_5116, wire_5107, wire_5101, wire_14292, wire_14270, wire_14248, wire_14194, wire_10403, wire_5122, wire_5113, wire_5107, wire_5072, wire_14284, wire_14262, wire_14240, wire_14216, wire_10401, wire_5122, wire_5113, wire_5107, wire_5072, wire_14306, wire_14254, wire_14232, wire_14208, wire_10399, wire_5122, wire_5113, wire_5107, wire_5072, wire_14298, wire_14276, wire_14224, wire_14200, wire_10397, wire_5119, wire_5113, wire_5104, wire_5072, wire_14290, wire_14268, wire_14246, wire_14192, wire_10395, wire_5119, wire_5113, wire_5104, wire_5072, wire_14282, wire_14260, wire_14238, wire_14214, wire_10393, wire_5119, wire_5113, wire_5104, wire_5072, wire_14304, wire_14252, wire_14230, wire_14206, wire_10391, wire_5119, wire_5110, wire_5104, wire_5068, wire_14296, wire_14274, wire_14222, wire_14198, wire_10389, wire_5119, wire_5110, wire_5104, wire_5068, wire_14288, wire_14266, wire_14244, wire_14190, wire_10387, wire_5119, wire_5110, wire_5104, wire_5068, wire_14280, wire_14258, wire_14236, wire_14212, wire_10385, wire_5116, wire_5110, wire_5101, wire_5068, wire_14302, wire_14250, wire_14228, wire_14204, wire_10383, wire_5116, wire_5110, wire_5101, wire_5068, wire_14294, wire_14272, wire_14220, wire_14196, wire_10381, wire_5116, wire_5110, wire_5101, wire_5068};
    // CHNAXY TOTAL: 573
    assign wire_10261 = lut_tile_10_9_chanxy_out[0];
    assign wire_10263 = lut_tile_10_9_chanxy_out[1];
    assign wire_10265 = lut_tile_10_9_chanxy_out[2];
    assign wire_10267 = lut_tile_10_9_chanxy_out[3];
    assign wire_10269 = lut_tile_10_9_chanxy_out[4];
    assign wire_10271 = lut_tile_10_9_chanxy_out[5];
    assign wire_10273 = lut_tile_10_9_chanxy_out[6];
    assign wire_10275 = lut_tile_10_9_chanxy_out[7];
    assign wire_10277 = lut_tile_10_9_chanxy_out[8];
    assign wire_10279 = lut_tile_10_9_chanxy_out[9];
    assign wire_10281 = lut_tile_10_9_chanxy_out[10];
    assign wire_10283 = lut_tile_10_9_chanxy_out[11];
    assign wire_10285 = lut_tile_10_9_chanxy_out[12];
    assign wire_10287 = lut_tile_10_9_chanxy_out[13];
    assign wire_10289 = lut_tile_10_9_chanxy_out[14];
    assign wire_10350 = lut_tile_10_9_chanxy_out[15];
    assign wire_10352 = lut_tile_10_9_chanxy_out[16];
    assign wire_10354 = lut_tile_10_9_chanxy_out[17];
    assign wire_10356 = lut_tile_10_9_chanxy_out[18];
    assign wire_10358 = lut_tile_10_9_chanxy_out[19];
    assign wire_10360 = lut_tile_10_9_chanxy_out[20];
    assign wire_10362 = lut_tile_10_9_chanxy_out[21];
    assign wire_10364 = lut_tile_10_9_chanxy_out[22];
    assign wire_10366 = lut_tile_10_9_chanxy_out[23];
    assign wire_10368 = lut_tile_10_9_chanxy_out[24];
    assign wire_10370 = lut_tile_10_9_chanxy_out[25];
    assign wire_10372 = lut_tile_10_9_chanxy_out[26];
    assign wire_10374 = lut_tile_10_9_chanxy_out[27];
    assign wire_10376 = lut_tile_10_9_chanxy_out[28];
    assign wire_10378 = lut_tile_10_9_chanxy_out[29];
    assign wire_14191 = lut_tile_10_9_chanxy_out[30];
    assign wire_14193 = lut_tile_10_9_chanxy_out[31];
    assign wire_14195 = lut_tile_10_9_chanxy_out[32];
    assign wire_14197 = lut_tile_10_9_chanxy_out[33];
    assign wire_14199 = lut_tile_10_9_chanxy_out[34];
    assign wire_14201 = lut_tile_10_9_chanxy_out[35];
    assign wire_14203 = lut_tile_10_9_chanxy_out[36];
    assign wire_14205 = lut_tile_10_9_chanxy_out[37];
    assign wire_14207 = lut_tile_10_9_chanxy_out[38];
    assign wire_14209 = lut_tile_10_9_chanxy_out[39];
    assign wire_14211 = lut_tile_10_9_chanxy_out[40];
    assign wire_14213 = lut_tile_10_9_chanxy_out[41];
    assign wire_14215 = lut_tile_10_9_chanxy_out[42];
    assign wire_14217 = lut_tile_10_9_chanxy_out[43];
    assign wire_14219 = lut_tile_10_9_chanxy_out[44];
    assign wire_14221 = lut_tile_10_9_chanxy_out[45];
    assign wire_14223 = lut_tile_10_9_chanxy_out[46];
    assign wire_14225 = lut_tile_10_9_chanxy_out[47];
    assign wire_14227 = lut_tile_10_9_chanxy_out[48];
    assign wire_14229 = lut_tile_10_9_chanxy_out[49];
    assign wire_14231 = lut_tile_10_9_chanxy_out[50];
    assign wire_14233 = lut_tile_10_9_chanxy_out[51];
    assign wire_14235 = lut_tile_10_9_chanxy_out[52];
    assign wire_14237 = lut_tile_10_9_chanxy_out[53];
    assign wire_14239 = lut_tile_10_9_chanxy_out[54];
    assign wire_14241 = lut_tile_10_9_chanxy_out[55];
    assign wire_14243 = lut_tile_10_9_chanxy_out[56];
    assign wire_14245 = lut_tile_10_9_chanxy_out[57];
    assign wire_14247 = lut_tile_10_9_chanxy_out[58];
    assign wire_14249 = lut_tile_10_9_chanxy_out[59];
    assign wire_14251 = lut_tile_10_9_chanxy_out[60];
    assign wire_14253 = lut_tile_10_9_chanxy_out[61];
    assign wire_14255 = lut_tile_10_9_chanxy_out[62];
    assign wire_14257 = lut_tile_10_9_chanxy_out[63];
    assign wire_14259 = lut_tile_10_9_chanxy_out[64];
    assign wire_14261 = lut_tile_10_9_chanxy_out[65];
    assign wire_14263 = lut_tile_10_9_chanxy_out[66];
    assign wire_14265 = lut_tile_10_9_chanxy_out[67];
    assign wire_14267 = lut_tile_10_9_chanxy_out[68];
    assign wire_14269 = lut_tile_10_9_chanxy_out[69];
    assign wire_14271 = lut_tile_10_9_chanxy_out[70];
    assign wire_14273 = lut_tile_10_9_chanxy_out[71];
    assign wire_14275 = lut_tile_10_9_chanxy_out[72];
    assign wire_14277 = lut_tile_10_9_chanxy_out[73];
    assign wire_14279 = lut_tile_10_9_chanxy_out[74];
    assign wire_14280 = lut_tile_10_9_chanxy_out[75];
    assign wire_14281 = lut_tile_10_9_chanxy_out[76];
    assign wire_14282 = lut_tile_10_9_chanxy_out[77];
    assign wire_14283 = lut_tile_10_9_chanxy_out[78];
    assign wire_14284 = lut_tile_10_9_chanxy_out[79];
    assign wire_14285 = lut_tile_10_9_chanxy_out[80];
    assign wire_14286 = lut_tile_10_9_chanxy_out[81];
    assign wire_14287 = lut_tile_10_9_chanxy_out[82];
    assign wire_14288 = lut_tile_10_9_chanxy_out[83];
    assign wire_14289 = lut_tile_10_9_chanxy_out[84];
    assign wire_14290 = lut_tile_10_9_chanxy_out[85];
    assign wire_14291 = lut_tile_10_9_chanxy_out[86];
    assign wire_14292 = lut_tile_10_9_chanxy_out[87];
    assign wire_14293 = lut_tile_10_9_chanxy_out[88];
    assign wire_14294 = lut_tile_10_9_chanxy_out[89];
    assign wire_14295 = lut_tile_10_9_chanxy_out[90];
    assign wire_14296 = lut_tile_10_9_chanxy_out[91];
    assign wire_14297 = lut_tile_10_9_chanxy_out[92];
    assign wire_14298 = lut_tile_10_9_chanxy_out[93];
    assign wire_14299 = lut_tile_10_9_chanxy_out[94];
    assign wire_14300 = lut_tile_10_9_chanxy_out[95];
    assign wire_14301 = lut_tile_10_9_chanxy_out[96];
    assign wire_14302 = lut_tile_10_9_chanxy_out[97];
    assign wire_14303 = lut_tile_10_9_chanxy_out[98];
    assign wire_14304 = lut_tile_10_9_chanxy_out[99];
    assign wire_14305 = lut_tile_10_9_chanxy_out[100];
    assign wire_14306 = lut_tile_10_9_chanxy_out[101];
    assign wire_14307 = lut_tile_10_9_chanxy_out[102];
    assign wire_14308 = lut_tile_10_9_chanxy_out[103];
    assign wire_14309 = lut_tile_10_9_chanxy_out[104];
   // CHANXY OUT
    assign lut_tile_10_10_chanxy_in = {wire_10290, wire_6118, wire_14578, wire_9996, wire_9974, wire_9952, wire_9928, wire_6118, wire_6112, wire_6103, wire_6097, wire_10318, wire_6118, wire_14576, wire_10018, wire_9966, wire_9944, wire_9920, wire_6118, wire_6112, wire_6103, wire_6097, wire_10316, wire_6115, wire_14574, wire_10010, wire_9988, wire_9936, wire_9912, wire_6118, wire_6112, wire_6103, wire_6097, wire_10314, wire_6112, wire_14572, wire_10002, wire_9980, wire_9958, wire_9904, wire_6118, wire_6109, wire_6103, wire_5589, wire_10312, wire_6112, wire_14570, wire_9994, wire_9972, wire_9950, wire_9926, wire_6118, wire_6109, wire_6103, wire_5589, wire_10310, wire_6109, wire_14568, wire_10016, wire_9964, wire_9942, wire_9918, wire_6118, wire_6109, wire_6103, wire_5589, wire_10308, wire_6106, wire_14566, wire_10008, wire_9986, wire_9934, wire_9910, wire_6115, wire_6109, wire_6100, wire_5589, wire_10306, wire_6106, wire_14564, wire_10000, wire_9978, wire_9956, wire_9902, wire_6115, wire_6109, wire_6100, wire_5589, wire_10304, wire_6103, wire_14562, wire_9992, wire_9970, wire_9948, wire_9924, wire_6115, wire_6109, wire_6100, wire_5589, wire_10302, wire_6100, wire_14560, wire_10014, wire_9962, wire_9940, wire_9916, wire_6115, wire_6106, wire_6100, wire_5585, wire_10300, wire_6100, wire_14558, wire_10006, wire_9984, wire_9932, wire_9908, wire_6115, wire_6106, wire_6100, wire_5585, wire_10298, wire_6097, wire_14556, wire_9998, wire_9976, wire_9954, wire_9900, wire_6115, wire_6106, wire_6100, wire_5585, wire_10296, wire_5589, wire_14554, wire_9990, wire_9968, wire_9946, wire_9922, wire_6112, wire_6106, wire_6097, wire_5585, wire_10294, wire_5589, wire_14552, wire_10012, wire_9960, wire_9938, wire_9914, wire_6112, wire_6106, wire_6097, wire_5585, wire_10292, wire_5585, wire_14550, wire_10004, wire_9982, wire_9930, wire_9906, wire_6112, wire_6106, wire_6097, wire_5585, wire_10408, wire_6118, wire_10406, wire_6118, wire_10404, wire_6115, wire_10402, wire_6112, wire_10400, wire_6112, wire_10398, wire_6109, wire_10396, wire_6106, wire_10394, wire_6106, wire_10392, wire_6103, wire_10390, wire_6100, wire_10388, wire_6100, wire_10386, wire_6097, wire_10384, wire_5589, wire_10382, wire_5589, wire_10380, wire_5585, wire_10378, wire_6118, wire_10376, wire_6115, wire_10374, wire_6115, wire_10372, wire_6112, wire_10370, wire_6109, wire_10368, wire_6109, wire_10366, wire_6106, wire_10364, wire_6103, wire_10362, wire_6103, wire_10360, wire_6100, wire_10358, wire_6097, wire_10356, wire_6097, wire_10354, wire_5589, wire_10352, wire_5585, wire_10350, wire_5585, wire_10348, wire_6118, wire_10346, wire_6115, wire_10344, wire_6115, wire_10342, wire_6112, wire_10340, wire_6109, wire_10338, wire_6109, wire_10336, wire_6106, wire_10334, wire_6103, wire_10332, wire_6103, wire_10330, wire_6100, wire_10328, wire_6097, wire_10326, wire_6097, wire_10324, wire_5589, wire_10322, wire_5585, wire_10320, wire_5585, wire_14668, wire_5638, wire_14286, wire_14264, wire_14242, wire_14218, wire_10288, wire_5638, wire_5632, wire_5623, wire_5617, wire_14666, wire_5638, wire_14308, wire_14256, wire_14234, wire_14210, wire_10286, wire_5638, wire_5632, wire_5623, wire_5617, wire_14664, wire_5635, wire_14300, wire_14278, wire_14226, wire_14202, wire_10284, wire_5638, wire_5632, wire_5623, wire_5617, wire_14662, wire_5632, wire_14292, wire_14270, wire_14248, wire_14194, wire_10282, wire_5638, wire_5629, wire_5623, wire_5588, wire_14660, wire_5632, wire_14284, wire_14262, wire_14240, wire_14216, wire_10280, wire_5638, wire_5629, wire_5623, wire_5588, wire_14658, wire_5629, wire_14306, wire_14254, wire_14232, wire_14208, wire_10278, wire_5638, wire_5629, wire_5623, wire_5588, wire_14656, wire_5626, wire_14298, wire_14276, wire_14224, wire_14200, wire_10276, wire_5635, wire_5629, wire_5620, wire_5588, wire_14654, wire_5626, wire_14290, wire_14268, wire_14246, wire_14192, wire_10274, wire_5635, wire_5629, wire_5620, wire_5588, wire_14652, wire_5623, wire_14282, wire_14260, wire_14238, wire_14214, wire_10272, wire_5635, wire_5629, wire_5620, wire_5588, wire_14650, wire_5620, wire_14304, wire_14252, wire_14230, wire_14206, wire_10270, wire_5635, wire_5626, wire_5620, wire_5584, wire_14648, wire_5620, wire_14296, wire_14274, wire_14222, wire_14198, wire_10268, wire_5635, wire_5626, wire_5620, wire_5584, wire_14646, wire_5617, wire_14288, wire_14266, wire_14244, wire_14190, wire_10266, wire_5635, wire_5626, wire_5620, wire_5584, wire_14644, wire_5588, wire_14280, wire_14258, wire_14236, wire_14212, wire_10264, wire_5632, wire_5626, wire_5617, wire_5584, wire_14642, wire_5588, wire_14302, wire_14250, wire_14228, wire_14204, wire_10262, wire_5632, wire_5626, wire_5617, wire_5584, wire_14640, wire_5584, wire_14294, wire_14272, wire_14220, wire_14196, wire_10260, wire_5632, wire_5626, wire_5617, wire_5584, wire_14638, wire_5638, wire_14636, wire_5638, wire_14634, wire_5635, wire_14632, wire_5632, wire_14630, wire_5632, wire_14628, wire_5629, wire_14626, wire_5626, wire_14624, wire_5626, wire_14622, wire_5623, wire_14620, wire_5620, wire_14618, wire_5620, wire_14616, wire_5617, wire_14614, wire_5588, wire_14612, wire_5588, wire_14610, wire_5584, wire_14608, wire_5638, wire_14606, wire_5635, wire_14604, wire_5635, wire_14602, wire_5632, wire_14600, wire_5629, wire_14598, wire_5629, wire_14596, wire_5626, wire_14594, wire_5623, wire_14592, wire_5623, wire_14590, wire_5620, wire_14588, wire_5617, wire_14586, wire_5617, wire_14584, wire_5588, wire_14582, wire_5584, wire_14580, wire_5584, wire_14696, wire_5638, wire_14694, wire_5635, wire_14692, wire_5635, wire_14690, wire_5632, wire_14688, wire_5629, wire_14686, wire_5629, wire_14684, wire_5626, wire_14682, wire_5623, wire_14680, wire_5623, wire_14678, wire_5620, wire_14676, wire_5617, wire_14674, wire_5617, wire_14672, wire_5588, wire_14670, wire_5584, wire_14698, wire_5584};
    // CHNAXY TOTAL: 510
    assign wire_10291 = lut_tile_10_10_chanxy_out[0];
    assign wire_10293 = lut_tile_10_10_chanxy_out[1];
    assign wire_10295 = lut_tile_10_10_chanxy_out[2];
    assign wire_10297 = lut_tile_10_10_chanxy_out[3];
    assign wire_10299 = lut_tile_10_10_chanxy_out[4];
    assign wire_10301 = lut_tile_10_10_chanxy_out[5];
    assign wire_10303 = lut_tile_10_10_chanxy_out[6];
    assign wire_10305 = lut_tile_10_10_chanxy_out[7];
    assign wire_10307 = lut_tile_10_10_chanxy_out[8];
    assign wire_10309 = lut_tile_10_10_chanxy_out[9];
    assign wire_10311 = lut_tile_10_10_chanxy_out[10];
    assign wire_10313 = lut_tile_10_10_chanxy_out[11];
    assign wire_10315 = lut_tile_10_10_chanxy_out[12];
    assign wire_10317 = lut_tile_10_10_chanxy_out[13];
    assign wire_10319 = lut_tile_10_10_chanxy_out[14];
    assign wire_10321 = lut_tile_10_10_chanxy_out[15];
    assign wire_10323 = lut_tile_10_10_chanxy_out[16];
    assign wire_10325 = lut_tile_10_10_chanxy_out[17];
    assign wire_10327 = lut_tile_10_10_chanxy_out[18];
    assign wire_10329 = lut_tile_10_10_chanxy_out[19];
    assign wire_10331 = lut_tile_10_10_chanxy_out[20];
    assign wire_10333 = lut_tile_10_10_chanxy_out[21];
    assign wire_10335 = lut_tile_10_10_chanxy_out[22];
    assign wire_10337 = lut_tile_10_10_chanxy_out[23];
    assign wire_10339 = lut_tile_10_10_chanxy_out[24];
    assign wire_10341 = lut_tile_10_10_chanxy_out[25];
    assign wire_10343 = lut_tile_10_10_chanxy_out[26];
    assign wire_10345 = lut_tile_10_10_chanxy_out[27];
    assign wire_10347 = lut_tile_10_10_chanxy_out[28];
    assign wire_10349 = lut_tile_10_10_chanxy_out[29];
    assign wire_10351 = lut_tile_10_10_chanxy_out[30];
    assign wire_10353 = lut_tile_10_10_chanxy_out[31];
    assign wire_10355 = lut_tile_10_10_chanxy_out[32];
    assign wire_10357 = lut_tile_10_10_chanxy_out[33];
    assign wire_10359 = lut_tile_10_10_chanxy_out[34];
    assign wire_10361 = lut_tile_10_10_chanxy_out[35];
    assign wire_10363 = lut_tile_10_10_chanxy_out[36];
    assign wire_10365 = lut_tile_10_10_chanxy_out[37];
    assign wire_10367 = lut_tile_10_10_chanxy_out[38];
    assign wire_10369 = lut_tile_10_10_chanxy_out[39];
    assign wire_10371 = lut_tile_10_10_chanxy_out[40];
    assign wire_10373 = lut_tile_10_10_chanxy_out[41];
    assign wire_10375 = lut_tile_10_10_chanxy_out[42];
    assign wire_10377 = lut_tile_10_10_chanxy_out[43];
    assign wire_10379 = lut_tile_10_10_chanxy_out[44];
    assign wire_10380 = lut_tile_10_10_chanxy_out[45];
    assign wire_10381 = lut_tile_10_10_chanxy_out[46];
    assign wire_10382 = lut_tile_10_10_chanxy_out[47];
    assign wire_10383 = lut_tile_10_10_chanxy_out[48];
    assign wire_10384 = lut_tile_10_10_chanxy_out[49];
    assign wire_10385 = lut_tile_10_10_chanxy_out[50];
    assign wire_10386 = lut_tile_10_10_chanxy_out[51];
    assign wire_10387 = lut_tile_10_10_chanxy_out[52];
    assign wire_10388 = lut_tile_10_10_chanxy_out[53];
    assign wire_10389 = lut_tile_10_10_chanxy_out[54];
    assign wire_10390 = lut_tile_10_10_chanxy_out[55];
    assign wire_10391 = lut_tile_10_10_chanxy_out[56];
    assign wire_10392 = lut_tile_10_10_chanxy_out[57];
    assign wire_10393 = lut_tile_10_10_chanxy_out[58];
    assign wire_10394 = lut_tile_10_10_chanxy_out[59];
    assign wire_10395 = lut_tile_10_10_chanxy_out[60];
    assign wire_10396 = lut_tile_10_10_chanxy_out[61];
    assign wire_10397 = lut_tile_10_10_chanxy_out[62];
    assign wire_10398 = lut_tile_10_10_chanxy_out[63];
    assign wire_10399 = lut_tile_10_10_chanxy_out[64];
    assign wire_10400 = lut_tile_10_10_chanxy_out[65];
    assign wire_10401 = lut_tile_10_10_chanxy_out[66];
    assign wire_10402 = lut_tile_10_10_chanxy_out[67];
    assign wire_10403 = lut_tile_10_10_chanxy_out[68];
    assign wire_10404 = lut_tile_10_10_chanxy_out[69];
    assign wire_10405 = lut_tile_10_10_chanxy_out[70];
    assign wire_10406 = lut_tile_10_10_chanxy_out[71];
    assign wire_10407 = lut_tile_10_10_chanxy_out[72];
    assign wire_10408 = lut_tile_10_10_chanxy_out[73];
    assign wire_10409 = lut_tile_10_10_chanxy_out[74];
    assign wire_14581 = lut_tile_10_10_chanxy_out[75];
    assign wire_14583 = lut_tile_10_10_chanxy_out[76];
    assign wire_14585 = lut_tile_10_10_chanxy_out[77];
    assign wire_14587 = lut_tile_10_10_chanxy_out[78];
    assign wire_14589 = lut_tile_10_10_chanxy_out[79];
    assign wire_14591 = lut_tile_10_10_chanxy_out[80];
    assign wire_14593 = lut_tile_10_10_chanxy_out[81];
    assign wire_14595 = lut_tile_10_10_chanxy_out[82];
    assign wire_14597 = lut_tile_10_10_chanxy_out[83];
    assign wire_14599 = lut_tile_10_10_chanxy_out[84];
    assign wire_14601 = lut_tile_10_10_chanxy_out[85];
    assign wire_14603 = lut_tile_10_10_chanxy_out[86];
    assign wire_14605 = lut_tile_10_10_chanxy_out[87];
    assign wire_14607 = lut_tile_10_10_chanxy_out[88];
    assign wire_14609 = lut_tile_10_10_chanxy_out[89];
    assign wire_14611 = lut_tile_10_10_chanxy_out[90];
    assign wire_14613 = lut_tile_10_10_chanxy_out[91];
    assign wire_14615 = lut_tile_10_10_chanxy_out[92];
    assign wire_14617 = lut_tile_10_10_chanxy_out[93];
    assign wire_14619 = lut_tile_10_10_chanxy_out[94];
    assign wire_14621 = lut_tile_10_10_chanxy_out[95];
    assign wire_14623 = lut_tile_10_10_chanxy_out[96];
    assign wire_14625 = lut_tile_10_10_chanxy_out[97];
    assign wire_14627 = lut_tile_10_10_chanxy_out[98];
    assign wire_14629 = lut_tile_10_10_chanxy_out[99];
    assign wire_14631 = lut_tile_10_10_chanxy_out[100];
    assign wire_14633 = lut_tile_10_10_chanxy_out[101];
    assign wire_14635 = lut_tile_10_10_chanxy_out[102];
    assign wire_14637 = lut_tile_10_10_chanxy_out[103];
    assign wire_14639 = lut_tile_10_10_chanxy_out[104];
    assign wire_14641 = lut_tile_10_10_chanxy_out[105];
    assign wire_14643 = lut_tile_10_10_chanxy_out[106];
    assign wire_14645 = lut_tile_10_10_chanxy_out[107];
    assign wire_14647 = lut_tile_10_10_chanxy_out[108];
    assign wire_14649 = lut_tile_10_10_chanxy_out[109];
    assign wire_14651 = lut_tile_10_10_chanxy_out[110];
    assign wire_14653 = lut_tile_10_10_chanxy_out[111];
    assign wire_14655 = lut_tile_10_10_chanxy_out[112];
    assign wire_14657 = lut_tile_10_10_chanxy_out[113];
    assign wire_14659 = lut_tile_10_10_chanxy_out[114];
    assign wire_14661 = lut_tile_10_10_chanxy_out[115];
    assign wire_14663 = lut_tile_10_10_chanxy_out[116];
    assign wire_14665 = lut_tile_10_10_chanxy_out[117];
    assign wire_14667 = lut_tile_10_10_chanxy_out[118];
    assign wire_14669 = lut_tile_10_10_chanxy_out[119];
    assign wire_14670 = lut_tile_10_10_chanxy_out[120];
    assign wire_14671 = lut_tile_10_10_chanxy_out[121];
    assign wire_14672 = lut_tile_10_10_chanxy_out[122];
    assign wire_14673 = lut_tile_10_10_chanxy_out[123];
    assign wire_14674 = lut_tile_10_10_chanxy_out[124];
    assign wire_14675 = lut_tile_10_10_chanxy_out[125];
    assign wire_14676 = lut_tile_10_10_chanxy_out[126];
    assign wire_14677 = lut_tile_10_10_chanxy_out[127];
    assign wire_14678 = lut_tile_10_10_chanxy_out[128];
    assign wire_14679 = lut_tile_10_10_chanxy_out[129];
    assign wire_14680 = lut_tile_10_10_chanxy_out[130];
    assign wire_14681 = lut_tile_10_10_chanxy_out[131];
    assign wire_14682 = lut_tile_10_10_chanxy_out[132];
    assign wire_14683 = lut_tile_10_10_chanxy_out[133];
    assign wire_14684 = lut_tile_10_10_chanxy_out[134];
    assign wire_14685 = lut_tile_10_10_chanxy_out[135];
    assign wire_14686 = lut_tile_10_10_chanxy_out[136];
    assign wire_14687 = lut_tile_10_10_chanxy_out[137];
    assign wire_14688 = lut_tile_10_10_chanxy_out[138];
    assign wire_14689 = lut_tile_10_10_chanxy_out[139];
    assign wire_14690 = lut_tile_10_10_chanxy_out[140];
    assign wire_14691 = lut_tile_10_10_chanxy_out[141];
    assign wire_14692 = lut_tile_10_10_chanxy_out[142];
    assign wire_14693 = lut_tile_10_10_chanxy_out[143];
    assign wire_14694 = lut_tile_10_10_chanxy_out[144];
    assign wire_14695 = lut_tile_10_10_chanxy_out[145];
    assign wire_14696 = lut_tile_10_10_chanxy_out[146];
    assign wire_14697 = lut_tile_10_10_chanxy_out[147];
    assign wire_14698 = lut_tile_10_10_chanxy_out[148];
    assign wire_14699 = lut_tile_10_10_chanxy_out[149];
   // CHANXY OUT
    // FPGA IO IPIN
    assign io_tile_1_0_ipin_in = {wire_10529, wire_10528, wire_10509, wire_10508, wire_10489, wire_10488, wire_10469, wire_10468, wire_10449, wire_10448, wire_10429, wire_10428, wire_10525, wire_10524, wire_10505, wire_10504, wire_10485, wire_10484, wire_10465, wire_10464, wire_10445, wire_10444, wire_10425, wire_10424, wire_10523, wire_10522, wire_10503, wire_10502, wire_10483, wire_10482, wire_10463, wire_10462, wire_10443, wire_10442, wire_10423, wire_10422, wire_10521, wire_10520, wire_10501, wire_10500, wire_10481, wire_10480, wire_10461, wire_10460, wire_10441, wire_10440, wire_10421, wire_10420, wire_10519, wire_10518, wire_10499, wire_10498, wire_10479, wire_10478, wire_10459, wire_10458, wire_10439, wire_10438, wire_10419, wire_10418, wire_10515, wire_10514, wire_10495, wire_10494, wire_10475, wire_10474, wire_10455, wire_10454, wire_10435, wire_10434, wire_10415, wire_10414, wire_10513, wire_10512, wire_10493, wire_10492, wire_10473, wire_10472, wire_10453, wire_10452, wire_10433, wire_10432, wire_10413, wire_10412, wire_10511, wire_10510, wire_10491, wire_10490, wire_10471, wire_10470, wire_10451, wire_10450, wire_10431, wire_10430, wire_10411, wire_10410};
    // FPGA IPIN IN
    assign io_tile_2_0_ipin_in = {wire_10527, wire_10526, wire_10507, wire_10506, wire_10487, wire_10486, wire_10467, wire_10466, wire_10447, wire_10446, wire_10427, wire_10426, wire_10523, wire_10522, wire_10503, wire_10502, wire_10483, wire_10482, wire_10463, wire_10462, wire_10443, wire_10442, wire_10423, wire_10422, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_10529, wire_10528, wire_10489, wire_10488, wire_10449, wire_10448, wire_10519, wire_10518, wire_10499, wire_10498, wire_10479, wire_10478, wire_10459, wire_10458, wire_10439, wire_10438, wire_10419, wire_10418, wire_10557, wire_10556, wire_10547, wire_10546, wire_10537, wire_10536, wire_10505, wire_10504, wire_10465, wire_10464, wire_10425, wire_10424, wire_10551, wire_10550, wire_10541, wire_10540, wire_10531, wire_10530, wire_10521, wire_10520, wire_10481, wire_10480, wire_10441, wire_10440, wire_10511, wire_10510, wire_10491, wire_10490, wire_10471, wire_10470, wire_10451, wire_10450, wire_10431, wire_10430, wire_10411, wire_10410, wire_10555, wire_10554, wire_10545, wire_10544, wire_10535, wire_10534, wire_10497, wire_10496, wire_10457, wire_10456, wire_10417, wire_10416};
    // FPGA IPIN IN
    assign io_tile_3_0_ipin_in = {wire_10559, wire_10558, wire_10549, wire_10548, wire_10539, wire_10538, wire_10513, wire_10512, wire_10473, wire_10472, wire_10433, wire_10432, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_10529, wire_10528, wire_10489, wire_10488, wire_10449, wire_10448, wire_10589, wire_10588, wire_10579, wire_10578, wire_10569, wire_10568, wire_10499, wire_10498, wire_10459, wire_10458, wire_10419, wire_10418, wire_10557, wire_10556, wire_10547, wire_10546, wire_10537, wire_10536, wire_10505, wire_10504, wire_10465, wire_10464, wire_10425, wire_10424, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_10515, wire_10514, wire_10475, wire_10474, wire_10435, wire_10434, wire_10587, wire_10586, wire_10577, wire_10576, wire_10567, wire_10566, wire_10491, wire_10490, wire_10451, wire_10450, wire_10411, wire_10410, wire_10555, wire_10554, wire_10545, wire_10544, wire_10535, wire_10534, wire_10497, wire_10496, wire_10457, wire_10456, wire_10417, wire_10416, wire_10581, wire_10580, wire_10571, wire_10570, wire_10561, wire_10560, wire_10507, wire_10506, wire_10467, wire_10466, wire_10427, wire_10426};
    // FPGA IPIN IN
    assign io_tile_4_0_ipin_in = {wire_10585, wire_10584, wire_10575, wire_10574, wire_10565, wire_10564, wire_10523, wire_10522, wire_10483, wire_10482, wire_10443, wire_10442, wire_10589, wire_10588, wire_10579, wire_10578, wire_10569, wire_10568, wire_10499, wire_10498, wire_10459, wire_10458, wire_10419, wire_10418, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_10559, wire_10558, wire_10549, wire_10548, wire_10539, wire_10538, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_10515, wire_10514, wire_10475, wire_10474, wire_10435, wire_10434, wire_10617, wire_10616, wire_10607, wire_10606, wire_10597, wire_10596, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_10611, wire_10610, wire_10601, wire_10600, wire_10591, wire_10590, wire_10557, wire_10556, wire_10547, wire_10546, wire_10537, wire_10536, wire_10581, wire_10580, wire_10571, wire_10570, wire_10561, wire_10560, wire_10507, wire_10506, wire_10467, wire_10466, wire_10427, wire_10426, wire_10615, wire_10614, wire_10605, wire_10604, wire_10595, wire_10594, wire_10551, wire_10550, wire_10541, wire_10540, wire_10531, wire_10530};
    // FPGA IPIN IN
    assign io_tile_5_0_ipin_in = {wire_10619, wire_10618, wire_10609, wire_10608, wire_10599, wire_10598, wire_10555, wire_10554, wire_10545, wire_10544, wire_10535, wire_10534, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_10559, wire_10558, wire_10549, wire_10548, wire_10539, wire_10538, wire_10649, wire_10648, wire_10639, wire_10638, wire_10629, wire_10628, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_10617, wire_10616, wire_10607, wire_10606, wire_10597, wire_10596, wire_10553, wire_10552, wire_10543, wire_10542, wire_10533, wire_10532, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_10587, wire_10586, wire_10577, wire_10576, wire_10567, wire_10566, wire_10647, wire_10646, wire_10637, wire_10636, wire_10627, wire_10626, wire_10581, wire_10580, wire_10571, wire_10570, wire_10561, wire_10560, wire_10615, wire_10614, wire_10605, wire_10604, wire_10595, wire_10594, wire_10551, wire_10550, wire_10541, wire_10540, wire_10531, wire_10530, wire_10641, wire_10640, wire_10631, wire_10630, wire_10621, wire_10620, wire_10585, wire_10584, wire_10575, wire_10574, wire_10565, wire_10564};
    // FPGA IPIN IN
    assign io_tile_6_0_ipin_in = {wire_10645, wire_10644, wire_10635, wire_10634, wire_10625, wire_10624, wire_10589, wire_10588, wire_10579, wire_10578, wire_10569, wire_10568, wire_10649, wire_10648, wire_10639, wire_10638, wire_10629, wire_10628, wire_10583, wire_10582, wire_10573, wire_10572, wire_10563, wire_10562, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_10619, wire_10618, wire_10609, wire_10608, wire_10599, wire_10598, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_10587, wire_10586, wire_10577, wire_10576, wire_10567, wire_10566, wire_10677, wire_10676, wire_10667, wire_10666, wire_10657, wire_10656, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_10671, wire_10670, wire_10661, wire_10660, wire_10651, wire_10650, wire_10617, wire_10616, wire_10607, wire_10606, wire_10597, wire_10596, wire_10641, wire_10640, wire_10631, wire_10630, wire_10621, wire_10620, wire_10585, wire_10584, wire_10575, wire_10574, wire_10565, wire_10564, wire_10675, wire_10674, wire_10665, wire_10664, wire_10655, wire_10654, wire_10611, wire_10610, wire_10601, wire_10600, wire_10591, wire_10590};
    // FPGA IPIN IN
    assign io_tile_7_0_ipin_in = {wire_10679, wire_10678, wire_10669, wire_10668, wire_10659, wire_10658, wire_10615, wire_10614, wire_10605, wire_10604, wire_10595, wire_10594, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_10619, wire_10618, wire_10609, wire_10608, wire_10599, wire_10598, wire_10709, wire_10708, wire_10699, wire_10698, wire_10689, wire_10688, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_10677, wire_10676, wire_10667, wire_10666, wire_10657, wire_10656, wire_10613, wire_10612, wire_10603, wire_10602, wire_10593, wire_10592, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_10647, wire_10646, wire_10637, wire_10636, wire_10627, wire_10626, wire_10707, wire_10706, wire_10697, wire_10696, wire_10687, wire_10686, wire_10641, wire_10640, wire_10631, wire_10630, wire_10621, wire_10620, wire_10675, wire_10674, wire_10665, wire_10664, wire_10655, wire_10654, wire_10611, wire_10610, wire_10601, wire_10600, wire_10591, wire_10590, wire_10701, wire_10700, wire_10691, wire_10690, wire_10681, wire_10680, wire_10645, wire_10644, wire_10635, wire_10634, wire_10625, wire_10624};
    // FPGA IPIN IN
    assign io_tile_8_0_ipin_in = {wire_10705, wire_10704, wire_10695, wire_10694, wire_10685, wire_10684, wire_10649, wire_10648, wire_10639, wire_10638, wire_10629, wire_10628, wire_10709, wire_10708, wire_10699, wire_10698, wire_10689, wire_10688, wire_10643, wire_10642, wire_10633, wire_10632, wire_10623, wire_10622, wire_10733, wire_10732, wire_10723, wire_10722, wire_10713, wire_10712, wire_10679, wire_10678, wire_10669, wire_10668, wire_10659, wire_10658, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_10647, wire_10646, wire_10637, wire_10636, wire_10627, wire_10626, wire_10737, wire_10736, wire_10727, wire_10726, wire_10717, wire_10716, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_10731, wire_10730, wire_10721, wire_10720, wire_10711, wire_10710, wire_10677, wire_10676, wire_10667, wire_10666, wire_10657, wire_10656, wire_10701, wire_10700, wire_10691, wire_10690, wire_10681, wire_10680, wire_10645, wire_10644, wire_10635, wire_10634, wire_10625, wire_10624, wire_10735, wire_10734, wire_10725, wire_10724, wire_10715, wire_10714, wire_10671, wire_10670, wire_10661, wire_10660, wire_10651, wire_10650};
    // FPGA IPIN IN
    assign io_tile_9_0_ipin_in = {wire_10739, wire_10738, wire_10729, wire_10728, wire_10719, wire_10718, wire_10675, wire_10674, wire_10665, wire_10664, wire_10655, wire_10654, wire_10733, wire_10732, wire_10723, wire_10722, wire_10713, wire_10712, wire_10679, wire_10678, wire_10669, wire_10668, wire_10659, wire_10658, wire_10769, wire_10768, wire_10759, wire_10758, wire_10749, wire_10748, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_10737, wire_10736, wire_10727, wire_10726, wire_10717, wire_10716, wire_10673, wire_10672, wire_10663, wire_10662, wire_10653, wire_10652, wire_10763, wire_10762, wire_10753, wire_10752, wire_10743, wire_10742, wire_10707, wire_10706, wire_10697, wire_10696, wire_10687, wire_10686, wire_10767, wire_10766, wire_10757, wire_10756, wire_10747, wire_10746, wire_10701, wire_10700, wire_10691, wire_10690, wire_10681, wire_10680, wire_10735, wire_10734, wire_10725, wire_10724, wire_10715, wire_10714, wire_10671, wire_10670, wire_10661, wire_10660, wire_10651, wire_10650, wire_10761, wire_10760, wire_10751, wire_10750, wire_10741, wire_10740, wire_10705, wire_10704, wire_10695, wire_10694, wire_10685, wire_10684};
    // FPGA IPIN IN
    assign io_tile_10_0_ipin_in = {wire_10765, wire_10764, wire_10755, wire_10754, wire_10745, wire_10744, wire_10709, wire_10708, wire_10699, wire_10698, wire_10689, wire_10688, wire_10769, wire_10768, wire_10759, wire_10758, wire_10749, wire_10748, wire_10703, wire_10702, wire_10693, wire_10692, wire_10683, wire_10682, wire_10793, wire_10792, wire_10783, wire_10782, wire_10773, wire_10772, wire_10739, wire_10738, wire_10729, wire_10728, wire_10719, wire_10718, wire_10763, wire_10762, wire_10753, wire_10752, wire_10743, wire_10742, wire_10707, wire_10706, wire_10697, wire_10696, wire_10687, wire_10686, wire_10797, wire_10796, wire_10787, wire_10786, wire_10777, wire_10776, wire_10733, wire_10732, wire_10723, wire_10722, wire_10713, wire_10712, wire_10791, wire_10790, wire_10781, wire_10780, wire_10771, wire_10770, wire_10737, wire_10736, wire_10727, wire_10726, wire_10717, wire_10716, wire_10761, wire_10760, wire_10751, wire_10750, wire_10741, wire_10740, wire_10705, wire_10704, wire_10695, wire_10694, wire_10685, wire_10684, wire_10795, wire_10794, wire_10785, wire_10784, wire_10775, wire_10774, wire_10731, wire_10730, wire_10721, wire_10720, wire_10711, wire_10710};
    // FPGA IPIN IN
    assign io_tile_1_11_ipin_in = {wire_14425, wire_14424, wire_14413, wire_14412, wire_14385, wire_14384, wire_14373, wire_14372, wire_14345, wire_14344, wire_14333, wire_14332, wire_14423, wire_14422, wire_14411, wire_14410, wire_14383, wire_14382, wire_14371, wire_14370, wire_14343, wire_14342, wire_14331, wire_14330, wire_14429, wire_14428, wire_14401, wire_14400, wire_14389, wire_14388, wire_14361, wire_14360, wire_14349, wire_14348, wire_14321, wire_14320, wire_14417, wire_14416, wire_14405, wire_14404, wire_14377, wire_14376, wire_14365, wire_14364, wire_14337, wire_14336, wire_14325, wire_14324, wire_14415, wire_14414, wire_14403, wire_14402, wire_14375, wire_14374, wire_14363, wire_14362, wire_14335, wire_14334, wire_14323, wire_14322, wire_14421, wire_14420, wire_14393, wire_14392, wire_14381, wire_14380, wire_14353, wire_14352, wire_14341, wire_14340, wire_14313, wire_14312, wire_14419, wire_14418, wire_14391, wire_14390, wire_14379, wire_14378, wire_14351, wire_14350, wire_14339, wire_14338, wire_14311, wire_14310, wire_14407, wire_14406, wire_14395, wire_14394, wire_14367, wire_14366, wire_14355, wire_14354, wire_14327, wire_14326, wire_14315, wire_14314};
    // FPGA IPIN IN
    assign io_tile_2_11_ipin_in = {wire_14423, wire_14422, wire_14411, wire_14410, wire_14383, wire_14382, wire_14371, wire_14370, wire_14343, wire_14342, wire_14331, wire_14330, wire_14459, wire_14458, wire_14449, wire_14448, wire_14439, wire_14438, wire_14409, wire_14408, wire_14369, wire_14368, wire_14329, wire_14328, wire_14427, wire_14426, wire_14399, wire_14398, wire_14387, wire_14386, wire_14359, wire_14358, wire_14347, wire_14346, wire_14319, wire_14318, wire_14415, wire_14414, wire_14403, wire_14402, wire_14375, wire_14374, wire_14363, wire_14362, wire_14335, wire_14334, wire_14323, wire_14322, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_14401, wire_14400, wire_14361, wire_14360, wire_14321, wire_14320, wire_14419, wire_14418, wire_14391, wire_14390, wire_14379, wire_14378, wire_14351, wire_14350, wire_14339, wire_14338, wire_14311, wire_14310, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430, wire_14417, wire_14416, wire_14377, wire_14376, wire_14337, wire_14336, wire_14455, wire_14454, wire_14445, wire_14444, wire_14435, wire_14434, wire_14393, wire_14392, wire_14353, wire_14352, wire_14313, wire_14312};
    // FPGA IPIN IN
    assign io_tile_3_11_ipin_in = {wire_14459, wire_14458, wire_14449, wire_14448, wire_14439, wire_14438, wire_14409, wire_14408, wire_14369, wire_14368, wire_14329, wire_14328, wire_14485, wire_14484, wire_14475, wire_14474, wire_14465, wire_14464, wire_14427, wire_14426, wire_14387, wire_14386, wire_14347, wire_14346, wire_14453, wire_14452, wire_14443, wire_14442, wire_14433, wire_14432, wire_14425, wire_14424, wire_14385, wire_14384, wire_14345, wire_14344, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_14401, wire_14400, wire_14361, wire_14360, wire_14321, wire_14320, wire_14483, wire_14482, wire_14473, wire_14472, wire_14463, wire_14462, wire_14419, wire_14418, wire_14379, wire_14378, wire_14339, wire_14338, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430, wire_14417, wire_14416, wire_14377, wire_14376, wire_14337, wire_14336, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14395, wire_14394, wire_14355, wire_14354, wire_14315, wire_14314, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_14411, wire_14410, wire_14371, wire_14370, wire_14331, wire_14330};
    // FPGA IPIN IN
    assign io_tile_4_11_ipin_in = {wire_14485, wire_14484, wire_14475, wire_14474, wire_14465, wire_14464, wire_14427, wire_14426, wire_14387, wire_14386, wire_14347, wire_14346, wire_14519, wire_14518, wire_14509, wire_14508, wire_14499, wire_14498, wire_14455, wire_14454, wire_14445, wire_14444, wire_14435, wire_14434, wire_14489, wire_14488, wire_14479, wire_14478, wire_14469, wire_14468, wire_14403, wire_14402, wire_14363, wire_14362, wire_14323, wire_14322, wire_14483, wire_14482, wire_14473, wire_14472, wire_14463, wire_14462, wire_14419, wire_14418, wire_14379, wire_14378, wire_14339, wire_14338, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_14453, wire_14452, wire_14443, wire_14442, wire_14433, wire_14432, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14395, wire_14394, wire_14355, wire_14354, wire_14315, wire_14314, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_14515, wire_14514, wire_14505, wire_14504, wire_14495, wire_14494, wire_14451, wire_14450, wire_14441, wire_14440, wire_14431, wire_14430};
    // FPGA IPIN IN
    assign io_tile_5_11_ipin_in = {wire_14519, wire_14518, wire_14509, wire_14508, wire_14499, wire_14498, wire_14455, wire_14454, wire_14445, wire_14444, wire_14435, wire_14434, wire_14545, wire_14544, wire_14535, wire_14534, wire_14525, wire_14524, wire_14489, wire_14488, wire_14479, wire_14478, wire_14469, wire_14468, wire_14513, wire_14512, wire_14503, wire_14502, wire_14493, wire_14492, wire_14459, wire_14458, wire_14449, wire_14448, wire_14439, wire_14438, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_14453, wire_14452, wire_14443, wire_14442, wire_14433, wire_14432, wire_14543, wire_14542, wire_14533, wire_14532, wire_14523, wire_14522, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490, wire_14457, wire_14456, wire_14447, wire_14446, wire_14437, wire_14436, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_14485, wire_14484, wire_14475, wire_14474, wire_14465, wire_14464};
    // FPGA IPIN IN
    assign io_tile_6_11_ipin_in = {wire_14545, wire_14544, wire_14535, wire_14534, wire_14525, wire_14524, wire_14489, wire_14488, wire_14479, wire_14478, wire_14469, wire_14468, wire_14579, wire_14578, wire_14569, wire_14568, wire_14559, wire_14558, wire_14515, wire_14514, wire_14505, wire_14504, wire_14495, wire_14494, wire_14549, wire_14548, wire_14539, wire_14538, wire_14529, wire_14528, wire_14483, wire_14482, wire_14473, wire_14472, wire_14463, wire_14462, wire_14543, wire_14542, wire_14533, wire_14532, wire_14523, wire_14522, wire_14487, wire_14486, wire_14477, wire_14476, wire_14467, wire_14466, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_14513, wire_14512, wire_14503, wire_14502, wire_14493, wire_14492, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14481, wire_14480, wire_14471, wire_14470, wire_14461, wire_14460, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_14575, wire_14574, wire_14565, wire_14564, wire_14555, wire_14554, wire_14511, wire_14510, wire_14501, wire_14500, wire_14491, wire_14490};
    // FPGA IPIN IN
    assign io_tile_7_11_ipin_in = {wire_14579, wire_14578, wire_14569, wire_14568, wire_14559, wire_14558, wire_14515, wire_14514, wire_14505, wire_14504, wire_14495, wire_14494, wire_14605, wire_14604, wire_14595, wire_14594, wire_14585, wire_14584, wire_14549, wire_14548, wire_14539, wire_14538, wire_14529, wire_14528, wire_14573, wire_14572, wire_14563, wire_14562, wire_14553, wire_14552, wire_14519, wire_14518, wire_14509, wire_14508, wire_14499, wire_14498, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_14513, wire_14512, wire_14503, wire_14502, wire_14493, wire_14492, wire_14603, wire_14602, wire_14593, wire_14592, wire_14583, wire_14582, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550, wire_14517, wire_14516, wire_14507, wire_14506, wire_14497, wire_14496, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_14545, wire_14544, wire_14535, wire_14534, wire_14525, wire_14524};
    // FPGA IPIN IN
    assign io_tile_8_11_ipin_in = {wire_14605, wire_14604, wire_14595, wire_14594, wire_14585, wire_14584, wire_14549, wire_14548, wire_14539, wire_14538, wire_14529, wire_14528, wire_14639, wire_14638, wire_14629, wire_14628, wire_14619, wire_14618, wire_14575, wire_14574, wire_14565, wire_14564, wire_14555, wire_14554, wire_14609, wire_14608, wire_14599, wire_14598, wire_14589, wire_14588, wire_14543, wire_14542, wire_14533, wire_14532, wire_14523, wire_14522, wire_14603, wire_14602, wire_14593, wire_14592, wire_14583, wire_14582, wire_14547, wire_14546, wire_14537, wire_14536, wire_14527, wire_14526, wire_14637, wire_14636, wire_14627, wire_14626, wire_14617, wire_14616, wire_14573, wire_14572, wire_14563, wire_14562, wire_14553, wire_14552, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14541, wire_14540, wire_14531, wire_14530, wire_14521, wire_14520, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_14635, wire_14634, wire_14625, wire_14624, wire_14615, wire_14614, wire_14571, wire_14570, wire_14561, wire_14560, wire_14551, wire_14550};
    // FPGA IPIN IN
    assign io_tile_9_11_ipin_in = {wire_14639, wire_14638, wire_14629, wire_14628, wire_14619, wire_14618, wire_14575, wire_14574, wire_14565, wire_14564, wire_14555, wire_14554, wire_14665, wire_14664, wire_14655, wire_14654, wire_14645, wire_14644, wire_14609, wire_14608, wire_14599, wire_14598, wire_14589, wire_14588, wire_14633, wire_14632, wire_14623, wire_14622, wire_14613, wire_14612, wire_14579, wire_14578, wire_14569, wire_14568, wire_14559, wire_14558, wire_14637, wire_14636, wire_14627, wire_14626, wire_14617, wire_14616, wire_14573, wire_14572, wire_14563, wire_14562, wire_14553, wire_14552, wire_14663, wire_14662, wire_14653, wire_14652, wire_14643, wire_14642, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610, wire_14577, wire_14576, wire_14567, wire_14566, wire_14557, wire_14556, wire_14667, wire_14666, wire_14657, wire_14656, wire_14647, wire_14646, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_14661, wire_14660, wire_14651, wire_14650, wire_14641, wire_14640, wire_14605, wire_14604, wire_14595, wire_14594, wire_14585, wire_14584};
    // FPGA IPIN IN
    assign io_tile_10_11_ipin_in = {wire_14665, wire_14664, wire_14655, wire_14654, wire_14645, wire_14644, wire_14609, wire_14608, wire_14599, wire_14598, wire_14589, wire_14588, wire_14699, wire_14698, wire_14689, wire_14688, wire_14679, wire_14678, wire_14635, wire_14634, wire_14625, wire_14624, wire_14615, wire_14614, wire_14669, wire_14668, wire_14659, wire_14658, wire_14649, wire_14648, wire_14603, wire_14602, wire_14593, wire_14592, wire_14583, wire_14582, wire_14663, wire_14662, wire_14653, wire_14652, wire_14643, wire_14642, wire_14607, wire_14606, wire_14597, wire_14596, wire_14587, wire_14586, wire_14697, wire_14696, wire_14687, wire_14686, wire_14677, wire_14676, wire_14633, wire_14632, wire_14623, wire_14622, wire_14613, wire_14612, wire_14667, wire_14666, wire_14657, wire_14656, wire_14647, wire_14646, wire_14601, wire_14600, wire_14591, wire_14590, wire_14581, wire_14580, wire_14691, wire_14690, wire_14681, wire_14680, wire_14671, wire_14670, wire_14637, wire_14636, wire_14627, wire_14626, wire_14617, wire_14616, wire_14695, wire_14694, wire_14685, wire_14684, wire_14675, wire_14674, wire_14631, wire_14630, wire_14621, wire_14620, wire_14611, wire_14610};
    // FPGA IPIN IN
    assign io_tile_0_1_ipin_in = {wire_6237, wire_6236, wire_6217, wire_6216, wire_6197, wire_6196, wire_6177, wire_6176, wire_6157, wire_6156, wire_6137, wire_6136, wire_6235, wire_6234, wire_6215, wire_6214, wire_6195, wire_6194, wire_6175, wire_6174, wire_6155, wire_6154, wire_6135, wire_6134, wire_6233, wire_6232, wire_6213, wire_6212, wire_6193, wire_6192, wire_6173, wire_6172, wire_6153, wire_6152, wire_6133, wire_6132, wire_6231, wire_6230, wire_6211, wire_6210, wire_6191, wire_6190, wire_6171, wire_6170, wire_6151, wire_6150, wire_6131, wire_6130, wire_6227, wire_6226, wire_6207, wire_6206, wire_6187, wire_6186, wire_6167, wire_6166, wire_6147, wire_6146, wire_6127, wire_6126, wire_6225, wire_6224, wire_6205, wire_6204, wire_6185, wire_6184, wire_6165, wire_6164, wire_6145, wire_6144, wire_6125, wire_6124, wire_6223, wire_6222, wire_6203, wire_6202, wire_6183, wire_6182, wire_6163, wire_6162, wire_6143, wire_6142, wire_6123, wire_6122, wire_6221, wire_6220, wire_6201, wire_6200, wire_6181, wire_6180, wire_6161, wire_6160, wire_6141, wire_6140, wire_6121, wire_6120};
    // FPGA IPIN IN
    assign io_tile_0_2_ipin_in = {wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_6223, wire_6222, wire_6183, wire_6182, wire_6143, wire_6142, wire_6233, wire_6232, wire_6213, wire_6212, wire_6193, wire_6192, wire_6173, wire_6172, wire_6153, wire_6152, wire_6133, wire_6132, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_6239, wire_6238, wire_6199, wire_6198, wire_6159, wire_6158, wire_6229, wire_6228, wire_6209, wire_6208, wire_6189, wire_6188, wire_6169, wire_6168, wire_6149, wire_6148, wire_6129, wire_6128, wire_6225, wire_6224, wire_6205, wire_6204, wire_6185, wire_6184, wire_6165, wire_6164, wire_6145, wire_6144, wire_6125, wire_6124, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240, wire_6231, wire_6230, wire_6191, wire_6190, wire_6151, wire_6150, wire_6221, wire_6220, wire_6201, wire_6200, wire_6181, wire_6180, wire_6161, wire_6160, wire_6141, wire_6140, wire_6121, wire_6120, wire_6265, wire_6264, wire_6255, wire_6254, wire_6245, wire_6244, wire_6207, wire_6206, wire_6167, wire_6166, wire_6127, wire_6126};
    // FPGA IPIN IN
    assign io_tile_0_3_ipin_in = {wire_6295, wire_6294, wire_6285, wire_6284, wire_6275, wire_6274, wire_6233, wire_6232, wire_6193, wire_6192, wire_6153, wire_6152, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_6239, wire_6238, wire_6199, wire_6198, wire_6159, wire_6158, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_6209, wire_6208, wire_6169, wire_6168, wire_6129, wire_6128, wire_6267, wire_6266, wire_6257, wire_6256, wire_6247, wire_6246, wire_6215, wire_6214, wire_6175, wire_6174, wire_6135, wire_6134, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240, wire_6231, wire_6230, wire_6191, wire_6190, wire_6151, wire_6150, wire_6297, wire_6296, wire_6287, wire_6286, wire_6277, wire_6276, wire_6201, wire_6200, wire_6161, wire_6160, wire_6121, wire_6120, wire_6265, wire_6264, wire_6255, wire_6254, wire_6245, wire_6244, wire_6207, wire_6206, wire_6167, wire_6166, wire_6127, wire_6126, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_6217, wire_6216, wire_6177, wire_6176, wire_6137, wire_6136};
    // FPGA IPIN IN
    assign io_tile_0_4_ipin_in = {wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_6265, wire_6264, wire_6255, wire_6254, wire_6245, wire_6244, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_6209, wire_6208, wire_6169, wire_6168, wire_6129, wire_6128, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_6225, wire_6224, wire_6185, wire_6184, wire_6145, wire_6144, wire_6297, wire_6296, wire_6287, wire_6286, wire_6277, wire_6276, wire_6201, wire_6200, wire_6161, wire_6160, wire_6121, wire_6120, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300, wire_6267, wire_6266, wire_6257, wire_6256, wire_6247, wire_6246, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_6217, wire_6216, wire_6177, wire_6176, wire_6137, wire_6136, wire_6325, wire_6324, wire_6315, wire_6314, wire_6305, wire_6304, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240};
    // FPGA IPIN IN
    assign io_tile_0_5_ipin_in = {wire_6355, wire_6354, wire_6345, wire_6344, wire_6335, wire_6334, wire_6299, wire_6298, wire_6289, wire_6288, wire_6279, wire_6278, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_6269, wire_6268, wire_6259, wire_6258, wire_6249, wire_6248, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_6327, wire_6326, wire_6317, wire_6316, wire_6307, wire_6306, wire_6263, wire_6262, wire_6253, wire_6252, wire_6243, wire_6242, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300, wire_6267, wire_6266, wire_6257, wire_6256, wire_6247, wire_6246, wire_6357, wire_6356, wire_6347, wire_6346, wire_6337, wire_6336, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_6325, wire_6324, wire_6315, wire_6314, wire_6305, wire_6304, wire_6261, wire_6260, wire_6251, wire_6250, wire_6241, wire_6240, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_6295, wire_6294, wire_6285, wire_6284, wire_6275, wire_6274};
    // FPGA IPIN IN
    assign io_tile_0_6_ipin_in = {wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_6325, wire_6324, wire_6315, wire_6314, wire_6305, wire_6304, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_6293, wire_6292, wire_6283, wire_6282, wire_6273, wire_6272, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_6297, wire_6296, wire_6287, wire_6286, wire_6277, wire_6276, wire_6357, wire_6356, wire_6347, wire_6346, wire_6337, wire_6336, wire_6291, wire_6290, wire_6281, wire_6280, wire_6271, wire_6270, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360, wire_6327, wire_6326, wire_6317, wire_6316, wire_6307, wire_6306, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_6295, wire_6294, wire_6285, wire_6284, wire_6275, wire_6274, wire_6385, wire_6384, wire_6375, wire_6374, wire_6365, wire_6364, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300};
    // FPGA IPIN IN
    assign io_tile_0_7_ipin_in = {wire_6415, wire_6414, wire_6405, wire_6404, wire_6395, wire_6394, wire_6359, wire_6358, wire_6349, wire_6348, wire_6339, wire_6338, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_6329, wire_6328, wire_6319, wire_6318, wire_6309, wire_6308, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_6387, wire_6386, wire_6377, wire_6376, wire_6367, wire_6366, wire_6323, wire_6322, wire_6313, wire_6312, wire_6303, wire_6302, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360, wire_6327, wire_6326, wire_6317, wire_6316, wire_6307, wire_6306, wire_6417, wire_6416, wire_6407, wire_6406, wire_6397, wire_6396, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_6385, wire_6384, wire_6375, wire_6374, wire_6365, wire_6364, wire_6321, wire_6320, wire_6311, wire_6310, wire_6301, wire_6300, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_6355, wire_6354, wire_6345, wire_6344, wire_6335, wire_6334};
    // FPGA IPIN IN
    assign io_tile_0_8_ipin_in = {wire_6449, wire_6448, wire_6439, wire_6438, wire_6429, wire_6428, wire_6385, wire_6384, wire_6375, wire_6374, wire_6365, wire_6364, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_6353, wire_6352, wire_6343, wire_6342, wire_6333, wire_6332, wire_6443, wire_6442, wire_6433, wire_6432, wire_6423, wire_6422, wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_6357, wire_6356, wire_6347, wire_6346, wire_6337, wire_6336, wire_6417, wire_6416, wire_6407, wire_6406, wire_6397, wire_6396, wire_6351, wire_6350, wire_6341, wire_6340, wire_6331, wire_6330, wire_6441, wire_6440, wire_6431, wire_6430, wire_6421, wire_6420, wire_6387, wire_6386, wire_6377, wire_6376, wire_6367, wire_6366, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_6355, wire_6354, wire_6345, wire_6344, wire_6335, wire_6334, wire_6445, wire_6444, wire_6435, wire_6434, wire_6425, wire_6424, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360};
    // FPGA IPIN IN
    assign io_tile_0_9_ipin_in = {wire_6475, wire_6474, wire_6465, wire_6464, wire_6455, wire_6454, wire_6419, wire_6418, wire_6409, wire_6408, wire_6399, wire_6398, wire_6443, wire_6442, wire_6433, wire_6432, wire_6423, wire_6422, wire_6389, wire_6388, wire_6379, wire_6378, wire_6369, wire_6368, wire_6479, wire_6478, wire_6469, wire_6468, wire_6459, wire_6458, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_6447, wire_6446, wire_6437, wire_6436, wire_6427, wire_6426, wire_6383, wire_6382, wire_6373, wire_6372, wire_6363, wire_6362, wire_6441, wire_6440, wire_6431, wire_6430, wire_6421, wire_6420, wire_6387, wire_6386, wire_6377, wire_6376, wire_6367, wire_6366, wire_6477, wire_6476, wire_6467, wire_6466, wire_6457, wire_6456, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_6445, wire_6444, wire_6435, wire_6434, wire_6425, wire_6424, wire_6381, wire_6380, wire_6371, wire_6370, wire_6361, wire_6360, wire_6471, wire_6470, wire_6461, wire_6460, wire_6451, wire_6450, wire_6415, wire_6414, wire_6405, wire_6404, wire_6395, wire_6394};
    // FPGA IPIN IN
    assign io_tile_0_10_ipin_in = {wire_6509, wire_6508, wire_6499, wire_6498, wire_6489, wire_6488, wire_6445, wire_6444, wire_6435, wire_6434, wire_6425, wire_6424, wire_6479, wire_6478, wire_6469, wire_6468, wire_6459, wire_6458, wire_6413, wire_6412, wire_6403, wire_6402, wire_6393, wire_6392, wire_6503, wire_6502, wire_6493, wire_6492, wire_6483, wire_6482, wire_6449, wire_6448, wire_6439, wire_6438, wire_6429, wire_6428, wire_6473, wire_6472, wire_6463, wire_6462, wire_6453, wire_6452, wire_6417, wire_6416, wire_6407, wire_6406, wire_6397, wire_6396, wire_6477, wire_6476, wire_6467, wire_6466, wire_6457, wire_6456, wire_6411, wire_6410, wire_6401, wire_6400, wire_6391, wire_6390, wire_6501, wire_6500, wire_6491, wire_6490, wire_6481, wire_6480, wire_6447, wire_6446, wire_6437, wire_6436, wire_6427, wire_6426, wire_6471, wire_6470, wire_6461, wire_6460, wire_6451, wire_6450, wire_6415, wire_6414, wire_6405, wire_6404, wire_6395, wire_6394, wire_6505, wire_6504, wire_6495, wire_6494, wire_6485, wire_6484, wire_6441, wire_6440, wire_6431, wire_6430, wire_6421, wire_6420};
    // FPGA IPIN IN
    assign io_tile_11_1_ipin_in = {wire_10135, wire_10134, wire_10123, wire_10122, wire_10095, wire_10094, wire_10083, wire_10082, wire_10055, wire_10054, wire_10043, wire_10042, wire_10133, wire_10132, wire_10121, wire_10120, wire_10093, wire_10092, wire_10081, wire_10080, wire_10053, wire_10052, wire_10041, wire_10040, wire_10137, wire_10136, wire_10109, wire_10108, wire_10097, wire_10096, wire_10069, wire_10068, wire_10057, wire_10056, wire_10029, wire_10028, wire_10127, wire_10126, wire_10115, wire_10114, wire_10087, wire_10086, wire_10075, wire_10074, wire_10047, wire_10046, wire_10035, wire_10034, wire_10125, wire_10124, wire_10113, wire_10112, wire_10085, wire_10084, wire_10073, wire_10072, wire_10045, wire_10044, wire_10033, wire_10032, wire_10131, wire_10130, wire_10103, wire_10102, wire_10091, wire_10090, wire_10063, wire_10062, wire_10051, wire_10050, wire_10023, wire_10022, wire_10119, wire_10118, wire_10107, wire_10106, wire_10079, wire_10078, wire_10067, wire_10066, wire_10039, wire_10038, wire_10027, wire_10026, wire_10117, wire_10116, wire_10105, wire_10104, wire_10077, wire_10076, wire_10065, wire_10064, wire_10037, wire_10036, wire_10025, wire_10024};
    // FPGA IPIN IN
    assign io_tile_11_2_ipin_in = {wire_10133, wire_10132, wire_10121, wire_10120, wire_10093, wire_10092, wire_10081, wire_10080, wire_10053, wire_10052, wire_10041, wire_10040, wire_10169, wire_10168, wire_10159, wire_10158, wire_10149, wire_10148, wire_10119, wire_10118, wire_10079, wire_10078, wire_10039, wire_10038, wire_10163, wire_10162, wire_10153, wire_10152, wire_10143, wire_10142, wire_10135, wire_10134, wire_10095, wire_10094, wire_10055, wire_10054, wire_10125, wire_10124, wire_10113, wire_10112, wire_10085, wire_10084, wire_10073, wire_10072, wire_10045, wire_10044, wire_10033, wire_10032, wire_10167, wire_10166, wire_10157, wire_10156, wire_10147, wire_10146, wire_10111, wire_10110, wire_10071, wire_10070, wire_10031, wire_10030, wire_10129, wire_10128, wire_10101, wire_10100, wire_10089, wire_10088, wire_10061, wire_10060, wire_10049, wire_10048, wire_10021, wire_10020, wire_10117, wire_10116, wire_10105, wire_10104, wire_10077, wire_10076, wire_10065, wire_10064, wire_10037, wire_10036, wire_10025, wire_10024, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10103, wire_10102, wire_10063, wire_10062, wire_10023, wire_10022};
    // FPGA IPIN IN
    assign io_tile_11_3_ipin_in = {wire_10169, wire_10168, wire_10159, wire_10158, wire_10149, wire_10148, wire_10119, wire_10118, wire_10079, wire_10078, wire_10039, wire_10038, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174, wire_10137, wire_10136, wire_10097, wire_10096, wire_10057, wire_10056, wire_10199, wire_10198, wire_10189, wire_10188, wire_10179, wire_10178, wire_10113, wire_10112, wire_10073, wire_10072, wire_10033, wire_10032, wire_10167, wire_10166, wire_10157, wire_10156, wire_10147, wire_10146, wire_10111, wire_10110, wire_10071, wire_10070, wire_10031, wire_10030, wire_10193, wire_10192, wire_10183, wire_10182, wire_10173, wire_10172, wire_10129, wire_10128, wire_10089, wire_10088, wire_10049, wire_10048, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140, wire_10127, wire_10126, wire_10087, wire_10086, wire_10047, wire_10046, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10103, wire_10102, wire_10063, wire_10062, wire_10023, wire_10022, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_10121, wire_10120, wire_10081, wire_10080, wire_10041, wire_10040};
    // FPGA IPIN IN
    assign io_tile_11_4_ipin_in = {wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174, wire_10137, wire_10136, wire_10097, wire_10096, wire_10057, wire_10056, wire_10229, wire_10228, wire_10219, wire_10218, wire_10209, wire_10208, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10223, wire_10222, wire_10213, wire_10212, wire_10203, wire_10202, wire_10169, wire_10168, wire_10159, wire_10158, wire_10149, wire_10148, wire_10193, wire_10192, wire_10183, wire_10182, wire_10173, wire_10172, wire_10129, wire_10128, wire_10089, wire_10088, wire_10049, wire_10048, wire_10227, wire_10226, wire_10217, wire_10216, wire_10207, wire_10206, wire_10163, wire_10162, wire_10153, wire_10152, wire_10143, wire_10142, wire_10197, wire_10196, wire_10187, wire_10186, wire_10177, wire_10176, wire_10105, wire_10104, wire_10065, wire_10064, wire_10025, wire_10024, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_10121, wire_10120, wire_10081, wire_10080, wire_10041, wire_10040, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140};
    // FPGA IPIN IN
    assign io_tile_11_5_ipin_in = {wire_10229, wire_10228, wire_10219, wire_10218, wire_10209, wire_10208, wire_10165, wire_10164, wire_10155, wire_10154, wire_10145, wire_10144, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234, wire_10199, wire_10198, wire_10189, wire_10188, wire_10179, wire_10178, wire_10259, wire_10258, wire_10249, wire_10248, wire_10239, wire_10238, wire_10193, wire_10192, wire_10183, wire_10182, wire_10173, wire_10172, wire_10227, wire_10226, wire_10217, wire_10216, wire_10207, wire_10206, wire_10163, wire_10162, wire_10153, wire_10152, wire_10143, wire_10142, wire_10253, wire_10252, wire_10243, wire_10242, wire_10233, wire_10232, wire_10197, wire_10196, wire_10187, wire_10186, wire_10177, wire_10176, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200, wire_10167, wire_10166, wire_10157, wire_10156, wire_10147, wire_10146, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10161, wire_10160, wire_10151, wire_10150, wire_10141, wire_10140, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174};
    // FPGA IPIN IN
    assign io_tile_11_6_ipin_in = {wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234, wire_10199, wire_10198, wire_10189, wire_10188, wire_10179, wire_10178, wire_10289, wire_10288, wire_10279, wire_10278, wire_10269, wire_10268, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10283, wire_10282, wire_10273, wire_10272, wire_10263, wire_10262, wire_10229, wire_10228, wire_10219, wire_10218, wire_10209, wire_10208, wire_10253, wire_10252, wire_10243, wire_10242, wire_10233, wire_10232, wire_10197, wire_10196, wire_10187, wire_10186, wire_10177, wire_10176, wire_10287, wire_10286, wire_10277, wire_10276, wire_10267, wire_10266, wire_10223, wire_10222, wire_10213, wire_10212, wire_10203, wire_10202, wire_10257, wire_10256, wire_10247, wire_10246, wire_10237, wire_10236, wire_10191, wire_10190, wire_10181, wire_10180, wire_10171, wire_10170, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_10195, wire_10194, wire_10185, wire_10184, wire_10175, wire_10174, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200};
    // FPGA IPIN IN
    assign io_tile_11_7_ipin_in = {wire_10289, wire_10288, wire_10279, wire_10278, wire_10269, wire_10268, wire_10225, wire_10224, wire_10215, wire_10214, wire_10205, wire_10204, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294, wire_10259, wire_10258, wire_10249, wire_10248, wire_10239, wire_10238, wire_10319, wire_10318, wire_10309, wire_10308, wire_10299, wire_10298, wire_10253, wire_10252, wire_10243, wire_10242, wire_10233, wire_10232, wire_10287, wire_10286, wire_10277, wire_10276, wire_10267, wire_10266, wire_10223, wire_10222, wire_10213, wire_10212, wire_10203, wire_10202, wire_10313, wire_10312, wire_10303, wire_10302, wire_10293, wire_10292, wire_10257, wire_10256, wire_10247, wire_10246, wire_10237, wire_10236, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260, wire_10227, wire_10226, wire_10217, wire_10216, wire_10207, wire_10206, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10221, wire_10220, wire_10211, wire_10210, wire_10201, wire_10200, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234};
    // FPGA IPIN IN
    assign io_tile_11_8_ipin_in = {wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294, wire_10259, wire_10258, wire_10249, wire_10248, wire_10239, wire_10238, wire_10349, wire_10348, wire_10339, wire_10338, wire_10329, wire_10328, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10343, wire_10342, wire_10333, wire_10332, wire_10323, wire_10322, wire_10289, wire_10288, wire_10279, wire_10278, wire_10269, wire_10268, wire_10313, wire_10312, wire_10303, wire_10302, wire_10293, wire_10292, wire_10257, wire_10256, wire_10247, wire_10246, wire_10237, wire_10236, wire_10347, wire_10346, wire_10337, wire_10336, wire_10327, wire_10326, wire_10283, wire_10282, wire_10273, wire_10272, wire_10263, wire_10262, wire_10317, wire_10316, wire_10307, wire_10306, wire_10297, wire_10296, wire_10251, wire_10250, wire_10241, wire_10240, wire_10231, wire_10230, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_10255, wire_10254, wire_10245, wire_10244, wire_10235, wire_10234, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260};
    // FPGA IPIN IN
    assign io_tile_11_9_ipin_in = {wire_10349, wire_10348, wire_10339, wire_10338, wire_10329, wire_10328, wire_10285, wire_10284, wire_10275, wire_10274, wire_10265, wire_10264, wire_10375, wire_10374, wire_10365, wire_10364, wire_10355, wire_10354, wire_10319, wire_10318, wire_10309, wire_10308, wire_10299, wire_10298, wire_10379, wire_10378, wire_10369, wire_10368, wire_10359, wire_10358, wire_10313, wire_10312, wire_10303, wire_10302, wire_10293, wire_10292, wire_10347, wire_10346, wire_10337, wire_10336, wire_10327, wire_10326, wire_10283, wire_10282, wire_10273, wire_10272, wire_10263, wire_10262, wire_10373, wire_10372, wire_10363, wire_10362, wire_10353, wire_10352, wire_10317, wire_10316, wire_10307, wire_10306, wire_10297, wire_10296, wire_10341, wire_10340, wire_10331, wire_10330, wire_10321, wire_10320, wire_10287, wire_10286, wire_10277, wire_10276, wire_10267, wire_10266, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_10281, wire_10280, wire_10271, wire_10270, wire_10261, wire_10260, wire_10371, wire_10370, wire_10361, wire_10360, wire_10351, wire_10350, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294};
    // FPGA IPIN IN
    assign io_tile_11_10_ipin_in = {wire_10375, wire_10374, wire_10365, wire_10364, wire_10355, wire_10354, wire_10319, wire_10318, wire_10309, wire_10308, wire_10299, wire_10298, wire_10409, wire_10408, wire_10399, wire_10398, wire_10389, wire_10388, wire_10345, wire_10344, wire_10335, wire_10334, wire_10325, wire_10324, wire_10403, wire_10402, wire_10393, wire_10392, wire_10383, wire_10382, wire_10349, wire_10348, wire_10339, wire_10338, wire_10329, wire_10328, wire_10373, wire_10372, wire_10363, wire_10362, wire_10353, wire_10352, wire_10317, wire_10316, wire_10307, wire_10306, wire_10297, wire_10296, wire_10407, wire_10406, wire_10397, wire_10396, wire_10387, wire_10386, wire_10343, wire_10342, wire_10333, wire_10332, wire_10323, wire_10322, wire_10377, wire_10376, wire_10367, wire_10366, wire_10357, wire_10356, wire_10311, wire_10310, wire_10301, wire_10300, wire_10291, wire_10290, wire_10371, wire_10370, wire_10361, wire_10360, wire_10351, wire_10350, wire_10315, wire_10314, wire_10305, wire_10304, wire_10295, wire_10294, wire_10405, wire_10404, wire_10395, wire_10394, wire_10385, wire_10384, wire_10341, wire_10340, wire_10331, wire_10330, wire_10321, wire_10320};
    // FPGA IPIN IN


    // FPGA IO OPIN
    assign wire_25 = io_tile_1_0_opin_out[0];
    assign wire_28 = io_tile_1_0_opin_out[1];
    assign wire_31 = io_tile_1_0_opin_out[2];
    assign wire_34 = io_tile_1_0_opin_out[3];
    assign wire_37 = io_tile_1_0_opin_out[4];
    assign wire_40 = io_tile_1_0_opin_out[5];
    assign wire_43 = io_tile_1_0_opin_out[6];
    assign wire_46 = io_tile_1_0_opin_out[7];
    assign wire_73 = io_tile_2_0_opin_out[0];
    assign wire_76 = io_tile_2_0_opin_out[1];
    assign wire_79 = io_tile_2_0_opin_out[2];
    assign wire_82 = io_tile_2_0_opin_out[3];
    assign wire_85 = io_tile_2_0_opin_out[4];
    assign wire_88 = io_tile_2_0_opin_out[5];
    assign wire_91 = io_tile_2_0_opin_out[6];
    assign wire_94 = io_tile_2_0_opin_out[7];
    assign wire_121 = io_tile_3_0_opin_out[0];
    assign wire_124 = io_tile_3_0_opin_out[1];
    assign wire_127 = io_tile_3_0_opin_out[2];
    assign wire_130 = io_tile_3_0_opin_out[3];
    assign wire_133 = io_tile_3_0_opin_out[4];
    assign wire_136 = io_tile_3_0_opin_out[5];
    assign wire_139 = io_tile_3_0_opin_out[6];
    assign wire_142 = io_tile_3_0_opin_out[7];
    assign wire_169 = io_tile_4_0_opin_out[0];
    assign wire_172 = io_tile_4_0_opin_out[1];
    assign wire_175 = io_tile_4_0_opin_out[2];
    assign wire_178 = io_tile_4_0_opin_out[3];
    assign wire_181 = io_tile_4_0_opin_out[4];
    assign wire_184 = io_tile_4_0_opin_out[5];
    assign wire_187 = io_tile_4_0_opin_out[6];
    assign wire_190 = io_tile_4_0_opin_out[7];
    assign wire_217 = io_tile_5_0_opin_out[0];
    assign wire_220 = io_tile_5_0_opin_out[1];
    assign wire_223 = io_tile_5_0_opin_out[2];
    assign wire_226 = io_tile_5_0_opin_out[3];
    assign wire_229 = io_tile_5_0_opin_out[4];
    assign wire_232 = io_tile_5_0_opin_out[5];
    assign wire_235 = io_tile_5_0_opin_out[6];
    assign wire_238 = io_tile_5_0_opin_out[7];
    assign wire_265 = io_tile_6_0_opin_out[0];
    assign wire_268 = io_tile_6_0_opin_out[1];
    assign wire_271 = io_tile_6_0_opin_out[2];
    assign wire_274 = io_tile_6_0_opin_out[3];
    assign wire_277 = io_tile_6_0_opin_out[4];
    assign wire_280 = io_tile_6_0_opin_out[5];
    assign wire_283 = io_tile_6_0_opin_out[6];
    assign wire_286 = io_tile_6_0_opin_out[7];
    assign wire_313 = io_tile_7_0_opin_out[0];
    assign wire_316 = io_tile_7_0_opin_out[1];
    assign wire_319 = io_tile_7_0_opin_out[2];
    assign wire_322 = io_tile_7_0_opin_out[3];
    assign wire_325 = io_tile_7_0_opin_out[4];
    assign wire_328 = io_tile_7_0_opin_out[5];
    assign wire_331 = io_tile_7_0_opin_out[6];
    assign wire_334 = io_tile_7_0_opin_out[7];
    assign wire_361 = io_tile_8_0_opin_out[0];
    assign wire_364 = io_tile_8_0_opin_out[1];
    assign wire_367 = io_tile_8_0_opin_out[2];
    assign wire_370 = io_tile_8_0_opin_out[3];
    assign wire_373 = io_tile_8_0_opin_out[4];
    assign wire_376 = io_tile_8_0_opin_out[5];
    assign wire_379 = io_tile_8_0_opin_out[6];
    assign wire_382 = io_tile_8_0_opin_out[7];
    assign wire_409 = io_tile_9_0_opin_out[0];
    assign wire_412 = io_tile_9_0_opin_out[1];
    assign wire_415 = io_tile_9_0_opin_out[2];
    assign wire_418 = io_tile_9_0_opin_out[3];
    assign wire_421 = io_tile_9_0_opin_out[4];
    assign wire_424 = io_tile_9_0_opin_out[5];
    assign wire_427 = io_tile_9_0_opin_out[6];
    assign wire_430 = io_tile_9_0_opin_out[7];
    assign wire_457 = io_tile_10_0_opin_out[0];
    assign wire_460 = io_tile_10_0_opin_out[1];
    assign wire_463 = io_tile_10_0_opin_out[2];
    assign wire_466 = io_tile_10_0_opin_out[3];
    assign wire_469 = io_tile_10_0_opin_out[4];
    assign wire_472 = io_tile_10_0_opin_out[5];
    assign wire_475 = io_tile_10_0_opin_out[6];
    assign wire_478 = io_tile_10_0_opin_out[7];
    assign wire_5665 = io_tile_1_11_opin_out[0];
    assign wire_5668 = io_tile_1_11_opin_out[1];
    assign wire_5671 = io_tile_1_11_opin_out[2];
    assign wire_5674 = io_tile_1_11_opin_out[3];
    assign wire_5677 = io_tile_1_11_opin_out[4];
    assign wire_5680 = io_tile_1_11_opin_out[5];
    assign wire_5683 = io_tile_1_11_opin_out[6];
    assign wire_5686 = io_tile_1_11_opin_out[7];
    assign wire_5713 = io_tile_2_11_opin_out[0];
    assign wire_5716 = io_tile_2_11_opin_out[1];
    assign wire_5719 = io_tile_2_11_opin_out[2];
    assign wire_5722 = io_tile_2_11_opin_out[3];
    assign wire_5725 = io_tile_2_11_opin_out[4];
    assign wire_5728 = io_tile_2_11_opin_out[5];
    assign wire_5731 = io_tile_2_11_opin_out[6];
    assign wire_5734 = io_tile_2_11_opin_out[7];
    assign wire_5761 = io_tile_3_11_opin_out[0];
    assign wire_5764 = io_tile_3_11_opin_out[1];
    assign wire_5767 = io_tile_3_11_opin_out[2];
    assign wire_5770 = io_tile_3_11_opin_out[3];
    assign wire_5773 = io_tile_3_11_opin_out[4];
    assign wire_5776 = io_tile_3_11_opin_out[5];
    assign wire_5779 = io_tile_3_11_opin_out[6];
    assign wire_5782 = io_tile_3_11_opin_out[7];
    assign wire_5809 = io_tile_4_11_opin_out[0];
    assign wire_5812 = io_tile_4_11_opin_out[1];
    assign wire_5815 = io_tile_4_11_opin_out[2];
    assign wire_5818 = io_tile_4_11_opin_out[3];
    assign wire_5821 = io_tile_4_11_opin_out[4];
    assign wire_5824 = io_tile_4_11_opin_out[5];
    assign wire_5827 = io_tile_4_11_opin_out[6];
    assign wire_5830 = io_tile_4_11_opin_out[7];
    assign wire_5857 = io_tile_5_11_opin_out[0];
    assign wire_5860 = io_tile_5_11_opin_out[1];
    assign wire_5863 = io_tile_5_11_opin_out[2];
    assign wire_5866 = io_tile_5_11_opin_out[3];
    assign wire_5869 = io_tile_5_11_opin_out[4];
    assign wire_5872 = io_tile_5_11_opin_out[5];
    assign wire_5875 = io_tile_5_11_opin_out[6];
    assign wire_5878 = io_tile_5_11_opin_out[7];
    assign wire_5905 = io_tile_6_11_opin_out[0];
    assign wire_5908 = io_tile_6_11_opin_out[1];
    assign wire_5911 = io_tile_6_11_opin_out[2];
    assign wire_5914 = io_tile_6_11_opin_out[3];
    assign wire_5917 = io_tile_6_11_opin_out[4];
    assign wire_5920 = io_tile_6_11_opin_out[5];
    assign wire_5923 = io_tile_6_11_opin_out[6];
    assign wire_5926 = io_tile_6_11_opin_out[7];
    assign wire_5953 = io_tile_7_11_opin_out[0];
    assign wire_5956 = io_tile_7_11_opin_out[1];
    assign wire_5959 = io_tile_7_11_opin_out[2];
    assign wire_5962 = io_tile_7_11_opin_out[3];
    assign wire_5965 = io_tile_7_11_opin_out[4];
    assign wire_5968 = io_tile_7_11_opin_out[5];
    assign wire_5971 = io_tile_7_11_opin_out[6];
    assign wire_5974 = io_tile_7_11_opin_out[7];
    assign wire_6001 = io_tile_8_11_opin_out[0];
    assign wire_6004 = io_tile_8_11_opin_out[1];
    assign wire_6007 = io_tile_8_11_opin_out[2];
    assign wire_6010 = io_tile_8_11_opin_out[3];
    assign wire_6013 = io_tile_8_11_opin_out[4];
    assign wire_6016 = io_tile_8_11_opin_out[5];
    assign wire_6019 = io_tile_8_11_opin_out[6];
    assign wire_6022 = io_tile_8_11_opin_out[7];
    assign wire_6049 = io_tile_9_11_opin_out[0];
    assign wire_6052 = io_tile_9_11_opin_out[1];
    assign wire_6055 = io_tile_9_11_opin_out[2];
    assign wire_6058 = io_tile_9_11_opin_out[3];
    assign wire_6061 = io_tile_9_11_opin_out[4];
    assign wire_6064 = io_tile_9_11_opin_out[5];
    assign wire_6067 = io_tile_9_11_opin_out[6];
    assign wire_6070 = io_tile_9_11_opin_out[7];
    assign wire_6097 = io_tile_10_11_opin_out[0];
    assign wire_6100 = io_tile_10_11_opin_out[1];
    assign wire_6103 = io_tile_10_11_opin_out[2];
    assign wire_6106 = io_tile_10_11_opin_out[3];
    assign wire_6109 = io_tile_10_11_opin_out[4];
    assign wire_6112 = io_tile_10_11_opin_out[5];
    assign wire_6115 = io_tile_10_11_opin_out[6];
    assign wire_6118 = io_tile_10_11_opin_out[7];
    assign wire_505 = io_tile_0_1_opin_out[0];
    assign wire_508 = io_tile_0_1_opin_out[1];
    assign wire_511 = io_tile_0_1_opin_out[2];
    assign wire_514 = io_tile_0_1_opin_out[3];
    assign wire_517 = io_tile_0_1_opin_out[4];
    assign wire_520 = io_tile_0_1_opin_out[5];
    assign wire_523 = io_tile_0_1_opin_out[6];
    assign wire_526 = io_tile_0_1_opin_out[7];
    assign wire_1021 = io_tile_0_2_opin_out[0];
    assign wire_1024 = io_tile_0_2_opin_out[1];
    assign wire_1027 = io_tile_0_2_opin_out[2];
    assign wire_1030 = io_tile_0_2_opin_out[3];
    assign wire_1033 = io_tile_0_2_opin_out[4];
    assign wire_1036 = io_tile_0_2_opin_out[5];
    assign wire_1039 = io_tile_0_2_opin_out[6];
    assign wire_1042 = io_tile_0_2_opin_out[7];
    assign wire_1537 = io_tile_0_3_opin_out[0];
    assign wire_1540 = io_tile_0_3_opin_out[1];
    assign wire_1543 = io_tile_0_3_opin_out[2];
    assign wire_1546 = io_tile_0_3_opin_out[3];
    assign wire_1549 = io_tile_0_3_opin_out[4];
    assign wire_1552 = io_tile_0_3_opin_out[5];
    assign wire_1555 = io_tile_0_3_opin_out[6];
    assign wire_1558 = io_tile_0_3_opin_out[7];
    assign wire_2053 = io_tile_0_4_opin_out[0];
    assign wire_2056 = io_tile_0_4_opin_out[1];
    assign wire_2059 = io_tile_0_4_opin_out[2];
    assign wire_2062 = io_tile_0_4_opin_out[3];
    assign wire_2065 = io_tile_0_4_opin_out[4];
    assign wire_2068 = io_tile_0_4_opin_out[5];
    assign wire_2071 = io_tile_0_4_opin_out[6];
    assign wire_2074 = io_tile_0_4_opin_out[7];
    assign wire_2569 = io_tile_0_5_opin_out[0];
    assign wire_2572 = io_tile_0_5_opin_out[1];
    assign wire_2575 = io_tile_0_5_opin_out[2];
    assign wire_2578 = io_tile_0_5_opin_out[3];
    assign wire_2581 = io_tile_0_5_opin_out[4];
    assign wire_2584 = io_tile_0_5_opin_out[5];
    assign wire_2587 = io_tile_0_5_opin_out[6];
    assign wire_2590 = io_tile_0_5_opin_out[7];
    assign wire_3085 = io_tile_0_6_opin_out[0];
    assign wire_3088 = io_tile_0_6_opin_out[1];
    assign wire_3091 = io_tile_0_6_opin_out[2];
    assign wire_3094 = io_tile_0_6_opin_out[3];
    assign wire_3097 = io_tile_0_6_opin_out[4];
    assign wire_3100 = io_tile_0_6_opin_out[5];
    assign wire_3103 = io_tile_0_6_opin_out[6];
    assign wire_3106 = io_tile_0_6_opin_out[7];
    assign wire_3601 = io_tile_0_7_opin_out[0];
    assign wire_3604 = io_tile_0_7_opin_out[1];
    assign wire_3607 = io_tile_0_7_opin_out[2];
    assign wire_3610 = io_tile_0_7_opin_out[3];
    assign wire_3613 = io_tile_0_7_opin_out[4];
    assign wire_3616 = io_tile_0_7_opin_out[5];
    assign wire_3619 = io_tile_0_7_opin_out[6];
    assign wire_3622 = io_tile_0_7_opin_out[7];
    assign wire_4117 = io_tile_0_8_opin_out[0];
    assign wire_4120 = io_tile_0_8_opin_out[1];
    assign wire_4123 = io_tile_0_8_opin_out[2];
    assign wire_4126 = io_tile_0_8_opin_out[3];
    assign wire_4129 = io_tile_0_8_opin_out[4];
    assign wire_4132 = io_tile_0_8_opin_out[5];
    assign wire_4135 = io_tile_0_8_opin_out[6];
    assign wire_4138 = io_tile_0_8_opin_out[7];
    assign wire_4633 = io_tile_0_9_opin_out[0];
    assign wire_4636 = io_tile_0_9_opin_out[1];
    assign wire_4639 = io_tile_0_9_opin_out[2];
    assign wire_4642 = io_tile_0_9_opin_out[3];
    assign wire_4645 = io_tile_0_9_opin_out[4];
    assign wire_4648 = io_tile_0_9_opin_out[5];
    assign wire_4651 = io_tile_0_9_opin_out[6];
    assign wire_4654 = io_tile_0_9_opin_out[7];
    assign wire_5149 = io_tile_0_10_opin_out[0];
    assign wire_5152 = io_tile_0_10_opin_out[1];
    assign wire_5155 = io_tile_0_10_opin_out[2];
    assign wire_5158 = io_tile_0_10_opin_out[3];
    assign wire_5161 = io_tile_0_10_opin_out[4];
    assign wire_5164 = io_tile_0_10_opin_out[5];
    assign wire_5167 = io_tile_0_10_opin_out[6];
    assign wire_5170 = io_tile_0_10_opin_out[7];
    assign wire_973 = io_tile_11_1_opin_out[0];
    assign wire_976 = io_tile_11_1_opin_out[1];
    assign wire_979 = io_tile_11_1_opin_out[2];
    assign wire_982 = io_tile_11_1_opin_out[3];
    assign wire_985 = io_tile_11_1_opin_out[4];
    assign wire_988 = io_tile_11_1_opin_out[5];
    assign wire_991 = io_tile_11_1_opin_out[6];
    assign wire_994 = io_tile_11_1_opin_out[7];
    assign wire_1489 = io_tile_11_2_opin_out[0];
    assign wire_1492 = io_tile_11_2_opin_out[1];
    assign wire_1495 = io_tile_11_2_opin_out[2];
    assign wire_1498 = io_tile_11_2_opin_out[3];
    assign wire_1501 = io_tile_11_2_opin_out[4];
    assign wire_1504 = io_tile_11_2_opin_out[5];
    assign wire_1507 = io_tile_11_2_opin_out[6];
    assign wire_1510 = io_tile_11_2_opin_out[7];
    assign wire_2005 = io_tile_11_3_opin_out[0];
    assign wire_2008 = io_tile_11_3_opin_out[1];
    assign wire_2011 = io_tile_11_3_opin_out[2];
    assign wire_2014 = io_tile_11_3_opin_out[3];
    assign wire_2017 = io_tile_11_3_opin_out[4];
    assign wire_2020 = io_tile_11_3_opin_out[5];
    assign wire_2023 = io_tile_11_3_opin_out[6];
    assign wire_2026 = io_tile_11_3_opin_out[7];
    assign wire_2521 = io_tile_11_4_opin_out[0];
    assign wire_2524 = io_tile_11_4_opin_out[1];
    assign wire_2527 = io_tile_11_4_opin_out[2];
    assign wire_2530 = io_tile_11_4_opin_out[3];
    assign wire_2533 = io_tile_11_4_opin_out[4];
    assign wire_2536 = io_tile_11_4_opin_out[5];
    assign wire_2539 = io_tile_11_4_opin_out[6];
    assign wire_2542 = io_tile_11_4_opin_out[7];
    assign wire_3037 = io_tile_11_5_opin_out[0];
    assign wire_3040 = io_tile_11_5_opin_out[1];
    assign wire_3043 = io_tile_11_5_opin_out[2];
    assign wire_3046 = io_tile_11_5_opin_out[3];
    assign wire_3049 = io_tile_11_5_opin_out[4];
    assign wire_3052 = io_tile_11_5_opin_out[5];
    assign wire_3055 = io_tile_11_5_opin_out[6];
    assign wire_3058 = io_tile_11_5_opin_out[7];
    assign wire_3553 = io_tile_11_6_opin_out[0];
    assign wire_3556 = io_tile_11_6_opin_out[1];
    assign wire_3559 = io_tile_11_6_opin_out[2];
    assign wire_3562 = io_tile_11_6_opin_out[3];
    assign wire_3565 = io_tile_11_6_opin_out[4];
    assign wire_3568 = io_tile_11_6_opin_out[5];
    assign wire_3571 = io_tile_11_6_opin_out[6];
    assign wire_3574 = io_tile_11_6_opin_out[7];
    assign wire_4069 = io_tile_11_7_opin_out[0];
    assign wire_4072 = io_tile_11_7_opin_out[1];
    assign wire_4075 = io_tile_11_7_opin_out[2];
    assign wire_4078 = io_tile_11_7_opin_out[3];
    assign wire_4081 = io_tile_11_7_opin_out[4];
    assign wire_4084 = io_tile_11_7_opin_out[5];
    assign wire_4087 = io_tile_11_7_opin_out[6];
    assign wire_4090 = io_tile_11_7_opin_out[7];
    assign wire_4585 = io_tile_11_8_opin_out[0];
    assign wire_4588 = io_tile_11_8_opin_out[1];
    assign wire_4591 = io_tile_11_8_opin_out[2];
    assign wire_4594 = io_tile_11_8_opin_out[3];
    assign wire_4597 = io_tile_11_8_opin_out[4];
    assign wire_4600 = io_tile_11_8_opin_out[5];
    assign wire_4603 = io_tile_11_8_opin_out[6];
    assign wire_4606 = io_tile_11_8_opin_out[7];
    assign wire_5101 = io_tile_11_9_opin_out[0];
    assign wire_5104 = io_tile_11_9_opin_out[1];
    assign wire_5107 = io_tile_11_9_opin_out[2];
    assign wire_5110 = io_tile_11_9_opin_out[3];
    assign wire_5113 = io_tile_11_9_opin_out[4];
    assign wire_5116 = io_tile_11_9_opin_out[5];
    assign wire_5119 = io_tile_11_9_opin_out[6];
    assign wire_5122 = io_tile_11_9_opin_out[7];
    assign wire_5617 = io_tile_11_10_opin_out[0];
    assign wire_5620 = io_tile_11_10_opin_out[1];
    assign wire_5623 = io_tile_11_10_opin_out[2];
    assign wire_5626 = io_tile_11_10_opin_out[3];
    assign wire_5629 = io_tile_11_10_opin_out[4];
    assign wire_5632 = io_tile_11_10_opin_out[5];
    assign wire_5635 = io_tile_11_10_opin_out[6];
    assign wire_5638 = io_tile_11_10_opin_out[7];
    // FPGA IO CHANXY
    assign io_tile_1_0_chanxy_in = {wire_6121, wire_565, wire_6239, wire_565, wire_10559, wire_6629, wire_6599, wire_6569, wire_6539, wire_565, wire_46, wire_37, wire_31, wire_6237, wire_565, wire_6235, wire_565, wire_6233, wire_565, wire_6231, wire_565, wire_10557, wire_6627, wire_6597, wire_6567, wire_6537, wire_565, wire_46, wire_37, wire_31, wire_6229, wire_561, wire_6227, wire_561, wire_6225, wire_561, wire_6223, wire_561, wire_10555, wire_6625, wire_6595, wire_6565, wire_6535, wire_565, wire_46, wire_37, wire_31, wire_6221, wire_561, wire_6219, wire_561, wire_6217, wire_46, wire_6215, wire_46, wire_10553, wire_6623, wire_6593, wire_6563, wire_6533, wire_565, wire_43, wire_37, wire_28, wire_6213, wire_46, wire_6211, wire_46, wire_6209, wire_46, wire_6207, wire_46, wire_10551, wire_6621, wire_6591, wire_6561, wire_6531, wire_565, wire_43, wire_37, wire_28, wire_6205, wire_43, wire_6203, wire_43, wire_6201, wire_43, wire_6199, wire_43, wire_10549, wire_6619, wire_6589, wire_6559, wire_6529, wire_565, wire_43, wire_37, wire_28, wire_6197, wire_43, wire_6195, wire_43, wire_6193, wire_40, wire_6191, wire_40, wire_10547, wire_6617, wire_6587, wire_6557, wire_6527, wire_561, wire_43, wire_34, wire_28, wire_6189, wire_40, wire_6187, wire_40, wire_6185, wire_40, wire_6183, wire_40, wire_10545, wire_6615, wire_6585, wire_6555, wire_6525, wire_561, wire_43, wire_34, wire_28, wire_6181, wire_37, wire_6179, wire_37, wire_6177, wire_37, wire_6175, wire_37, wire_10543, wire_6613, wire_6583, wire_6553, wire_6523, wire_561, wire_43, wire_34, wire_28, wire_6173, wire_37, wire_6171, wire_37, wire_6169, wire_34, wire_6167, wire_34, wire_10541, wire_6611, wire_6581, wire_6551, wire_6521, wire_561, wire_40, wire_34, wire_25, wire_6165, wire_34, wire_6163, wire_34, wire_6161, wire_34, wire_6159, wire_34, wire_10539, wire_6609, wire_6579, wire_6549, wire_6519, wire_561, wire_40, wire_34, wire_25, wire_6157, wire_31, wire_6155, wire_31, wire_6153, wire_31, wire_6151, wire_31, wire_10537, wire_6607, wire_6577, wire_6547, wire_6517, wire_561, wire_40, wire_34, wire_25, wire_6149, wire_31, wire_6147, wire_31, wire_6145, wire_28, wire_6143, wire_28, wire_10535, wire_6605, wire_6575, wire_6545, wire_6515, wire_46, wire_40, wire_31, wire_25, wire_6141, wire_28, wire_6139, wire_28, wire_6137, wire_28, wire_6135, wire_28, wire_10533, wire_6603, wire_6573, wire_6543, wire_6513, wire_46, wire_40, wire_31, wire_25, wire_6133, wire_25, wire_6131, wire_25, wire_6129, wire_25, wire_6127, wire_25, wire_10531, wire_6601, wire_6571, wire_6541, wire_6511, wire_46, wire_40, wire_31, wire_25, wire_6125, wire_25, wire_6123, wire_25};
    // CHNAXY TOTAL: 75
    assign wire_10410 = io_tile_1_0_chanxy_out[0];
    assign wire_10412 = io_tile_1_0_chanxy_out[1];
    assign wire_10413 = io_tile_1_0_chanxy_out[2];
    assign wire_10414 = io_tile_1_0_chanxy_out[3];
    assign wire_10416 = io_tile_1_0_chanxy_out[4];
    assign wire_10418 = io_tile_1_0_chanxy_out[5];
    assign wire_10420 = io_tile_1_0_chanxy_out[6];
    assign wire_10421 = io_tile_1_0_chanxy_out[7];
    assign wire_10422 = io_tile_1_0_chanxy_out[8];
    assign wire_10424 = io_tile_1_0_chanxy_out[9];
    assign wire_10426 = io_tile_1_0_chanxy_out[10];
    assign wire_10428 = io_tile_1_0_chanxy_out[11];
    assign wire_10429 = io_tile_1_0_chanxy_out[12];
    assign wire_10430 = io_tile_1_0_chanxy_out[13];
    assign wire_10432 = io_tile_1_0_chanxy_out[14];
    assign wire_10434 = io_tile_1_0_chanxy_out[15];
    assign wire_10436 = io_tile_1_0_chanxy_out[16];
    assign wire_10437 = io_tile_1_0_chanxy_out[17];
    assign wire_10438 = io_tile_1_0_chanxy_out[18];
    assign wire_10440 = io_tile_1_0_chanxy_out[19];
    assign wire_10442 = io_tile_1_0_chanxy_out[20];
    assign wire_10444 = io_tile_1_0_chanxy_out[21];
    assign wire_10445 = io_tile_1_0_chanxy_out[22];
    assign wire_10446 = io_tile_1_0_chanxy_out[23];
    assign wire_10448 = io_tile_1_0_chanxy_out[24];
    assign wire_10450 = io_tile_1_0_chanxy_out[25];
    assign wire_10452 = io_tile_1_0_chanxy_out[26];
    assign wire_10453 = io_tile_1_0_chanxy_out[27];
    assign wire_10454 = io_tile_1_0_chanxy_out[28];
    assign wire_10456 = io_tile_1_0_chanxy_out[29];
    assign wire_10458 = io_tile_1_0_chanxy_out[30];
    assign wire_10460 = io_tile_1_0_chanxy_out[31];
    assign wire_10461 = io_tile_1_0_chanxy_out[32];
    assign wire_10462 = io_tile_1_0_chanxy_out[33];
    assign wire_10464 = io_tile_1_0_chanxy_out[34];
    assign wire_10466 = io_tile_1_0_chanxy_out[35];
    assign wire_10468 = io_tile_1_0_chanxy_out[36];
    assign wire_10469 = io_tile_1_0_chanxy_out[37];
    assign wire_10470 = io_tile_1_0_chanxy_out[38];
    assign wire_10472 = io_tile_1_0_chanxy_out[39];
    assign wire_10474 = io_tile_1_0_chanxy_out[40];
    assign wire_10476 = io_tile_1_0_chanxy_out[41];
    assign wire_10477 = io_tile_1_0_chanxy_out[42];
    assign wire_10478 = io_tile_1_0_chanxy_out[43];
    assign wire_10480 = io_tile_1_0_chanxy_out[44];
    assign wire_10482 = io_tile_1_0_chanxy_out[45];
    assign wire_10484 = io_tile_1_0_chanxy_out[46];
    assign wire_10485 = io_tile_1_0_chanxy_out[47];
    assign wire_10486 = io_tile_1_0_chanxy_out[48];
    assign wire_10488 = io_tile_1_0_chanxy_out[49];
    assign wire_10490 = io_tile_1_0_chanxy_out[50];
    assign wire_10492 = io_tile_1_0_chanxy_out[51];
    assign wire_10493 = io_tile_1_0_chanxy_out[52];
    assign wire_10494 = io_tile_1_0_chanxy_out[53];
    assign wire_10496 = io_tile_1_0_chanxy_out[54];
    assign wire_10498 = io_tile_1_0_chanxy_out[55];
    assign wire_10500 = io_tile_1_0_chanxy_out[56];
    assign wire_10501 = io_tile_1_0_chanxy_out[57];
    assign wire_10502 = io_tile_1_0_chanxy_out[58];
    assign wire_10504 = io_tile_1_0_chanxy_out[59];
    assign wire_10506 = io_tile_1_0_chanxy_out[60];
    assign wire_10508 = io_tile_1_0_chanxy_out[61];
    assign wire_10509 = io_tile_1_0_chanxy_out[62];
    assign wire_10510 = io_tile_1_0_chanxy_out[63];
    assign wire_10512 = io_tile_1_0_chanxy_out[64];
    assign wire_10514 = io_tile_1_0_chanxy_out[65];
    assign wire_10516 = io_tile_1_0_chanxy_out[66];
    assign wire_10517 = io_tile_1_0_chanxy_out[67];
    assign wire_10518 = io_tile_1_0_chanxy_out[68];
    assign wire_10520 = io_tile_1_0_chanxy_out[69];
    assign wire_10522 = io_tile_1_0_chanxy_out[70];
    assign wire_10524 = io_tile_1_0_chanxy_out[71];
    assign wire_10525 = io_tile_1_0_chanxy_out[72];
    assign wire_10526 = io_tile_1_0_chanxy_out[73];
    assign wire_10528 = io_tile_1_0_chanxy_out[74];
    assign io_tile_2_0_chanxy_in = {wire_10524, wire_6629, wire_6599, wire_6569, wire_6539, wire_607, wire_94, wire_85, wire_79, wire_10516, wire_6627, wire_6597, wire_6567, wire_6537, wire_607, wire_94, wire_85, wire_79, wire_10508, wire_6625, wire_6595, wire_6565, wire_6535, wire_607, wire_94, wire_85, wire_79, wire_10500, wire_6623, wire_6593, wire_6563, wire_6533, wire_607, wire_91, wire_85, wire_76, wire_10492, wire_6621, wire_6591, wire_6561, wire_6531, wire_607, wire_91, wire_85, wire_76, wire_10484, wire_6619, wire_6589, wire_6559, wire_6529, wire_607, wire_91, wire_85, wire_76, wire_10476, wire_6617, wire_6587, wire_6557, wire_6527, wire_603, wire_91, wire_82, wire_76, wire_10468, wire_6615, wire_6585, wire_6555, wire_6525, wire_603, wire_91, wire_82, wire_76, wire_10460, wire_6613, wire_6583, wire_6553, wire_6523, wire_603, wire_91, wire_82, wire_76, wire_10452, wire_6611, wire_6581, wire_6551, wire_6521, wire_603, wire_88, wire_82, wire_73, wire_10444, wire_6609, wire_6579, wire_6549, wire_6519, wire_603, wire_88, wire_82, wire_73, wire_10436, wire_6607, wire_6577, wire_6547, wire_6517, wire_603, wire_88, wire_82, wire_73, wire_10428, wire_6605, wire_6575, wire_6545, wire_6515, wire_94, wire_88, wire_79, wire_73, wire_10420, wire_6603, wire_6573, wire_6543, wire_6513, wire_94, wire_88, wire_79, wire_73, wire_10412, wire_6601, wire_6571, wire_6541, wire_6511, wire_94, wire_88, wire_79, wire_73, wire_10589, wire_7019, wire_6989, wire_6959, wire_6929, wire_607, wire_94, wire_85, wire_79, wire_10587, wire_7017, wire_6987, wire_6957, wire_6927, wire_607, wire_94, wire_85, wire_79, wire_10585, wire_7015, wire_6985, wire_6955, wire_6925, wire_607, wire_94, wire_85, wire_79, wire_10583, wire_7013, wire_6983, wire_6953, wire_6923, wire_607, wire_91, wire_85, wire_76, wire_10581, wire_7011, wire_6981, wire_6951, wire_6921, wire_607, wire_91, wire_85, wire_76, wire_10579, wire_7009, wire_6979, wire_6949, wire_6919, wire_607, wire_91, wire_85, wire_76, wire_10577, wire_7007, wire_6977, wire_6947, wire_6917, wire_603, wire_91, wire_82, wire_76, wire_10575, wire_7005, wire_6975, wire_6945, wire_6915, wire_603, wire_91, wire_82, wire_76, wire_10573, wire_7003, wire_6973, wire_6943, wire_6913, wire_603, wire_91, wire_82, wire_76, wire_10571, wire_7001, wire_6971, wire_6941, wire_6911, wire_603, wire_88, wire_82, wire_73, wire_10569, wire_6999, wire_6969, wire_6939, wire_6909, wire_603, wire_88, wire_82, wire_73, wire_10567, wire_6997, wire_6967, wire_6937, wire_6907, wire_603, wire_88, wire_82, wire_73, wire_10565, wire_6995, wire_6965, wire_6935, wire_6905, wire_94, wire_88, wire_79, wire_73, wire_10563, wire_6993, wire_6963, wire_6933, wire_6903, wire_94, wire_88, wire_79, wire_73, wire_10561, wire_6991, wire_6961, wire_6931, wire_6901, wire_94, wire_88, wire_79, wire_73};
    // CHNAXY TOTAL: 30
    assign wire_10415 = io_tile_2_0_chanxy_out[0];
    assign wire_10423 = io_tile_2_0_chanxy_out[1];
    assign wire_10431 = io_tile_2_0_chanxy_out[2];
    assign wire_10439 = io_tile_2_0_chanxy_out[3];
    assign wire_10447 = io_tile_2_0_chanxy_out[4];
    assign wire_10455 = io_tile_2_0_chanxy_out[5];
    assign wire_10463 = io_tile_2_0_chanxy_out[6];
    assign wire_10471 = io_tile_2_0_chanxy_out[7];
    assign wire_10479 = io_tile_2_0_chanxy_out[8];
    assign wire_10487 = io_tile_2_0_chanxy_out[9];
    assign wire_10495 = io_tile_2_0_chanxy_out[10];
    assign wire_10503 = io_tile_2_0_chanxy_out[11];
    assign wire_10511 = io_tile_2_0_chanxy_out[12];
    assign wire_10519 = io_tile_2_0_chanxy_out[13];
    assign wire_10527 = io_tile_2_0_chanxy_out[14];
    assign wire_10530 = io_tile_2_0_chanxy_out[15];
    assign wire_10532 = io_tile_2_0_chanxy_out[16];
    assign wire_10534 = io_tile_2_0_chanxy_out[17];
    assign wire_10536 = io_tile_2_0_chanxy_out[18];
    assign wire_10538 = io_tile_2_0_chanxy_out[19];
    assign wire_10540 = io_tile_2_0_chanxy_out[20];
    assign wire_10542 = io_tile_2_0_chanxy_out[21];
    assign wire_10544 = io_tile_2_0_chanxy_out[22];
    assign wire_10546 = io_tile_2_0_chanxy_out[23];
    assign wire_10548 = io_tile_2_0_chanxy_out[24];
    assign wire_10550 = io_tile_2_0_chanxy_out[25];
    assign wire_10552 = io_tile_2_0_chanxy_out[26];
    assign wire_10554 = io_tile_2_0_chanxy_out[27];
    assign wire_10556 = io_tile_2_0_chanxy_out[28];
    assign wire_10558 = io_tile_2_0_chanxy_out[29];
    assign io_tile_3_0_chanxy_in = {wire_10526, wire_7019, wire_6989, wire_6959, wire_6929, wire_649, wire_142, wire_133, wire_127, wire_10518, wire_7017, wire_6987, wire_6957, wire_6927, wire_649, wire_142, wire_133, wire_127, wire_10510, wire_7015, wire_6985, wire_6955, wire_6925, wire_649, wire_142, wire_133, wire_127, wire_10502, wire_7013, wire_6983, wire_6953, wire_6923, wire_649, wire_139, wire_133, wire_124, wire_10494, wire_7011, wire_6981, wire_6951, wire_6921, wire_649, wire_139, wire_133, wire_124, wire_10486, wire_7009, wire_6979, wire_6949, wire_6919, wire_649, wire_139, wire_133, wire_124, wire_10478, wire_7007, wire_6977, wire_6947, wire_6917, wire_645, wire_139, wire_130, wire_124, wire_10470, wire_7005, wire_6975, wire_6945, wire_6915, wire_645, wire_139, wire_130, wire_124, wire_10462, wire_7003, wire_6973, wire_6943, wire_6913, wire_645, wire_139, wire_130, wire_124, wire_10454, wire_7001, wire_6971, wire_6941, wire_6911, wire_645, wire_136, wire_130, wire_121, wire_10446, wire_6999, wire_6969, wire_6939, wire_6909, wire_645, wire_136, wire_130, wire_121, wire_10438, wire_6997, wire_6967, wire_6937, wire_6907, wire_645, wire_136, wire_130, wire_121, wire_10430, wire_6995, wire_6965, wire_6935, wire_6905, wire_142, wire_136, wire_127, wire_121, wire_10422, wire_6993, wire_6963, wire_6933, wire_6903, wire_142, wire_136, wire_127, wire_121, wire_10414, wire_6991, wire_6961, wire_6931, wire_6901, wire_142, wire_136, wire_127, wire_121, wire_10619, wire_7409, wire_7379, wire_7349, wire_7319, wire_649, wire_142, wire_133, wire_127, wire_10617, wire_7407, wire_7377, wire_7347, wire_7317, wire_649, wire_142, wire_133, wire_127, wire_10615, wire_7405, wire_7375, wire_7345, wire_7315, wire_649, wire_142, wire_133, wire_127, wire_10613, wire_7403, wire_7373, wire_7343, wire_7313, wire_649, wire_139, wire_133, wire_124, wire_10611, wire_7401, wire_7371, wire_7341, wire_7311, wire_649, wire_139, wire_133, wire_124, wire_10609, wire_7399, wire_7369, wire_7339, wire_7309, wire_649, wire_139, wire_133, wire_124, wire_10607, wire_7397, wire_7367, wire_7337, wire_7307, wire_645, wire_139, wire_130, wire_124, wire_10605, wire_7395, wire_7365, wire_7335, wire_7305, wire_645, wire_139, wire_130, wire_124, wire_10603, wire_7393, wire_7363, wire_7333, wire_7303, wire_645, wire_139, wire_130, wire_124, wire_10601, wire_7391, wire_7361, wire_7331, wire_7301, wire_645, wire_136, wire_130, wire_121, wire_10599, wire_7389, wire_7359, wire_7329, wire_7299, wire_645, wire_136, wire_130, wire_121, wire_10597, wire_7387, wire_7357, wire_7327, wire_7297, wire_645, wire_136, wire_130, wire_121, wire_10595, wire_7385, wire_7355, wire_7325, wire_7295, wire_142, wire_136, wire_127, wire_121, wire_10593, wire_7383, wire_7353, wire_7323, wire_7293, wire_142, wire_136, wire_127, wire_121, wire_10591, wire_7381, wire_7351, wire_7321, wire_7291, wire_142, wire_136, wire_127, wire_121};
    // CHNAXY TOTAL: 30
    assign wire_10417 = io_tile_3_0_chanxy_out[0];
    assign wire_10425 = io_tile_3_0_chanxy_out[1];
    assign wire_10433 = io_tile_3_0_chanxy_out[2];
    assign wire_10441 = io_tile_3_0_chanxy_out[3];
    assign wire_10449 = io_tile_3_0_chanxy_out[4];
    assign wire_10457 = io_tile_3_0_chanxy_out[5];
    assign wire_10465 = io_tile_3_0_chanxy_out[6];
    assign wire_10473 = io_tile_3_0_chanxy_out[7];
    assign wire_10481 = io_tile_3_0_chanxy_out[8];
    assign wire_10489 = io_tile_3_0_chanxy_out[9];
    assign wire_10497 = io_tile_3_0_chanxy_out[10];
    assign wire_10505 = io_tile_3_0_chanxy_out[11];
    assign wire_10513 = io_tile_3_0_chanxy_out[12];
    assign wire_10521 = io_tile_3_0_chanxy_out[13];
    assign wire_10529 = io_tile_3_0_chanxy_out[14];
    assign wire_10560 = io_tile_3_0_chanxy_out[15];
    assign wire_10562 = io_tile_3_0_chanxy_out[16];
    assign wire_10564 = io_tile_3_0_chanxy_out[17];
    assign wire_10566 = io_tile_3_0_chanxy_out[18];
    assign wire_10568 = io_tile_3_0_chanxy_out[19];
    assign wire_10570 = io_tile_3_0_chanxy_out[20];
    assign wire_10572 = io_tile_3_0_chanxy_out[21];
    assign wire_10574 = io_tile_3_0_chanxy_out[22];
    assign wire_10576 = io_tile_3_0_chanxy_out[23];
    assign wire_10578 = io_tile_3_0_chanxy_out[24];
    assign wire_10580 = io_tile_3_0_chanxy_out[25];
    assign wire_10582 = io_tile_3_0_chanxy_out[26];
    assign wire_10584 = io_tile_3_0_chanxy_out[27];
    assign wire_10586 = io_tile_3_0_chanxy_out[28];
    assign wire_10588 = io_tile_3_0_chanxy_out[29];
    assign io_tile_4_0_chanxy_in = {wire_10528, wire_7409, wire_7379, wire_7349, wire_7319, wire_691, wire_190, wire_181, wire_175, wire_10520, wire_7407, wire_7377, wire_7347, wire_7317, wire_691, wire_190, wire_181, wire_175, wire_10512, wire_7405, wire_7375, wire_7345, wire_7315, wire_691, wire_190, wire_181, wire_175, wire_10504, wire_7403, wire_7373, wire_7343, wire_7313, wire_691, wire_187, wire_181, wire_172, wire_10496, wire_7401, wire_7371, wire_7341, wire_7311, wire_691, wire_187, wire_181, wire_172, wire_10488, wire_7399, wire_7369, wire_7339, wire_7309, wire_691, wire_187, wire_181, wire_172, wire_10480, wire_7397, wire_7367, wire_7337, wire_7307, wire_687, wire_187, wire_178, wire_172, wire_10472, wire_7395, wire_7365, wire_7335, wire_7305, wire_687, wire_187, wire_178, wire_172, wire_10464, wire_7393, wire_7363, wire_7333, wire_7303, wire_687, wire_187, wire_178, wire_172, wire_10456, wire_7391, wire_7361, wire_7331, wire_7301, wire_687, wire_184, wire_178, wire_169, wire_10448, wire_7389, wire_7359, wire_7329, wire_7299, wire_687, wire_184, wire_178, wire_169, wire_10440, wire_7387, wire_7357, wire_7327, wire_7297, wire_687, wire_184, wire_178, wire_169, wire_10432, wire_7385, wire_7355, wire_7325, wire_7295, wire_190, wire_184, wire_175, wire_169, wire_10424, wire_7383, wire_7353, wire_7323, wire_7293, wire_190, wire_184, wire_175, wire_169, wire_10416, wire_7381, wire_7351, wire_7321, wire_7291, wire_190, wire_184, wire_175, wire_169, wire_10649, wire_7799, wire_7769, wire_7739, wire_7709, wire_691, wire_190, wire_181, wire_175, wire_10647, wire_7797, wire_7767, wire_7737, wire_7707, wire_691, wire_190, wire_181, wire_175, wire_10645, wire_7795, wire_7765, wire_7735, wire_7705, wire_691, wire_190, wire_181, wire_175, wire_10643, wire_7793, wire_7763, wire_7733, wire_7703, wire_691, wire_187, wire_181, wire_172, wire_10641, wire_7791, wire_7761, wire_7731, wire_7701, wire_691, wire_187, wire_181, wire_172, wire_10639, wire_7789, wire_7759, wire_7729, wire_7699, wire_691, wire_187, wire_181, wire_172, wire_10637, wire_7787, wire_7757, wire_7727, wire_7697, wire_687, wire_187, wire_178, wire_172, wire_10635, wire_7785, wire_7755, wire_7725, wire_7695, wire_687, wire_187, wire_178, wire_172, wire_10633, wire_7783, wire_7753, wire_7723, wire_7693, wire_687, wire_187, wire_178, wire_172, wire_10631, wire_7781, wire_7751, wire_7721, wire_7691, wire_687, wire_184, wire_178, wire_169, wire_10629, wire_7779, wire_7749, wire_7719, wire_7689, wire_687, wire_184, wire_178, wire_169, wire_10627, wire_7777, wire_7747, wire_7717, wire_7687, wire_687, wire_184, wire_178, wire_169, wire_10625, wire_7775, wire_7745, wire_7715, wire_7685, wire_190, wire_184, wire_175, wire_169, wire_10623, wire_7773, wire_7743, wire_7713, wire_7683, wire_190, wire_184, wire_175, wire_169, wire_10621, wire_7771, wire_7741, wire_7711, wire_7681, wire_190, wire_184, wire_175, wire_169};
    // CHNAXY TOTAL: 30
    assign wire_10411 = io_tile_4_0_chanxy_out[0];
    assign wire_10419 = io_tile_4_0_chanxy_out[1];
    assign wire_10427 = io_tile_4_0_chanxy_out[2];
    assign wire_10435 = io_tile_4_0_chanxy_out[3];
    assign wire_10443 = io_tile_4_0_chanxy_out[4];
    assign wire_10451 = io_tile_4_0_chanxy_out[5];
    assign wire_10459 = io_tile_4_0_chanxy_out[6];
    assign wire_10467 = io_tile_4_0_chanxy_out[7];
    assign wire_10475 = io_tile_4_0_chanxy_out[8];
    assign wire_10483 = io_tile_4_0_chanxy_out[9];
    assign wire_10491 = io_tile_4_0_chanxy_out[10];
    assign wire_10499 = io_tile_4_0_chanxy_out[11];
    assign wire_10507 = io_tile_4_0_chanxy_out[12];
    assign wire_10515 = io_tile_4_0_chanxy_out[13];
    assign wire_10523 = io_tile_4_0_chanxy_out[14];
    assign wire_10590 = io_tile_4_0_chanxy_out[15];
    assign wire_10592 = io_tile_4_0_chanxy_out[16];
    assign wire_10594 = io_tile_4_0_chanxy_out[17];
    assign wire_10596 = io_tile_4_0_chanxy_out[18];
    assign wire_10598 = io_tile_4_0_chanxy_out[19];
    assign wire_10600 = io_tile_4_0_chanxy_out[20];
    assign wire_10602 = io_tile_4_0_chanxy_out[21];
    assign wire_10604 = io_tile_4_0_chanxy_out[22];
    assign wire_10606 = io_tile_4_0_chanxy_out[23];
    assign wire_10608 = io_tile_4_0_chanxy_out[24];
    assign wire_10610 = io_tile_4_0_chanxy_out[25];
    assign wire_10612 = io_tile_4_0_chanxy_out[26];
    assign wire_10614 = io_tile_4_0_chanxy_out[27];
    assign wire_10616 = io_tile_4_0_chanxy_out[28];
    assign wire_10618 = io_tile_4_0_chanxy_out[29];
    assign io_tile_5_0_chanxy_in = {wire_10522, wire_7799, wire_7769, wire_7739, wire_7709, wire_733, wire_238, wire_229, wire_223, wire_10514, wire_7797, wire_7767, wire_7737, wire_7707, wire_733, wire_238, wire_229, wire_223, wire_10506, wire_7795, wire_7765, wire_7735, wire_7705, wire_733, wire_238, wire_229, wire_223, wire_10498, wire_7793, wire_7763, wire_7733, wire_7703, wire_733, wire_235, wire_229, wire_220, wire_10490, wire_7791, wire_7761, wire_7731, wire_7701, wire_733, wire_235, wire_229, wire_220, wire_10482, wire_7789, wire_7759, wire_7729, wire_7699, wire_733, wire_235, wire_229, wire_220, wire_10474, wire_7787, wire_7757, wire_7727, wire_7697, wire_729, wire_235, wire_226, wire_220, wire_10466, wire_7785, wire_7755, wire_7725, wire_7695, wire_729, wire_235, wire_226, wire_220, wire_10458, wire_7783, wire_7753, wire_7723, wire_7693, wire_729, wire_235, wire_226, wire_220, wire_10450, wire_7781, wire_7751, wire_7721, wire_7691, wire_729, wire_232, wire_226, wire_217, wire_10442, wire_7779, wire_7749, wire_7719, wire_7689, wire_729, wire_232, wire_226, wire_217, wire_10434, wire_7777, wire_7747, wire_7717, wire_7687, wire_729, wire_232, wire_226, wire_217, wire_10426, wire_7775, wire_7745, wire_7715, wire_7685, wire_238, wire_232, wire_223, wire_217, wire_10418, wire_7773, wire_7743, wire_7713, wire_7683, wire_238, wire_232, wire_223, wire_217, wire_10410, wire_7771, wire_7741, wire_7711, wire_7681, wire_238, wire_232, wire_223, wire_217, wire_10679, wire_8189, wire_8159, wire_8129, wire_8099, wire_733, wire_238, wire_229, wire_223, wire_10677, wire_8187, wire_8157, wire_8127, wire_8097, wire_733, wire_238, wire_229, wire_223, wire_10675, wire_8185, wire_8155, wire_8125, wire_8095, wire_733, wire_238, wire_229, wire_223, wire_10673, wire_8183, wire_8153, wire_8123, wire_8093, wire_733, wire_235, wire_229, wire_220, wire_10671, wire_8181, wire_8151, wire_8121, wire_8091, wire_733, wire_235, wire_229, wire_220, wire_10669, wire_8179, wire_8149, wire_8119, wire_8089, wire_733, wire_235, wire_229, wire_220, wire_10667, wire_8177, wire_8147, wire_8117, wire_8087, wire_729, wire_235, wire_226, wire_220, wire_10665, wire_8175, wire_8145, wire_8115, wire_8085, wire_729, wire_235, wire_226, wire_220, wire_10663, wire_8173, wire_8143, wire_8113, wire_8083, wire_729, wire_235, wire_226, wire_220, wire_10661, wire_8171, wire_8141, wire_8111, wire_8081, wire_729, wire_232, wire_226, wire_217, wire_10659, wire_8169, wire_8139, wire_8109, wire_8079, wire_729, wire_232, wire_226, wire_217, wire_10657, wire_8167, wire_8137, wire_8107, wire_8077, wire_729, wire_232, wire_226, wire_217, wire_10655, wire_8165, wire_8135, wire_8105, wire_8075, wire_238, wire_232, wire_223, wire_217, wire_10653, wire_8163, wire_8133, wire_8103, wire_8073, wire_238, wire_232, wire_223, wire_217, wire_10651, wire_8161, wire_8131, wire_8101, wire_8071, wire_238, wire_232, wire_223, wire_217};
    // CHNAXY TOTAL: 30
    assign wire_10531 = io_tile_5_0_chanxy_out[0];
    assign wire_10533 = io_tile_5_0_chanxy_out[1];
    assign wire_10535 = io_tile_5_0_chanxy_out[2];
    assign wire_10537 = io_tile_5_0_chanxy_out[3];
    assign wire_10539 = io_tile_5_0_chanxy_out[4];
    assign wire_10541 = io_tile_5_0_chanxy_out[5];
    assign wire_10543 = io_tile_5_0_chanxy_out[6];
    assign wire_10545 = io_tile_5_0_chanxy_out[7];
    assign wire_10547 = io_tile_5_0_chanxy_out[8];
    assign wire_10549 = io_tile_5_0_chanxy_out[9];
    assign wire_10551 = io_tile_5_0_chanxy_out[10];
    assign wire_10553 = io_tile_5_0_chanxy_out[11];
    assign wire_10555 = io_tile_5_0_chanxy_out[12];
    assign wire_10557 = io_tile_5_0_chanxy_out[13];
    assign wire_10559 = io_tile_5_0_chanxy_out[14];
    assign wire_10620 = io_tile_5_0_chanxy_out[15];
    assign wire_10622 = io_tile_5_0_chanxy_out[16];
    assign wire_10624 = io_tile_5_0_chanxy_out[17];
    assign wire_10626 = io_tile_5_0_chanxy_out[18];
    assign wire_10628 = io_tile_5_0_chanxy_out[19];
    assign wire_10630 = io_tile_5_0_chanxy_out[20];
    assign wire_10632 = io_tile_5_0_chanxy_out[21];
    assign wire_10634 = io_tile_5_0_chanxy_out[22];
    assign wire_10636 = io_tile_5_0_chanxy_out[23];
    assign wire_10638 = io_tile_5_0_chanxy_out[24];
    assign wire_10640 = io_tile_5_0_chanxy_out[25];
    assign wire_10642 = io_tile_5_0_chanxy_out[26];
    assign wire_10644 = io_tile_5_0_chanxy_out[27];
    assign wire_10646 = io_tile_5_0_chanxy_out[28];
    assign wire_10648 = io_tile_5_0_chanxy_out[29];
    assign io_tile_6_0_chanxy_in = {wire_10558, wire_8189, wire_8159, wire_8129, wire_8099, wire_775, wire_286, wire_277, wire_271, wire_10556, wire_8187, wire_8157, wire_8127, wire_8097, wire_775, wire_286, wire_277, wire_271, wire_10554, wire_8185, wire_8155, wire_8125, wire_8095, wire_775, wire_286, wire_277, wire_271, wire_10552, wire_8183, wire_8153, wire_8123, wire_8093, wire_775, wire_283, wire_277, wire_268, wire_10550, wire_8181, wire_8151, wire_8121, wire_8091, wire_775, wire_283, wire_277, wire_268, wire_10548, wire_8179, wire_8149, wire_8119, wire_8089, wire_775, wire_283, wire_277, wire_268, wire_10546, wire_8177, wire_8147, wire_8117, wire_8087, wire_771, wire_283, wire_274, wire_268, wire_10544, wire_8175, wire_8145, wire_8115, wire_8085, wire_771, wire_283, wire_274, wire_268, wire_10542, wire_8173, wire_8143, wire_8113, wire_8083, wire_771, wire_283, wire_274, wire_268, wire_10540, wire_8171, wire_8141, wire_8111, wire_8081, wire_771, wire_280, wire_274, wire_265, wire_10538, wire_8169, wire_8139, wire_8109, wire_8079, wire_771, wire_280, wire_274, wire_265, wire_10536, wire_8167, wire_8137, wire_8107, wire_8077, wire_771, wire_280, wire_274, wire_265, wire_10534, wire_8165, wire_8135, wire_8105, wire_8075, wire_286, wire_280, wire_271, wire_265, wire_10532, wire_8163, wire_8133, wire_8103, wire_8073, wire_286, wire_280, wire_271, wire_265, wire_10530, wire_8161, wire_8131, wire_8101, wire_8071, wire_286, wire_280, wire_271, wire_265, wire_10709, wire_8579, wire_8549, wire_8519, wire_8489, wire_775, wire_286, wire_277, wire_271, wire_10707, wire_8577, wire_8547, wire_8517, wire_8487, wire_775, wire_286, wire_277, wire_271, wire_10705, wire_8575, wire_8545, wire_8515, wire_8485, wire_775, wire_286, wire_277, wire_271, wire_10703, wire_8573, wire_8543, wire_8513, wire_8483, wire_775, wire_283, wire_277, wire_268, wire_10701, wire_8571, wire_8541, wire_8511, wire_8481, wire_775, wire_283, wire_277, wire_268, wire_10699, wire_8569, wire_8539, wire_8509, wire_8479, wire_775, wire_283, wire_277, wire_268, wire_10697, wire_8567, wire_8537, wire_8507, wire_8477, wire_771, wire_283, wire_274, wire_268, wire_10695, wire_8565, wire_8535, wire_8505, wire_8475, wire_771, wire_283, wire_274, wire_268, wire_10693, wire_8563, wire_8533, wire_8503, wire_8473, wire_771, wire_283, wire_274, wire_268, wire_10691, wire_8561, wire_8531, wire_8501, wire_8471, wire_771, wire_280, wire_274, wire_265, wire_10689, wire_8559, wire_8529, wire_8499, wire_8469, wire_771, wire_280, wire_274, wire_265, wire_10687, wire_8557, wire_8527, wire_8497, wire_8467, wire_771, wire_280, wire_274, wire_265, wire_10685, wire_8555, wire_8525, wire_8495, wire_8465, wire_286, wire_280, wire_271, wire_265, wire_10683, wire_8553, wire_8523, wire_8493, wire_8463, wire_286, wire_280, wire_271, wire_265, wire_10681, wire_8551, wire_8521, wire_8491, wire_8461, wire_286, wire_280, wire_271, wire_265};
    // CHNAXY TOTAL: 30
    assign wire_10561 = io_tile_6_0_chanxy_out[0];
    assign wire_10563 = io_tile_6_0_chanxy_out[1];
    assign wire_10565 = io_tile_6_0_chanxy_out[2];
    assign wire_10567 = io_tile_6_0_chanxy_out[3];
    assign wire_10569 = io_tile_6_0_chanxy_out[4];
    assign wire_10571 = io_tile_6_0_chanxy_out[5];
    assign wire_10573 = io_tile_6_0_chanxy_out[6];
    assign wire_10575 = io_tile_6_0_chanxy_out[7];
    assign wire_10577 = io_tile_6_0_chanxy_out[8];
    assign wire_10579 = io_tile_6_0_chanxy_out[9];
    assign wire_10581 = io_tile_6_0_chanxy_out[10];
    assign wire_10583 = io_tile_6_0_chanxy_out[11];
    assign wire_10585 = io_tile_6_0_chanxy_out[12];
    assign wire_10587 = io_tile_6_0_chanxy_out[13];
    assign wire_10589 = io_tile_6_0_chanxy_out[14];
    assign wire_10650 = io_tile_6_0_chanxy_out[15];
    assign wire_10652 = io_tile_6_0_chanxy_out[16];
    assign wire_10654 = io_tile_6_0_chanxy_out[17];
    assign wire_10656 = io_tile_6_0_chanxy_out[18];
    assign wire_10658 = io_tile_6_0_chanxy_out[19];
    assign wire_10660 = io_tile_6_0_chanxy_out[20];
    assign wire_10662 = io_tile_6_0_chanxy_out[21];
    assign wire_10664 = io_tile_6_0_chanxy_out[22];
    assign wire_10666 = io_tile_6_0_chanxy_out[23];
    assign wire_10668 = io_tile_6_0_chanxy_out[24];
    assign wire_10670 = io_tile_6_0_chanxy_out[25];
    assign wire_10672 = io_tile_6_0_chanxy_out[26];
    assign wire_10674 = io_tile_6_0_chanxy_out[27];
    assign wire_10676 = io_tile_6_0_chanxy_out[28];
    assign wire_10678 = io_tile_6_0_chanxy_out[29];
    assign io_tile_7_0_chanxy_in = {wire_10588, wire_8579, wire_8549, wire_8519, wire_8489, wire_817, wire_334, wire_325, wire_319, wire_10586, wire_8577, wire_8547, wire_8517, wire_8487, wire_817, wire_334, wire_325, wire_319, wire_10584, wire_8575, wire_8545, wire_8515, wire_8485, wire_817, wire_334, wire_325, wire_319, wire_10582, wire_8573, wire_8543, wire_8513, wire_8483, wire_817, wire_331, wire_325, wire_316, wire_10580, wire_8571, wire_8541, wire_8511, wire_8481, wire_817, wire_331, wire_325, wire_316, wire_10578, wire_8569, wire_8539, wire_8509, wire_8479, wire_817, wire_331, wire_325, wire_316, wire_10576, wire_8567, wire_8537, wire_8507, wire_8477, wire_813, wire_331, wire_322, wire_316, wire_10574, wire_8565, wire_8535, wire_8505, wire_8475, wire_813, wire_331, wire_322, wire_316, wire_10572, wire_8563, wire_8533, wire_8503, wire_8473, wire_813, wire_331, wire_322, wire_316, wire_10570, wire_8561, wire_8531, wire_8501, wire_8471, wire_813, wire_328, wire_322, wire_313, wire_10568, wire_8559, wire_8529, wire_8499, wire_8469, wire_813, wire_328, wire_322, wire_313, wire_10566, wire_8557, wire_8527, wire_8497, wire_8467, wire_813, wire_328, wire_322, wire_313, wire_10564, wire_8555, wire_8525, wire_8495, wire_8465, wire_334, wire_328, wire_319, wire_313, wire_10562, wire_8553, wire_8523, wire_8493, wire_8463, wire_334, wire_328, wire_319, wire_313, wire_10560, wire_8551, wire_8521, wire_8491, wire_8461, wire_334, wire_328, wire_319, wire_313, wire_10739, wire_8969, wire_8939, wire_8909, wire_8879, wire_817, wire_334, wire_325, wire_319, wire_10737, wire_8967, wire_8937, wire_8907, wire_8877, wire_817, wire_334, wire_325, wire_319, wire_10735, wire_8965, wire_8935, wire_8905, wire_8875, wire_817, wire_334, wire_325, wire_319, wire_10733, wire_8963, wire_8933, wire_8903, wire_8873, wire_817, wire_331, wire_325, wire_316, wire_10731, wire_8961, wire_8931, wire_8901, wire_8871, wire_817, wire_331, wire_325, wire_316, wire_10729, wire_8959, wire_8929, wire_8899, wire_8869, wire_817, wire_331, wire_325, wire_316, wire_10727, wire_8957, wire_8927, wire_8897, wire_8867, wire_813, wire_331, wire_322, wire_316, wire_10725, wire_8955, wire_8925, wire_8895, wire_8865, wire_813, wire_331, wire_322, wire_316, wire_10723, wire_8953, wire_8923, wire_8893, wire_8863, wire_813, wire_331, wire_322, wire_316, wire_10721, wire_8951, wire_8921, wire_8891, wire_8861, wire_813, wire_328, wire_322, wire_313, wire_10719, wire_8949, wire_8919, wire_8889, wire_8859, wire_813, wire_328, wire_322, wire_313, wire_10717, wire_8947, wire_8917, wire_8887, wire_8857, wire_813, wire_328, wire_322, wire_313, wire_10715, wire_8945, wire_8915, wire_8885, wire_8855, wire_334, wire_328, wire_319, wire_313, wire_10713, wire_8943, wire_8913, wire_8883, wire_8853, wire_334, wire_328, wire_319, wire_313, wire_10711, wire_8941, wire_8911, wire_8881, wire_8851, wire_334, wire_328, wire_319, wire_313};
    // CHNAXY TOTAL: 30
    assign wire_10591 = io_tile_7_0_chanxy_out[0];
    assign wire_10593 = io_tile_7_0_chanxy_out[1];
    assign wire_10595 = io_tile_7_0_chanxy_out[2];
    assign wire_10597 = io_tile_7_0_chanxy_out[3];
    assign wire_10599 = io_tile_7_0_chanxy_out[4];
    assign wire_10601 = io_tile_7_0_chanxy_out[5];
    assign wire_10603 = io_tile_7_0_chanxy_out[6];
    assign wire_10605 = io_tile_7_0_chanxy_out[7];
    assign wire_10607 = io_tile_7_0_chanxy_out[8];
    assign wire_10609 = io_tile_7_0_chanxy_out[9];
    assign wire_10611 = io_tile_7_0_chanxy_out[10];
    assign wire_10613 = io_tile_7_0_chanxy_out[11];
    assign wire_10615 = io_tile_7_0_chanxy_out[12];
    assign wire_10617 = io_tile_7_0_chanxy_out[13];
    assign wire_10619 = io_tile_7_0_chanxy_out[14];
    assign wire_10680 = io_tile_7_0_chanxy_out[15];
    assign wire_10682 = io_tile_7_0_chanxy_out[16];
    assign wire_10684 = io_tile_7_0_chanxy_out[17];
    assign wire_10686 = io_tile_7_0_chanxy_out[18];
    assign wire_10688 = io_tile_7_0_chanxy_out[19];
    assign wire_10690 = io_tile_7_0_chanxy_out[20];
    assign wire_10692 = io_tile_7_0_chanxy_out[21];
    assign wire_10694 = io_tile_7_0_chanxy_out[22];
    assign wire_10696 = io_tile_7_0_chanxy_out[23];
    assign wire_10698 = io_tile_7_0_chanxy_out[24];
    assign wire_10700 = io_tile_7_0_chanxy_out[25];
    assign wire_10702 = io_tile_7_0_chanxy_out[26];
    assign wire_10704 = io_tile_7_0_chanxy_out[27];
    assign wire_10706 = io_tile_7_0_chanxy_out[28];
    assign wire_10708 = io_tile_7_0_chanxy_out[29];
    assign io_tile_8_0_chanxy_in = {wire_10618, wire_8969, wire_8939, wire_8909, wire_8879, wire_859, wire_382, wire_373, wire_367, wire_10616, wire_8967, wire_8937, wire_8907, wire_8877, wire_859, wire_382, wire_373, wire_367, wire_10614, wire_8965, wire_8935, wire_8905, wire_8875, wire_859, wire_382, wire_373, wire_367, wire_10612, wire_8963, wire_8933, wire_8903, wire_8873, wire_859, wire_379, wire_373, wire_364, wire_10610, wire_8961, wire_8931, wire_8901, wire_8871, wire_859, wire_379, wire_373, wire_364, wire_10608, wire_8959, wire_8929, wire_8899, wire_8869, wire_859, wire_379, wire_373, wire_364, wire_10606, wire_8957, wire_8927, wire_8897, wire_8867, wire_855, wire_379, wire_370, wire_364, wire_10604, wire_8955, wire_8925, wire_8895, wire_8865, wire_855, wire_379, wire_370, wire_364, wire_10602, wire_8953, wire_8923, wire_8893, wire_8863, wire_855, wire_379, wire_370, wire_364, wire_10600, wire_8951, wire_8921, wire_8891, wire_8861, wire_855, wire_376, wire_370, wire_361, wire_10598, wire_8949, wire_8919, wire_8889, wire_8859, wire_855, wire_376, wire_370, wire_361, wire_10596, wire_8947, wire_8917, wire_8887, wire_8857, wire_855, wire_376, wire_370, wire_361, wire_10594, wire_8945, wire_8915, wire_8885, wire_8855, wire_382, wire_376, wire_367, wire_361, wire_10592, wire_8943, wire_8913, wire_8883, wire_8853, wire_382, wire_376, wire_367, wire_361, wire_10590, wire_8941, wire_8911, wire_8881, wire_8851, wire_382, wire_376, wire_367, wire_361, wire_10769, wire_9359, wire_9329, wire_9299, wire_9269, wire_859, wire_382, wire_373, wire_367, wire_10767, wire_9357, wire_9327, wire_9297, wire_9267, wire_859, wire_382, wire_373, wire_367, wire_10765, wire_9355, wire_9325, wire_9295, wire_9265, wire_859, wire_382, wire_373, wire_367, wire_10763, wire_9353, wire_9323, wire_9293, wire_9263, wire_859, wire_379, wire_373, wire_364, wire_10761, wire_9351, wire_9321, wire_9291, wire_9261, wire_859, wire_379, wire_373, wire_364, wire_10759, wire_9349, wire_9319, wire_9289, wire_9259, wire_859, wire_379, wire_373, wire_364, wire_10757, wire_9347, wire_9317, wire_9287, wire_9257, wire_855, wire_379, wire_370, wire_364, wire_10755, wire_9345, wire_9315, wire_9285, wire_9255, wire_855, wire_379, wire_370, wire_364, wire_10753, wire_9343, wire_9313, wire_9283, wire_9253, wire_855, wire_379, wire_370, wire_364, wire_10751, wire_9341, wire_9311, wire_9281, wire_9251, wire_855, wire_376, wire_370, wire_361, wire_10749, wire_9339, wire_9309, wire_9279, wire_9249, wire_855, wire_376, wire_370, wire_361, wire_10747, wire_9337, wire_9307, wire_9277, wire_9247, wire_855, wire_376, wire_370, wire_361, wire_10745, wire_9335, wire_9305, wire_9275, wire_9245, wire_382, wire_376, wire_367, wire_361, wire_10743, wire_9333, wire_9303, wire_9273, wire_9243, wire_382, wire_376, wire_367, wire_361, wire_10741, wire_9331, wire_9301, wire_9271, wire_9241, wire_382, wire_376, wire_367, wire_361};
    // CHNAXY TOTAL: 30
    assign wire_10621 = io_tile_8_0_chanxy_out[0];
    assign wire_10623 = io_tile_8_0_chanxy_out[1];
    assign wire_10625 = io_tile_8_0_chanxy_out[2];
    assign wire_10627 = io_tile_8_0_chanxy_out[3];
    assign wire_10629 = io_tile_8_0_chanxy_out[4];
    assign wire_10631 = io_tile_8_0_chanxy_out[5];
    assign wire_10633 = io_tile_8_0_chanxy_out[6];
    assign wire_10635 = io_tile_8_0_chanxy_out[7];
    assign wire_10637 = io_tile_8_0_chanxy_out[8];
    assign wire_10639 = io_tile_8_0_chanxy_out[9];
    assign wire_10641 = io_tile_8_0_chanxy_out[10];
    assign wire_10643 = io_tile_8_0_chanxy_out[11];
    assign wire_10645 = io_tile_8_0_chanxy_out[12];
    assign wire_10647 = io_tile_8_0_chanxy_out[13];
    assign wire_10649 = io_tile_8_0_chanxy_out[14];
    assign wire_10710 = io_tile_8_0_chanxy_out[15];
    assign wire_10712 = io_tile_8_0_chanxy_out[16];
    assign wire_10714 = io_tile_8_0_chanxy_out[17];
    assign wire_10716 = io_tile_8_0_chanxy_out[18];
    assign wire_10718 = io_tile_8_0_chanxy_out[19];
    assign wire_10720 = io_tile_8_0_chanxy_out[20];
    assign wire_10722 = io_tile_8_0_chanxy_out[21];
    assign wire_10724 = io_tile_8_0_chanxy_out[22];
    assign wire_10726 = io_tile_8_0_chanxy_out[23];
    assign wire_10728 = io_tile_8_0_chanxy_out[24];
    assign wire_10730 = io_tile_8_0_chanxy_out[25];
    assign wire_10732 = io_tile_8_0_chanxy_out[26];
    assign wire_10734 = io_tile_8_0_chanxy_out[27];
    assign wire_10736 = io_tile_8_0_chanxy_out[28];
    assign wire_10738 = io_tile_8_0_chanxy_out[29];
    assign io_tile_9_0_chanxy_in = {wire_10648, wire_9359, wire_9329, wire_9299, wire_9269, wire_901, wire_430, wire_421, wire_415, wire_10646, wire_9357, wire_9327, wire_9297, wire_9267, wire_901, wire_430, wire_421, wire_415, wire_10644, wire_9355, wire_9325, wire_9295, wire_9265, wire_901, wire_430, wire_421, wire_415, wire_10642, wire_9353, wire_9323, wire_9293, wire_9263, wire_901, wire_427, wire_421, wire_412, wire_10640, wire_9351, wire_9321, wire_9291, wire_9261, wire_901, wire_427, wire_421, wire_412, wire_10638, wire_9349, wire_9319, wire_9289, wire_9259, wire_901, wire_427, wire_421, wire_412, wire_10636, wire_9347, wire_9317, wire_9287, wire_9257, wire_897, wire_427, wire_418, wire_412, wire_10634, wire_9345, wire_9315, wire_9285, wire_9255, wire_897, wire_427, wire_418, wire_412, wire_10632, wire_9343, wire_9313, wire_9283, wire_9253, wire_897, wire_427, wire_418, wire_412, wire_10630, wire_9341, wire_9311, wire_9281, wire_9251, wire_897, wire_424, wire_418, wire_409, wire_10628, wire_9339, wire_9309, wire_9279, wire_9249, wire_897, wire_424, wire_418, wire_409, wire_10626, wire_9337, wire_9307, wire_9277, wire_9247, wire_897, wire_424, wire_418, wire_409, wire_10624, wire_9335, wire_9305, wire_9275, wire_9245, wire_430, wire_424, wire_415, wire_409, wire_10622, wire_9333, wire_9303, wire_9273, wire_9243, wire_430, wire_424, wire_415, wire_409, wire_10620, wire_9331, wire_9301, wire_9271, wire_9241, wire_430, wire_424, wire_415, wire_409, wire_10799, wire_9749, wire_9719, wire_9689, wire_9659, wire_901, wire_430, wire_421, wire_415, wire_10797, wire_9747, wire_9717, wire_9687, wire_9657, wire_901, wire_430, wire_421, wire_415, wire_10795, wire_9745, wire_9715, wire_9685, wire_9655, wire_901, wire_430, wire_421, wire_415, wire_10793, wire_9743, wire_9713, wire_9683, wire_9653, wire_901, wire_427, wire_421, wire_412, wire_10791, wire_9741, wire_9711, wire_9681, wire_9651, wire_901, wire_427, wire_421, wire_412, wire_10789, wire_9739, wire_9709, wire_9679, wire_9649, wire_901, wire_427, wire_421, wire_412, wire_10787, wire_9737, wire_9707, wire_9677, wire_9647, wire_897, wire_427, wire_418, wire_412, wire_10785, wire_9735, wire_9705, wire_9675, wire_9645, wire_897, wire_427, wire_418, wire_412, wire_10783, wire_9733, wire_9703, wire_9673, wire_9643, wire_897, wire_427, wire_418, wire_412, wire_10781, wire_9731, wire_9701, wire_9671, wire_9641, wire_897, wire_424, wire_418, wire_409, wire_10779, wire_9729, wire_9699, wire_9669, wire_9639, wire_897, wire_424, wire_418, wire_409, wire_10777, wire_9727, wire_9697, wire_9667, wire_9637, wire_897, wire_424, wire_418, wire_409, wire_10775, wire_9725, wire_9695, wire_9665, wire_9635, wire_430, wire_424, wire_415, wire_409, wire_10773, wire_9723, wire_9693, wire_9663, wire_9633, wire_430, wire_424, wire_415, wire_409, wire_10771, wire_9721, wire_9691, wire_9661, wire_9631, wire_430, wire_424, wire_415, wire_409};
    // CHNAXY TOTAL: 30
    assign wire_10651 = io_tile_9_0_chanxy_out[0];
    assign wire_10653 = io_tile_9_0_chanxy_out[1];
    assign wire_10655 = io_tile_9_0_chanxy_out[2];
    assign wire_10657 = io_tile_9_0_chanxy_out[3];
    assign wire_10659 = io_tile_9_0_chanxy_out[4];
    assign wire_10661 = io_tile_9_0_chanxy_out[5];
    assign wire_10663 = io_tile_9_0_chanxy_out[6];
    assign wire_10665 = io_tile_9_0_chanxy_out[7];
    assign wire_10667 = io_tile_9_0_chanxy_out[8];
    assign wire_10669 = io_tile_9_0_chanxy_out[9];
    assign wire_10671 = io_tile_9_0_chanxy_out[10];
    assign wire_10673 = io_tile_9_0_chanxy_out[11];
    assign wire_10675 = io_tile_9_0_chanxy_out[12];
    assign wire_10677 = io_tile_9_0_chanxy_out[13];
    assign wire_10679 = io_tile_9_0_chanxy_out[14];
    assign wire_10740 = io_tile_9_0_chanxy_out[15];
    assign wire_10742 = io_tile_9_0_chanxy_out[16];
    assign wire_10744 = io_tile_9_0_chanxy_out[17];
    assign wire_10746 = io_tile_9_0_chanxy_out[18];
    assign wire_10748 = io_tile_9_0_chanxy_out[19];
    assign wire_10750 = io_tile_9_0_chanxy_out[20];
    assign wire_10752 = io_tile_9_0_chanxy_out[21];
    assign wire_10754 = io_tile_9_0_chanxy_out[22];
    assign wire_10756 = io_tile_9_0_chanxy_out[23];
    assign wire_10758 = io_tile_9_0_chanxy_out[24];
    assign wire_10760 = io_tile_9_0_chanxy_out[25];
    assign wire_10762 = io_tile_9_0_chanxy_out[26];
    assign wire_10764 = io_tile_9_0_chanxy_out[27];
    assign wire_10766 = io_tile_9_0_chanxy_out[28];
    assign wire_10768 = io_tile_9_0_chanxy_out[29];
    assign io_tile_10_0_chanxy_in = {wire_10023, wire_943, wire_10678, wire_9749, wire_9719, wire_9689, wire_9659, wire_943, wire_478, wire_469, wire_463, wire_10031, wire_939, wire_10676, wire_9747, wire_9717, wire_9687, wire_9657, wire_943, wire_478, wire_469, wire_463, wire_10039, wire_939, wire_10674, wire_9745, wire_9715, wire_9685, wire_9655, wire_943, wire_478, wire_469, wire_463, wire_10047, wire_478, wire_10672, wire_9743, wire_9713, wire_9683, wire_9653, wire_943, wire_475, wire_469, wire_460, wire_10055, wire_475, wire_10670, wire_9741, wire_9711, wire_9681, wire_9651, wire_943, wire_475, wire_469, wire_460, wire_10063, wire_475, wire_10668, wire_9739, wire_9709, wire_9679, wire_9649, wire_943, wire_475, wire_469, wire_460, wire_10071, wire_472, wire_10666, wire_9737, wire_9707, wire_9677, wire_9647, wire_939, wire_475, wire_466, wire_460, wire_10079, wire_469, wire_10664, wire_9735, wire_9705, wire_9675, wire_9645, wire_939, wire_475, wire_466, wire_460, wire_10087, wire_469, wire_10662, wire_9733, wire_9703, wire_9673, wire_9643, wire_939, wire_475, wire_466, wire_460, wire_10095, wire_466, wire_10660, wire_9731, wire_9701, wire_9671, wire_9641, wire_939, wire_472, wire_466, wire_457, wire_10103, wire_463, wire_10658, wire_9729, wire_9699, wire_9669, wire_9639, wire_939, wire_472, wire_466, wire_457, wire_10111, wire_463, wire_10656, wire_9727, wire_9697, wire_9667, wire_9637, wire_939, wire_472, wire_466, wire_457, wire_10119, wire_460, wire_10654, wire_9725, wire_9695, wire_9665, wire_9635, wire_478, wire_472, wire_463, wire_457, wire_10127, wire_457, wire_10652, wire_9723, wire_9693, wire_9663, wire_9633, wire_478, wire_472, wire_463, wire_457, wire_10135, wire_457, wire_10650, wire_9721, wire_9691, wire_9661, wire_9631, wire_478, wire_472, wire_463, wire_457, wire_10025, wire_943, wire_10033, wire_939, wire_10041, wire_939, wire_10049, wire_478, wire_10057, wire_475, wire_10065, wire_475, wire_10073, wire_472, wire_10081, wire_469, wire_10089, wire_469, wire_10097, wire_466, wire_10105, wire_463, wire_10113, wire_463, wire_10121, wire_460, wire_10129, wire_457, wire_10137, wire_457, wire_10139, wire_943, wire_10027, wire_943, wire_10035, wire_939, wire_10043, wire_478, wire_10051, wire_478, wire_10059, wire_475, wire_10067, wire_472, wire_10075, wire_472, wire_10083, wire_469, wire_10091, wire_466, wire_10099, wire_466, wire_10107, wire_463, wire_10115, wire_460, wire_10123, wire_460, wire_10131, wire_457, wire_10021, wire_943, wire_10029, wire_943, wire_10037, wire_939, wire_10045, wire_478, wire_10053, wire_478, wire_10061, wire_475, wire_10069, wire_472, wire_10077, wire_472, wire_10085, wire_469, wire_10093, wire_466, wire_10101, wire_466, wire_10109, wire_463, wire_10117, wire_460, wire_10125, wire_460, wire_10133, wire_457};
    // CHNAXY TOTAL: 75
    assign wire_10681 = io_tile_10_0_chanxy_out[0];
    assign wire_10683 = io_tile_10_0_chanxy_out[1];
    assign wire_10685 = io_tile_10_0_chanxy_out[2];
    assign wire_10687 = io_tile_10_0_chanxy_out[3];
    assign wire_10689 = io_tile_10_0_chanxy_out[4];
    assign wire_10691 = io_tile_10_0_chanxy_out[5];
    assign wire_10693 = io_tile_10_0_chanxy_out[6];
    assign wire_10695 = io_tile_10_0_chanxy_out[7];
    assign wire_10697 = io_tile_10_0_chanxy_out[8];
    assign wire_10699 = io_tile_10_0_chanxy_out[9];
    assign wire_10701 = io_tile_10_0_chanxy_out[10];
    assign wire_10703 = io_tile_10_0_chanxy_out[11];
    assign wire_10705 = io_tile_10_0_chanxy_out[12];
    assign wire_10707 = io_tile_10_0_chanxy_out[13];
    assign wire_10709 = io_tile_10_0_chanxy_out[14];
    assign wire_10711 = io_tile_10_0_chanxy_out[15];
    assign wire_10713 = io_tile_10_0_chanxy_out[16];
    assign wire_10715 = io_tile_10_0_chanxy_out[17];
    assign wire_10717 = io_tile_10_0_chanxy_out[18];
    assign wire_10719 = io_tile_10_0_chanxy_out[19];
    assign wire_10721 = io_tile_10_0_chanxy_out[20];
    assign wire_10723 = io_tile_10_0_chanxy_out[21];
    assign wire_10725 = io_tile_10_0_chanxy_out[22];
    assign wire_10727 = io_tile_10_0_chanxy_out[23];
    assign wire_10729 = io_tile_10_0_chanxy_out[24];
    assign wire_10731 = io_tile_10_0_chanxy_out[25];
    assign wire_10733 = io_tile_10_0_chanxy_out[26];
    assign wire_10735 = io_tile_10_0_chanxy_out[27];
    assign wire_10737 = io_tile_10_0_chanxy_out[28];
    assign wire_10739 = io_tile_10_0_chanxy_out[29];
    assign wire_10741 = io_tile_10_0_chanxy_out[30];
    assign wire_10743 = io_tile_10_0_chanxy_out[31];
    assign wire_10745 = io_tile_10_0_chanxy_out[32];
    assign wire_10747 = io_tile_10_0_chanxy_out[33];
    assign wire_10749 = io_tile_10_0_chanxy_out[34];
    assign wire_10751 = io_tile_10_0_chanxy_out[35];
    assign wire_10753 = io_tile_10_0_chanxy_out[36];
    assign wire_10755 = io_tile_10_0_chanxy_out[37];
    assign wire_10757 = io_tile_10_0_chanxy_out[38];
    assign wire_10759 = io_tile_10_0_chanxy_out[39];
    assign wire_10761 = io_tile_10_0_chanxy_out[40];
    assign wire_10763 = io_tile_10_0_chanxy_out[41];
    assign wire_10765 = io_tile_10_0_chanxy_out[42];
    assign wire_10767 = io_tile_10_0_chanxy_out[43];
    assign wire_10769 = io_tile_10_0_chanxy_out[44];
    assign wire_10770 = io_tile_10_0_chanxy_out[45];
    assign wire_10771 = io_tile_10_0_chanxy_out[46];
    assign wire_10772 = io_tile_10_0_chanxy_out[47];
    assign wire_10773 = io_tile_10_0_chanxy_out[48];
    assign wire_10774 = io_tile_10_0_chanxy_out[49];
    assign wire_10775 = io_tile_10_0_chanxy_out[50];
    assign wire_10776 = io_tile_10_0_chanxy_out[51];
    assign wire_10777 = io_tile_10_0_chanxy_out[52];
    assign wire_10778 = io_tile_10_0_chanxy_out[53];
    assign wire_10779 = io_tile_10_0_chanxy_out[54];
    assign wire_10780 = io_tile_10_0_chanxy_out[55];
    assign wire_10781 = io_tile_10_0_chanxy_out[56];
    assign wire_10782 = io_tile_10_0_chanxy_out[57];
    assign wire_10783 = io_tile_10_0_chanxy_out[58];
    assign wire_10784 = io_tile_10_0_chanxy_out[59];
    assign wire_10785 = io_tile_10_0_chanxy_out[60];
    assign wire_10786 = io_tile_10_0_chanxy_out[61];
    assign wire_10787 = io_tile_10_0_chanxy_out[62];
    assign wire_10788 = io_tile_10_0_chanxy_out[63];
    assign wire_10789 = io_tile_10_0_chanxy_out[64];
    assign wire_10790 = io_tile_10_0_chanxy_out[65];
    assign wire_10791 = io_tile_10_0_chanxy_out[66];
    assign wire_10792 = io_tile_10_0_chanxy_out[67];
    assign wire_10793 = io_tile_10_0_chanxy_out[68];
    assign wire_10794 = io_tile_10_0_chanxy_out[69];
    assign wire_10795 = io_tile_10_0_chanxy_out[70];
    assign wire_10796 = io_tile_10_0_chanxy_out[71];
    assign wire_10797 = io_tile_10_0_chanxy_out[72];
    assign wire_10798 = io_tile_10_0_chanxy_out[73];
    assign wire_10799 = io_tile_10_0_chanxy_out[74];
    assign io_tile_0_1_chanxy_in = {wire_10527, wire_568, wire_10525, wire_568, wire_10919, wire_10889, wire_10859, wire_10829, wire_6269, wire_568, wire_526, wire_517, wire_511, wire_10523, wire_568, wire_10521, wire_568, wire_10519, wire_568, wire_10517, wire_568, wire_10917, wire_10887, wire_10857, wire_10827, wire_6267, wire_568, wire_526, wire_517, wire_511, wire_10515, wire_564, wire_10513, wire_564, wire_10511, wire_564, wire_10509, wire_564, wire_10915, wire_10885, wire_10855, wire_10825, wire_6265, wire_568, wire_526, wire_517, wire_511, wire_10507, wire_564, wire_10505, wire_564, wire_10503, wire_526, wire_10501, wire_526, wire_10913, wire_10883, wire_10853, wire_10823, wire_6263, wire_568, wire_523, wire_517, wire_508, wire_10499, wire_526, wire_10497, wire_526, wire_10495, wire_526, wire_10493, wire_526, wire_10911, wire_10881, wire_10851, wire_10821, wire_6261, wire_568, wire_523, wire_517, wire_508, wire_10491, wire_523, wire_10489, wire_523, wire_10487, wire_523, wire_10485, wire_523, wire_10909, wire_10879, wire_10849, wire_10819, wire_6259, wire_568, wire_523, wire_517, wire_508, wire_10483, wire_523, wire_10481, wire_523, wire_10479, wire_520, wire_10477, wire_520, wire_10907, wire_10877, wire_10847, wire_10817, wire_6257, wire_564, wire_523, wire_514, wire_508, wire_10475, wire_520, wire_10473, wire_520, wire_10471, wire_520, wire_10469, wire_520, wire_10905, wire_10875, wire_10845, wire_10815, wire_6255, wire_564, wire_523, wire_514, wire_508, wire_10467, wire_517, wire_10465, wire_517, wire_10463, wire_517, wire_10461, wire_517, wire_10903, wire_10873, wire_10843, wire_10813, wire_6253, wire_564, wire_523, wire_514, wire_508, wire_10459, wire_517, wire_10457, wire_517, wire_10455, wire_514, wire_10453, wire_514, wire_10901, wire_10871, wire_10841, wire_10811, wire_6251, wire_564, wire_520, wire_514, wire_505, wire_10451, wire_514, wire_10449, wire_514, wire_10447, wire_514, wire_10445, wire_514, wire_10899, wire_10869, wire_10839, wire_10809, wire_6249, wire_564, wire_520, wire_514, wire_505, wire_10443, wire_511, wire_10441, wire_511, wire_10439, wire_511, wire_10437, wire_511, wire_10897, wire_10867, wire_10837, wire_10807, wire_6247, wire_564, wire_520, wire_514, wire_505, wire_10435, wire_511, wire_10433, wire_511, wire_10431, wire_508, wire_10429, wire_508, wire_10895, wire_10865, wire_10835, wire_10805, wire_6245, wire_526, wire_520, wire_511, wire_505, wire_10427, wire_508, wire_10425, wire_508, wire_10423, wire_508, wire_10421, wire_508, wire_10893, wire_10863, wire_10833, wire_10803, wire_6243, wire_526, wire_520, wire_511, wire_505, wire_10419, wire_505, wire_10417, wire_505, wire_10415, wire_505, wire_10413, wire_505, wire_10891, wire_10861, wire_10831, wire_10801, wire_6241, wire_526, wire_520, wire_511, wire_505, wire_10411, wire_505, wire_10529, wire_505};
    // CHNAXY TOTAL: 75
    assign wire_6120 = io_tile_0_1_chanxy_out[0];
    assign wire_6122 = io_tile_0_1_chanxy_out[1];
    assign wire_6123 = io_tile_0_1_chanxy_out[2];
    assign wire_6124 = io_tile_0_1_chanxy_out[3];
    assign wire_6126 = io_tile_0_1_chanxy_out[4];
    assign wire_6128 = io_tile_0_1_chanxy_out[5];
    assign wire_6130 = io_tile_0_1_chanxy_out[6];
    assign wire_6131 = io_tile_0_1_chanxy_out[7];
    assign wire_6132 = io_tile_0_1_chanxy_out[8];
    assign wire_6134 = io_tile_0_1_chanxy_out[9];
    assign wire_6136 = io_tile_0_1_chanxy_out[10];
    assign wire_6138 = io_tile_0_1_chanxy_out[11];
    assign wire_6139 = io_tile_0_1_chanxy_out[12];
    assign wire_6140 = io_tile_0_1_chanxy_out[13];
    assign wire_6142 = io_tile_0_1_chanxy_out[14];
    assign wire_6144 = io_tile_0_1_chanxy_out[15];
    assign wire_6146 = io_tile_0_1_chanxy_out[16];
    assign wire_6147 = io_tile_0_1_chanxy_out[17];
    assign wire_6148 = io_tile_0_1_chanxy_out[18];
    assign wire_6150 = io_tile_0_1_chanxy_out[19];
    assign wire_6152 = io_tile_0_1_chanxy_out[20];
    assign wire_6154 = io_tile_0_1_chanxy_out[21];
    assign wire_6155 = io_tile_0_1_chanxy_out[22];
    assign wire_6156 = io_tile_0_1_chanxy_out[23];
    assign wire_6158 = io_tile_0_1_chanxy_out[24];
    assign wire_6160 = io_tile_0_1_chanxy_out[25];
    assign wire_6162 = io_tile_0_1_chanxy_out[26];
    assign wire_6163 = io_tile_0_1_chanxy_out[27];
    assign wire_6164 = io_tile_0_1_chanxy_out[28];
    assign wire_6166 = io_tile_0_1_chanxy_out[29];
    assign wire_6168 = io_tile_0_1_chanxy_out[30];
    assign wire_6170 = io_tile_0_1_chanxy_out[31];
    assign wire_6171 = io_tile_0_1_chanxy_out[32];
    assign wire_6172 = io_tile_0_1_chanxy_out[33];
    assign wire_6174 = io_tile_0_1_chanxy_out[34];
    assign wire_6176 = io_tile_0_1_chanxy_out[35];
    assign wire_6178 = io_tile_0_1_chanxy_out[36];
    assign wire_6179 = io_tile_0_1_chanxy_out[37];
    assign wire_6180 = io_tile_0_1_chanxy_out[38];
    assign wire_6182 = io_tile_0_1_chanxy_out[39];
    assign wire_6184 = io_tile_0_1_chanxy_out[40];
    assign wire_6186 = io_tile_0_1_chanxy_out[41];
    assign wire_6187 = io_tile_0_1_chanxy_out[42];
    assign wire_6188 = io_tile_0_1_chanxy_out[43];
    assign wire_6190 = io_tile_0_1_chanxy_out[44];
    assign wire_6192 = io_tile_0_1_chanxy_out[45];
    assign wire_6194 = io_tile_0_1_chanxy_out[46];
    assign wire_6195 = io_tile_0_1_chanxy_out[47];
    assign wire_6196 = io_tile_0_1_chanxy_out[48];
    assign wire_6198 = io_tile_0_1_chanxy_out[49];
    assign wire_6200 = io_tile_0_1_chanxy_out[50];
    assign wire_6202 = io_tile_0_1_chanxy_out[51];
    assign wire_6203 = io_tile_0_1_chanxy_out[52];
    assign wire_6204 = io_tile_0_1_chanxy_out[53];
    assign wire_6206 = io_tile_0_1_chanxy_out[54];
    assign wire_6208 = io_tile_0_1_chanxy_out[55];
    assign wire_6210 = io_tile_0_1_chanxy_out[56];
    assign wire_6211 = io_tile_0_1_chanxy_out[57];
    assign wire_6212 = io_tile_0_1_chanxy_out[58];
    assign wire_6214 = io_tile_0_1_chanxy_out[59];
    assign wire_6216 = io_tile_0_1_chanxy_out[60];
    assign wire_6218 = io_tile_0_1_chanxy_out[61];
    assign wire_6219 = io_tile_0_1_chanxy_out[62];
    assign wire_6220 = io_tile_0_1_chanxy_out[63];
    assign wire_6222 = io_tile_0_1_chanxy_out[64];
    assign wire_6224 = io_tile_0_1_chanxy_out[65];
    assign wire_6226 = io_tile_0_1_chanxy_out[66];
    assign wire_6227 = io_tile_0_1_chanxy_out[67];
    assign wire_6228 = io_tile_0_1_chanxy_out[68];
    assign wire_6230 = io_tile_0_1_chanxy_out[69];
    assign wire_6232 = io_tile_0_1_chanxy_out[70];
    assign wire_6234 = io_tile_0_1_chanxy_out[71];
    assign wire_6235 = io_tile_0_1_chanxy_out[72];
    assign wire_6236 = io_tile_0_1_chanxy_out[73];
    assign wire_6238 = io_tile_0_1_chanxy_out[74];
    assign io_tile_0_2_chanxy_in = {wire_10919, wire_10889, wire_10859, wire_10829, wire_6234, wire_1084, wire_1042, wire_1033, wire_1027, wire_10917, wire_10887, wire_10857, wire_10827, wire_6226, wire_1084, wire_1042, wire_1033, wire_1027, wire_10915, wire_10885, wire_10855, wire_10825, wire_6218, wire_1084, wire_1042, wire_1033, wire_1027, wire_10913, wire_10883, wire_10853, wire_10823, wire_6210, wire_1084, wire_1039, wire_1033, wire_1024, wire_10911, wire_10881, wire_10851, wire_10821, wire_6202, wire_1084, wire_1039, wire_1033, wire_1024, wire_10909, wire_10879, wire_10849, wire_10819, wire_6194, wire_1084, wire_1039, wire_1033, wire_1024, wire_10907, wire_10877, wire_10847, wire_10817, wire_6186, wire_1080, wire_1039, wire_1030, wire_1024, wire_10905, wire_10875, wire_10845, wire_10815, wire_6178, wire_1080, wire_1039, wire_1030, wire_1024, wire_10903, wire_10873, wire_10843, wire_10813, wire_6170, wire_1080, wire_1039, wire_1030, wire_1024, wire_10901, wire_10871, wire_10841, wire_10811, wire_6162, wire_1080, wire_1036, wire_1030, wire_1021, wire_10899, wire_10869, wire_10839, wire_10809, wire_6154, wire_1080, wire_1036, wire_1030, wire_1021, wire_10897, wire_10867, wire_10837, wire_10807, wire_6146, wire_1080, wire_1036, wire_1030, wire_1021, wire_10895, wire_10865, wire_10835, wire_10805, wire_6138, wire_1042, wire_1036, wire_1027, wire_1021, wire_10893, wire_10863, wire_10833, wire_10803, wire_6130, wire_1042, wire_1036, wire_1027, wire_1021, wire_10891, wire_10861, wire_10831, wire_10801, wire_6122, wire_1042, wire_1036, wire_1027, wire_1021, wire_11309, wire_11279, wire_11249, wire_11219, wire_6299, wire_1084, wire_1042, wire_1033, wire_1027, wire_11307, wire_11277, wire_11247, wire_11217, wire_6297, wire_1084, wire_1042, wire_1033, wire_1027, wire_11305, wire_11275, wire_11245, wire_11215, wire_6295, wire_1084, wire_1042, wire_1033, wire_1027, wire_11303, wire_11273, wire_11243, wire_11213, wire_6293, wire_1084, wire_1039, wire_1033, wire_1024, wire_11301, wire_11271, wire_11241, wire_11211, wire_6291, wire_1084, wire_1039, wire_1033, wire_1024, wire_11299, wire_11269, wire_11239, wire_11209, wire_6289, wire_1084, wire_1039, wire_1033, wire_1024, wire_11297, wire_11267, wire_11237, wire_11207, wire_6287, wire_1080, wire_1039, wire_1030, wire_1024, wire_11295, wire_11265, wire_11235, wire_11205, wire_6285, wire_1080, wire_1039, wire_1030, wire_1024, wire_11293, wire_11263, wire_11233, wire_11203, wire_6283, wire_1080, wire_1039, wire_1030, wire_1024, wire_11291, wire_11261, wire_11231, wire_11201, wire_6281, wire_1080, wire_1036, wire_1030, wire_1021, wire_11289, wire_11259, wire_11229, wire_11199, wire_6279, wire_1080, wire_1036, wire_1030, wire_1021, wire_11287, wire_11257, wire_11227, wire_11197, wire_6277, wire_1080, wire_1036, wire_1030, wire_1021, wire_11285, wire_11255, wire_11225, wire_11195, wire_6275, wire_1042, wire_1036, wire_1027, wire_1021, wire_11283, wire_11253, wire_11223, wire_11193, wire_6273, wire_1042, wire_1036, wire_1027, wire_1021, wire_11281, wire_11251, wire_11221, wire_11191, wire_6271, wire_1042, wire_1036, wire_1027, wire_1021};
    // CHNAXY TOTAL: 30
    assign wire_6125 = io_tile_0_2_chanxy_out[0];
    assign wire_6133 = io_tile_0_2_chanxy_out[1];
    assign wire_6141 = io_tile_0_2_chanxy_out[2];
    assign wire_6149 = io_tile_0_2_chanxy_out[3];
    assign wire_6157 = io_tile_0_2_chanxy_out[4];
    assign wire_6165 = io_tile_0_2_chanxy_out[5];
    assign wire_6173 = io_tile_0_2_chanxy_out[6];
    assign wire_6181 = io_tile_0_2_chanxy_out[7];
    assign wire_6189 = io_tile_0_2_chanxy_out[8];
    assign wire_6197 = io_tile_0_2_chanxy_out[9];
    assign wire_6205 = io_tile_0_2_chanxy_out[10];
    assign wire_6213 = io_tile_0_2_chanxy_out[11];
    assign wire_6221 = io_tile_0_2_chanxy_out[12];
    assign wire_6229 = io_tile_0_2_chanxy_out[13];
    assign wire_6237 = io_tile_0_2_chanxy_out[14];
    assign wire_6240 = io_tile_0_2_chanxy_out[15];
    assign wire_6242 = io_tile_0_2_chanxy_out[16];
    assign wire_6244 = io_tile_0_2_chanxy_out[17];
    assign wire_6246 = io_tile_0_2_chanxy_out[18];
    assign wire_6248 = io_tile_0_2_chanxy_out[19];
    assign wire_6250 = io_tile_0_2_chanxy_out[20];
    assign wire_6252 = io_tile_0_2_chanxy_out[21];
    assign wire_6254 = io_tile_0_2_chanxy_out[22];
    assign wire_6256 = io_tile_0_2_chanxy_out[23];
    assign wire_6258 = io_tile_0_2_chanxy_out[24];
    assign wire_6260 = io_tile_0_2_chanxy_out[25];
    assign wire_6262 = io_tile_0_2_chanxy_out[26];
    assign wire_6264 = io_tile_0_2_chanxy_out[27];
    assign wire_6266 = io_tile_0_2_chanxy_out[28];
    assign wire_6268 = io_tile_0_2_chanxy_out[29];
    assign io_tile_0_3_chanxy_in = {wire_11309, wire_11279, wire_11249, wire_11219, wire_6236, wire_1600, wire_1558, wire_1549, wire_1543, wire_11307, wire_11277, wire_11247, wire_11217, wire_6228, wire_1600, wire_1558, wire_1549, wire_1543, wire_11305, wire_11275, wire_11245, wire_11215, wire_6220, wire_1600, wire_1558, wire_1549, wire_1543, wire_11303, wire_11273, wire_11243, wire_11213, wire_6212, wire_1600, wire_1555, wire_1549, wire_1540, wire_11301, wire_11271, wire_11241, wire_11211, wire_6204, wire_1600, wire_1555, wire_1549, wire_1540, wire_11299, wire_11269, wire_11239, wire_11209, wire_6196, wire_1600, wire_1555, wire_1549, wire_1540, wire_11297, wire_11267, wire_11237, wire_11207, wire_6188, wire_1596, wire_1555, wire_1546, wire_1540, wire_11295, wire_11265, wire_11235, wire_11205, wire_6180, wire_1596, wire_1555, wire_1546, wire_1540, wire_11293, wire_11263, wire_11233, wire_11203, wire_6172, wire_1596, wire_1555, wire_1546, wire_1540, wire_11291, wire_11261, wire_11231, wire_11201, wire_6164, wire_1596, wire_1552, wire_1546, wire_1537, wire_11289, wire_11259, wire_11229, wire_11199, wire_6156, wire_1596, wire_1552, wire_1546, wire_1537, wire_11287, wire_11257, wire_11227, wire_11197, wire_6148, wire_1596, wire_1552, wire_1546, wire_1537, wire_11285, wire_11255, wire_11225, wire_11195, wire_6140, wire_1558, wire_1552, wire_1543, wire_1537, wire_11283, wire_11253, wire_11223, wire_11193, wire_6132, wire_1558, wire_1552, wire_1543, wire_1537, wire_11281, wire_11251, wire_11221, wire_11191, wire_6124, wire_1558, wire_1552, wire_1543, wire_1537, wire_11699, wire_11669, wire_11639, wire_11609, wire_6329, wire_1600, wire_1558, wire_1549, wire_1543, wire_11697, wire_11667, wire_11637, wire_11607, wire_6327, wire_1600, wire_1558, wire_1549, wire_1543, wire_11695, wire_11665, wire_11635, wire_11605, wire_6325, wire_1600, wire_1558, wire_1549, wire_1543, wire_11693, wire_11663, wire_11633, wire_11603, wire_6323, wire_1600, wire_1555, wire_1549, wire_1540, wire_11691, wire_11661, wire_11631, wire_11601, wire_6321, wire_1600, wire_1555, wire_1549, wire_1540, wire_11689, wire_11659, wire_11629, wire_11599, wire_6319, wire_1600, wire_1555, wire_1549, wire_1540, wire_11687, wire_11657, wire_11627, wire_11597, wire_6317, wire_1596, wire_1555, wire_1546, wire_1540, wire_11685, wire_11655, wire_11625, wire_11595, wire_6315, wire_1596, wire_1555, wire_1546, wire_1540, wire_11683, wire_11653, wire_11623, wire_11593, wire_6313, wire_1596, wire_1555, wire_1546, wire_1540, wire_11681, wire_11651, wire_11621, wire_11591, wire_6311, wire_1596, wire_1552, wire_1546, wire_1537, wire_11679, wire_11649, wire_11619, wire_11589, wire_6309, wire_1596, wire_1552, wire_1546, wire_1537, wire_11677, wire_11647, wire_11617, wire_11587, wire_6307, wire_1596, wire_1552, wire_1546, wire_1537, wire_11675, wire_11645, wire_11615, wire_11585, wire_6305, wire_1558, wire_1552, wire_1543, wire_1537, wire_11673, wire_11643, wire_11613, wire_11583, wire_6303, wire_1558, wire_1552, wire_1543, wire_1537, wire_11671, wire_11641, wire_11611, wire_11581, wire_6301, wire_1558, wire_1552, wire_1543, wire_1537};
    // CHNAXY TOTAL: 30
    assign wire_6127 = io_tile_0_3_chanxy_out[0];
    assign wire_6135 = io_tile_0_3_chanxy_out[1];
    assign wire_6143 = io_tile_0_3_chanxy_out[2];
    assign wire_6151 = io_tile_0_3_chanxy_out[3];
    assign wire_6159 = io_tile_0_3_chanxy_out[4];
    assign wire_6167 = io_tile_0_3_chanxy_out[5];
    assign wire_6175 = io_tile_0_3_chanxy_out[6];
    assign wire_6183 = io_tile_0_3_chanxy_out[7];
    assign wire_6191 = io_tile_0_3_chanxy_out[8];
    assign wire_6199 = io_tile_0_3_chanxy_out[9];
    assign wire_6207 = io_tile_0_3_chanxy_out[10];
    assign wire_6215 = io_tile_0_3_chanxy_out[11];
    assign wire_6223 = io_tile_0_3_chanxy_out[12];
    assign wire_6231 = io_tile_0_3_chanxy_out[13];
    assign wire_6239 = io_tile_0_3_chanxy_out[14];
    assign wire_6270 = io_tile_0_3_chanxy_out[15];
    assign wire_6272 = io_tile_0_3_chanxy_out[16];
    assign wire_6274 = io_tile_0_3_chanxy_out[17];
    assign wire_6276 = io_tile_0_3_chanxy_out[18];
    assign wire_6278 = io_tile_0_3_chanxy_out[19];
    assign wire_6280 = io_tile_0_3_chanxy_out[20];
    assign wire_6282 = io_tile_0_3_chanxy_out[21];
    assign wire_6284 = io_tile_0_3_chanxy_out[22];
    assign wire_6286 = io_tile_0_3_chanxy_out[23];
    assign wire_6288 = io_tile_0_3_chanxy_out[24];
    assign wire_6290 = io_tile_0_3_chanxy_out[25];
    assign wire_6292 = io_tile_0_3_chanxy_out[26];
    assign wire_6294 = io_tile_0_3_chanxy_out[27];
    assign wire_6296 = io_tile_0_3_chanxy_out[28];
    assign wire_6298 = io_tile_0_3_chanxy_out[29];
    assign io_tile_0_4_chanxy_in = {wire_11699, wire_11669, wire_11639, wire_11609, wire_6238, wire_2116, wire_2074, wire_2065, wire_2059, wire_11697, wire_11667, wire_11637, wire_11607, wire_6230, wire_2116, wire_2074, wire_2065, wire_2059, wire_11695, wire_11665, wire_11635, wire_11605, wire_6222, wire_2116, wire_2074, wire_2065, wire_2059, wire_11693, wire_11663, wire_11633, wire_11603, wire_6214, wire_2116, wire_2071, wire_2065, wire_2056, wire_11691, wire_11661, wire_11631, wire_11601, wire_6206, wire_2116, wire_2071, wire_2065, wire_2056, wire_11689, wire_11659, wire_11629, wire_11599, wire_6198, wire_2116, wire_2071, wire_2065, wire_2056, wire_11687, wire_11657, wire_11627, wire_11597, wire_6190, wire_2112, wire_2071, wire_2062, wire_2056, wire_11685, wire_11655, wire_11625, wire_11595, wire_6182, wire_2112, wire_2071, wire_2062, wire_2056, wire_11683, wire_11653, wire_11623, wire_11593, wire_6174, wire_2112, wire_2071, wire_2062, wire_2056, wire_11681, wire_11651, wire_11621, wire_11591, wire_6166, wire_2112, wire_2068, wire_2062, wire_2053, wire_11679, wire_11649, wire_11619, wire_11589, wire_6158, wire_2112, wire_2068, wire_2062, wire_2053, wire_11677, wire_11647, wire_11617, wire_11587, wire_6150, wire_2112, wire_2068, wire_2062, wire_2053, wire_11675, wire_11645, wire_11615, wire_11585, wire_6142, wire_2074, wire_2068, wire_2059, wire_2053, wire_11673, wire_11643, wire_11613, wire_11583, wire_6134, wire_2074, wire_2068, wire_2059, wire_2053, wire_11671, wire_11641, wire_11611, wire_11581, wire_6126, wire_2074, wire_2068, wire_2059, wire_2053, wire_12089, wire_12059, wire_12029, wire_11999, wire_6359, wire_2116, wire_2074, wire_2065, wire_2059, wire_12087, wire_12057, wire_12027, wire_11997, wire_6357, wire_2116, wire_2074, wire_2065, wire_2059, wire_12085, wire_12055, wire_12025, wire_11995, wire_6355, wire_2116, wire_2074, wire_2065, wire_2059, wire_12083, wire_12053, wire_12023, wire_11993, wire_6353, wire_2116, wire_2071, wire_2065, wire_2056, wire_12081, wire_12051, wire_12021, wire_11991, wire_6351, wire_2116, wire_2071, wire_2065, wire_2056, wire_12079, wire_12049, wire_12019, wire_11989, wire_6349, wire_2116, wire_2071, wire_2065, wire_2056, wire_12077, wire_12047, wire_12017, wire_11987, wire_6347, wire_2112, wire_2071, wire_2062, wire_2056, wire_12075, wire_12045, wire_12015, wire_11985, wire_6345, wire_2112, wire_2071, wire_2062, wire_2056, wire_12073, wire_12043, wire_12013, wire_11983, wire_6343, wire_2112, wire_2071, wire_2062, wire_2056, wire_12071, wire_12041, wire_12011, wire_11981, wire_6341, wire_2112, wire_2068, wire_2062, wire_2053, wire_12069, wire_12039, wire_12009, wire_11979, wire_6339, wire_2112, wire_2068, wire_2062, wire_2053, wire_12067, wire_12037, wire_12007, wire_11977, wire_6337, wire_2112, wire_2068, wire_2062, wire_2053, wire_12065, wire_12035, wire_12005, wire_11975, wire_6335, wire_2074, wire_2068, wire_2059, wire_2053, wire_12063, wire_12033, wire_12003, wire_11973, wire_6333, wire_2074, wire_2068, wire_2059, wire_2053, wire_12061, wire_12031, wire_12001, wire_11971, wire_6331, wire_2074, wire_2068, wire_2059, wire_2053};
    // CHNAXY TOTAL: 30
    assign wire_6121 = io_tile_0_4_chanxy_out[0];
    assign wire_6129 = io_tile_0_4_chanxy_out[1];
    assign wire_6137 = io_tile_0_4_chanxy_out[2];
    assign wire_6145 = io_tile_0_4_chanxy_out[3];
    assign wire_6153 = io_tile_0_4_chanxy_out[4];
    assign wire_6161 = io_tile_0_4_chanxy_out[5];
    assign wire_6169 = io_tile_0_4_chanxy_out[6];
    assign wire_6177 = io_tile_0_4_chanxy_out[7];
    assign wire_6185 = io_tile_0_4_chanxy_out[8];
    assign wire_6193 = io_tile_0_4_chanxy_out[9];
    assign wire_6201 = io_tile_0_4_chanxy_out[10];
    assign wire_6209 = io_tile_0_4_chanxy_out[11];
    assign wire_6217 = io_tile_0_4_chanxy_out[12];
    assign wire_6225 = io_tile_0_4_chanxy_out[13];
    assign wire_6233 = io_tile_0_4_chanxy_out[14];
    assign wire_6300 = io_tile_0_4_chanxy_out[15];
    assign wire_6302 = io_tile_0_4_chanxy_out[16];
    assign wire_6304 = io_tile_0_4_chanxy_out[17];
    assign wire_6306 = io_tile_0_4_chanxy_out[18];
    assign wire_6308 = io_tile_0_4_chanxy_out[19];
    assign wire_6310 = io_tile_0_4_chanxy_out[20];
    assign wire_6312 = io_tile_0_4_chanxy_out[21];
    assign wire_6314 = io_tile_0_4_chanxy_out[22];
    assign wire_6316 = io_tile_0_4_chanxy_out[23];
    assign wire_6318 = io_tile_0_4_chanxy_out[24];
    assign wire_6320 = io_tile_0_4_chanxy_out[25];
    assign wire_6322 = io_tile_0_4_chanxy_out[26];
    assign wire_6324 = io_tile_0_4_chanxy_out[27];
    assign wire_6326 = io_tile_0_4_chanxy_out[28];
    assign wire_6328 = io_tile_0_4_chanxy_out[29];
    assign io_tile_0_5_chanxy_in = {wire_12089, wire_12059, wire_12029, wire_11999, wire_6232, wire_2632, wire_2590, wire_2581, wire_2575, wire_12087, wire_12057, wire_12027, wire_11997, wire_6224, wire_2632, wire_2590, wire_2581, wire_2575, wire_12085, wire_12055, wire_12025, wire_11995, wire_6216, wire_2632, wire_2590, wire_2581, wire_2575, wire_12083, wire_12053, wire_12023, wire_11993, wire_6208, wire_2632, wire_2587, wire_2581, wire_2572, wire_12081, wire_12051, wire_12021, wire_11991, wire_6200, wire_2632, wire_2587, wire_2581, wire_2572, wire_12079, wire_12049, wire_12019, wire_11989, wire_6192, wire_2632, wire_2587, wire_2581, wire_2572, wire_12077, wire_12047, wire_12017, wire_11987, wire_6184, wire_2628, wire_2587, wire_2578, wire_2572, wire_12075, wire_12045, wire_12015, wire_11985, wire_6176, wire_2628, wire_2587, wire_2578, wire_2572, wire_12073, wire_12043, wire_12013, wire_11983, wire_6168, wire_2628, wire_2587, wire_2578, wire_2572, wire_12071, wire_12041, wire_12011, wire_11981, wire_6160, wire_2628, wire_2584, wire_2578, wire_2569, wire_12069, wire_12039, wire_12009, wire_11979, wire_6152, wire_2628, wire_2584, wire_2578, wire_2569, wire_12067, wire_12037, wire_12007, wire_11977, wire_6144, wire_2628, wire_2584, wire_2578, wire_2569, wire_12065, wire_12035, wire_12005, wire_11975, wire_6136, wire_2590, wire_2584, wire_2575, wire_2569, wire_12063, wire_12033, wire_12003, wire_11973, wire_6128, wire_2590, wire_2584, wire_2575, wire_2569, wire_12061, wire_12031, wire_12001, wire_11971, wire_6120, wire_2590, wire_2584, wire_2575, wire_2569, wire_12479, wire_12449, wire_12419, wire_12389, wire_6389, wire_2632, wire_2590, wire_2581, wire_2575, wire_12477, wire_12447, wire_12417, wire_12387, wire_6387, wire_2632, wire_2590, wire_2581, wire_2575, wire_12475, wire_12445, wire_12415, wire_12385, wire_6385, wire_2632, wire_2590, wire_2581, wire_2575, wire_12473, wire_12443, wire_12413, wire_12383, wire_6383, wire_2632, wire_2587, wire_2581, wire_2572, wire_12471, wire_12441, wire_12411, wire_12381, wire_6381, wire_2632, wire_2587, wire_2581, wire_2572, wire_12469, wire_12439, wire_12409, wire_12379, wire_6379, wire_2632, wire_2587, wire_2581, wire_2572, wire_12467, wire_12437, wire_12407, wire_12377, wire_6377, wire_2628, wire_2587, wire_2578, wire_2572, wire_12465, wire_12435, wire_12405, wire_12375, wire_6375, wire_2628, wire_2587, wire_2578, wire_2572, wire_12463, wire_12433, wire_12403, wire_12373, wire_6373, wire_2628, wire_2587, wire_2578, wire_2572, wire_12461, wire_12431, wire_12401, wire_12371, wire_6371, wire_2628, wire_2584, wire_2578, wire_2569, wire_12459, wire_12429, wire_12399, wire_12369, wire_6369, wire_2628, wire_2584, wire_2578, wire_2569, wire_12457, wire_12427, wire_12397, wire_12367, wire_6367, wire_2628, wire_2584, wire_2578, wire_2569, wire_12455, wire_12425, wire_12395, wire_12365, wire_6365, wire_2590, wire_2584, wire_2575, wire_2569, wire_12453, wire_12423, wire_12393, wire_12363, wire_6363, wire_2590, wire_2584, wire_2575, wire_2569, wire_12451, wire_12421, wire_12391, wire_12361, wire_6361, wire_2590, wire_2584, wire_2575, wire_2569};
    // CHNAXY TOTAL: 30
    assign wire_6241 = io_tile_0_5_chanxy_out[0];
    assign wire_6243 = io_tile_0_5_chanxy_out[1];
    assign wire_6245 = io_tile_0_5_chanxy_out[2];
    assign wire_6247 = io_tile_0_5_chanxy_out[3];
    assign wire_6249 = io_tile_0_5_chanxy_out[4];
    assign wire_6251 = io_tile_0_5_chanxy_out[5];
    assign wire_6253 = io_tile_0_5_chanxy_out[6];
    assign wire_6255 = io_tile_0_5_chanxy_out[7];
    assign wire_6257 = io_tile_0_5_chanxy_out[8];
    assign wire_6259 = io_tile_0_5_chanxy_out[9];
    assign wire_6261 = io_tile_0_5_chanxy_out[10];
    assign wire_6263 = io_tile_0_5_chanxy_out[11];
    assign wire_6265 = io_tile_0_5_chanxy_out[12];
    assign wire_6267 = io_tile_0_5_chanxy_out[13];
    assign wire_6269 = io_tile_0_5_chanxy_out[14];
    assign wire_6330 = io_tile_0_5_chanxy_out[15];
    assign wire_6332 = io_tile_0_5_chanxy_out[16];
    assign wire_6334 = io_tile_0_5_chanxy_out[17];
    assign wire_6336 = io_tile_0_5_chanxy_out[18];
    assign wire_6338 = io_tile_0_5_chanxy_out[19];
    assign wire_6340 = io_tile_0_5_chanxy_out[20];
    assign wire_6342 = io_tile_0_5_chanxy_out[21];
    assign wire_6344 = io_tile_0_5_chanxy_out[22];
    assign wire_6346 = io_tile_0_5_chanxy_out[23];
    assign wire_6348 = io_tile_0_5_chanxy_out[24];
    assign wire_6350 = io_tile_0_5_chanxy_out[25];
    assign wire_6352 = io_tile_0_5_chanxy_out[26];
    assign wire_6354 = io_tile_0_5_chanxy_out[27];
    assign wire_6356 = io_tile_0_5_chanxy_out[28];
    assign wire_6358 = io_tile_0_5_chanxy_out[29];
    assign io_tile_0_6_chanxy_in = {wire_12479, wire_12449, wire_12419, wire_12389, wire_6268, wire_3148, wire_3106, wire_3097, wire_3091, wire_12477, wire_12447, wire_12417, wire_12387, wire_6266, wire_3148, wire_3106, wire_3097, wire_3091, wire_12475, wire_12445, wire_12415, wire_12385, wire_6264, wire_3148, wire_3106, wire_3097, wire_3091, wire_12473, wire_12443, wire_12413, wire_12383, wire_6262, wire_3148, wire_3103, wire_3097, wire_3088, wire_12471, wire_12441, wire_12411, wire_12381, wire_6260, wire_3148, wire_3103, wire_3097, wire_3088, wire_12469, wire_12439, wire_12409, wire_12379, wire_6258, wire_3148, wire_3103, wire_3097, wire_3088, wire_12467, wire_12437, wire_12407, wire_12377, wire_6256, wire_3144, wire_3103, wire_3094, wire_3088, wire_12465, wire_12435, wire_12405, wire_12375, wire_6254, wire_3144, wire_3103, wire_3094, wire_3088, wire_12463, wire_12433, wire_12403, wire_12373, wire_6252, wire_3144, wire_3103, wire_3094, wire_3088, wire_12461, wire_12431, wire_12401, wire_12371, wire_6250, wire_3144, wire_3100, wire_3094, wire_3085, wire_12459, wire_12429, wire_12399, wire_12369, wire_6248, wire_3144, wire_3100, wire_3094, wire_3085, wire_12457, wire_12427, wire_12397, wire_12367, wire_6246, wire_3144, wire_3100, wire_3094, wire_3085, wire_12455, wire_12425, wire_12395, wire_12365, wire_6244, wire_3106, wire_3100, wire_3091, wire_3085, wire_12453, wire_12423, wire_12393, wire_12363, wire_6242, wire_3106, wire_3100, wire_3091, wire_3085, wire_12451, wire_12421, wire_12391, wire_12361, wire_6240, wire_3106, wire_3100, wire_3091, wire_3085, wire_12869, wire_12839, wire_12809, wire_12779, wire_6419, wire_3148, wire_3106, wire_3097, wire_3091, wire_12867, wire_12837, wire_12807, wire_12777, wire_6417, wire_3148, wire_3106, wire_3097, wire_3091, wire_12865, wire_12835, wire_12805, wire_12775, wire_6415, wire_3148, wire_3106, wire_3097, wire_3091, wire_12863, wire_12833, wire_12803, wire_12773, wire_6413, wire_3148, wire_3103, wire_3097, wire_3088, wire_12861, wire_12831, wire_12801, wire_12771, wire_6411, wire_3148, wire_3103, wire_3097, wire_3088, wire_12859, wire_12829, wire_12799, wire_12769, wire_6409, wire_3148, wire_3103, wire_3097, wire_3088, wire_12857, wire_12827, wire_12797, wire_12767, wire_6407, wire_3144, wire_3103, wire_3094, wire_3088, wire_12855, wire_12825, wire_12795, wire_12765, wire_6405, wire_3144, wire_3103, wire_3094, wire_3088, wire_12853, wire_12823, wire_12793, wire_12763, wire_6403, wire_3144, wire_3103, wire_3094, wire_3088, wire_12851, wire_12821, wire_12791, wire_12761, wire_6401, wire_3144, wire_3100, wire_3094, wire_3085, wire_12849, wire_12819, wire_12789, wire_12759, wire_6399, wire_3144, wire_3100, wire_3094, wire_3085, wire_12847, wire_12817, wire_12787, wire_12757, wire_6397, wire_3144, wire_3100, wire_3094, wire_3085, wire_12845, wire_12815, wire_12785, wire_12755, wire_6395, wire_3106, wire_3100, wire_3091, wire_3085, wire_12843, wire_12813, wire_12783, wire_12753, wire_6393, wire_3106, wire_3100, wire_3091, wire_3085, wire_12841, wire_12811, wire_12781, wire_12751, wire_6391, wire_3106, wire_3100, wire_3091, wire_3085};
    // CHNAXY TOTAL: 30
    assign wire_6271 = io_tile_0_6_chanxy_out[0];
    assign wire_6273 = io_tile_0_6_chanxy_out[1];
    assign wire_6275 = io_tile_0_6_chanxy_out[2];
    assign wire_6277 = io_tile_0_6_chanxy_out[3];
    assign wire_6279 = io_tile_0_6_chanxy_out[4];
    assign wire_6281 = io_tile_0_6_chanxy_out[5];
    assign wire_6283 = io_tile_0_6_chanxy_out[6];
    assign wire_6285 = io_tile_0_6_chanxy_out[7];
    assign wire_6287 = io_tile_0_6_chanxy_out[8];
    assign wire_6289 = io_tile_0_6_chanxy_out[9];
    assign wire_6291 = io_tile_0_6_chanxy_out[10];
    assign wire_6293 = io_tile_0_6_chanxy_out[11];
    assign wire_6295 = io_tile_0_6_chanxy_out[12];
    assign wire_6297 = io_tile_0_6_chanxy_out[13];
    assign wire_6299 = io_tile_0_6_chanxy_out[14];
    assign wire_6360 = io_tile_0_6_chanxy_out[15];
    assign wire_6362 = io_tile_0_6_chanxy_out[16];
    assign wire_6364 = io_tile_0_6_chanxy_out[17];
    assign wire_6366 = io_tile_0_6_chanxy_out[18];
    assign wire_6368 = io_tile_0_6_chanxy_out[19];
    assign wire_6370 = io_tile_0_6_chanxy_out[20];
    assign wire_6372 = io_tile_0_6_chanxy_out[21];
    assign wire_6374 = io_tile_0_6_chanxy_out[22];
    assign wire_6376 = io_tile_0_6_chanxy_out[23];
    assign wire_6378 = io_tile_0_6_chanxy_out[24];
    assign wire_6380 = io_tile_0_6_chanxy_out[25];
    assign wire_6382 = io_tile_0_6_chanxy_out[26];
    assign wire_6384 = io_tile_0_6_chanxy_out[27];
    assign wire_6386 = io_tile_0_6_chanxy_out[28];
    assign wire_6388 = io_tile_0_6_chanxy_out[29];
    assign io_tile_0_7_chanxy_in = {wire_12869, wire_12839, wire_12809, wire_12779, wire_6298, wire_3664, wire_3622, wire_3613, wire_3607, wire_12867, wire_12837, wire_12807, wire_12777, wire_6296, wire_3664, wire_3622, wire_3613, wire_3607, wire_12865, wire_12835, wire_12805, wire_12775, wire_6294, wire_3664, wire_3622, wire_3613, wire_3607, wire_12863, wire_12833, wire_12803, wire_12773, wire_6292, wire_3664, wire_3619, wire_3613, wire_3604, wire_12861, wire_12831, wire_12801, wire_12771, wire_6290, wire_3664, wire_3619, wire_3613, wire_3604, wire_12859, wire_12829, wire_12799, wire_12769, wire_6288, wire_3664, wire_3619, wire_3613, wire_3604, wire_12857, wire_12827, wire_12797, wire_12767, wire_6286, wire_3660, wire_3619, wire_3610, wire_3604, wire_12855, wire_12825, wire_12795, wire_12765, wire_6284, wire_3660, wire_3619, wire_3610, wire_3604, wire_12853, wire_12823, wire_12793, wire_12763, wire_6282, wire_3660, wire_3619, wire_3610, wire_3604, wire_12851, wire_12821, wire_12791, wire_12761, wire_6280, wire_3660, wire_3616, wire_3610, wire_3601, wire_12849, wire_12819, wire_12789, wire_12759, wire_6278, wire_3660, wire_3616, wire_3610, wire_3601, wire_12847, wire_12817, wire_12787, wire_12757, wire_6276, wire_3660, wire_3616, wire_3610, wire_3601, wire_12845, wire_12815, wire_12785, wire_12755, wire_6274, wire_3622, wire_3616, wire_3607, wire_3601, wire_12843, wire_12813, wire_12783, wire_12753, wire_6272, wire_3622, wire_3616, wire_3607, wire_3601, wire_12841, wire_12811, wire_12781, wire_12751, wire_6270, wire_3622, wire_3616, wire_3607, wire_3601, wire_13259, wire_13229, wire_13199, wire_13169, wire_6449, wire_3664, wire_3622, wire_3613, wire_3607, wire_13257, wire_13227, wire_13197, wire_13167, wire_6447, wire_3664, wire_3622, wire_3613, wire_3607, wire_13255, wire_13225, wire_13195, wire_13165, wire_6445, wire_3664, wire_3622, wire_3613, wire_3607, wire_13253, wire_13223, wire_13193, wire_13163, wire_6443, wire_3664, wire_3619, wire_3613, wire_3604, wire_13251, wire_13221, wire_13191, wire_13161, wire_6441, wire_3664, wire_3619, wire_3613, wire_3604, wire_13249, wire_13219, wire_13189, wire_13159, wire_6439, wire_3664, wire_3619, wire_3613, wire_3604, wire_13247, wire_13217, wire_13187, wire_13157, wire_6437, wire_3660, wire_3619, wire_3610, wire_3604, wire_13245, wire_13215, wire_13185, wire_13155, wire_6435, wire_3660, wire_3619, wire_3610, wire_3604, wire_13243, wire_13213, wire_13183, wire_13153, wire_6433, wire_3660, wire_3619, wire_3610, wire_3604, wire_13241, wire_13211, wire_13181, wire_13151, wire_6431, wire_3660, wire_3616, wire_3610, wire_3601, wire_13239, wire_13209, wire_13179, wire_13149, wire_6429, wire_3660, wire_3616, wire_3610, wire_3601, wire_13237, wire_13207, wire_13177, wire_13147, wire_6427, wire_3660, wire_3616, wire_3610, wire_3601, wire_13235, wire_13205, wire_13175, wire_13145, wire_6425, wire_3622, wire_3616, wire_3607, wire_3601, wire_13233, wire_13203, wire_13173, wire_13143, wire_6423, wire_3622, wire_3616, wire_3607, wire_3601, wire_13231, wire_13201, wire_13171, wire_13141, wire_6421, wire_3622, wire_3616, wire_3607, wire_3601};
    // CHNAXY TOTAL: 30
    assign wire_6301 = io_tile_0_7_chanxy_out[0];
    assign wire_6303 = io_tile_0_7_chanxy_out[1];
    assign wire_6305 = io_tile_0_7_chanxy_out[2];
    assign wire_6307 = io_tile_0_7_chanxy_out[3];
    assign wire_6309 = io_tile_0_7_chanxy_out[4];
    assign wire_6311 = io_tile_0_7_chanxy_out[5];
    assign wire_6313 = io_tile_0_7_chanxy_out[6];
    assign wire_6315 = io_tile_0_7_chanxy_out[7];
    assign wire_6317 = io_tile_0_7_chanxy_out[8];
    assign wire_6319 = io_tile_0_7_chanxy_out[9];
    assign wire_6321 = io_tile_0_7_chanxy_out[10];
    assign wire_6323 = io_tile_0_7_chanxy_out[11];
    assign wire_6325 = io_tile_0_7_chanxy_out[12];
    assign wire_6327 = io_tile_0_7_chanxy_out[13];
    assign wire_6329 = io_tile_0_7_chanxy_out[14];
    assign wire_6390 = io_tile_0_7_chanxy_out[15];
    assign wire_6392 = io_tile_0_7_chanxy_out[16];
    assign wire_6394 = io_tile_0_7_chanxy_out[17];
    assign wire_6396 = io_tile_0_7_chanxy_out[18];
    assign wire_6398 = io_tile_0_7_chanxy_out[19];
    assign wire_6400 = io_tile_0_7_chanxy_out[20];
    assign wire_6402 = io_tile_0_7_chanxy_out[21];
    assign wire_6404 = io_tile_0_7_chanxy_out[22];
    assign wire_6406 = io_tile_0_7_chanxy_out[23];
    assign wire_6408 = io_tile_0_7_chanxy_out[24];
    assign wire_6410 = io_tile_0_7_chanxy_out[25];
    assign wire_6412 = io_tile_0_7_chanxy_out[26];
    assign wire_6414 = io_tile_0_7_chanxy_out[27];
    assign wire_6416 = io_tile_0_7_chanxy_out[28];
    assign wire_6418 = io_tile_0_7_chanxy_out[29];
    assign io_tile_0_8_chanxy_in = {wire_13259, wire_13229, wire_13199, wire_13169, wire_6328, wire_4180, wire_4138, wire_4129, wire_4123, wire_13257, wire_13227, wire_13197, wire_13167, wire_6326, wire_4180, wire_4138, wire_4129, wire_4123, wire_13255, wire_13225, wire_13195, wire_13165, wire_6324, wire_4180, wire_4138, wire_4129, wire_4123, wire_13253, wire_13223, wire_13193, wire_13163, wire_6322, wire_4180, wire_4135, wire_4129, wire_4120, wire_13251, wire_13221, wire_13191, wire_13161, wire_6320, wire_4180, wire_4135, wire_4129, wire_4120, wire_13249, wire_13219, wire_13189, wire_13159, wire_6318, wire_4180, wire_4135, wire_4129, wire_4120, wire_13247, wire_13217, wire_13187, wire_13157, wire_6316, wire_4176, wire_4135, wire_4126, wire_4120, wire_13245, wire_13215, wire_13185, wire_13155, wire_6314, wire_4176, wire_4135, wire_4126, wire_4120, wire_13243, wire_13213, wire_13183, wire_13153, wire_6312, wire_4176, wire_4135, wire_4126, wire_4120, wire_13241, wire_13211, wire_13181, wire_13151, wire_6310, wire_4176, wire_4132, wire_4126, wire_4117, wire_13239, wire_13209, wire_13179, wire_13149, wire_6308, wire_4176, wire_4132, wire_4126, wire_4117, wire_13237, wire_13207, wire_13177, wire_13147, wire_6306, wire_4176, wire_4132, wire_4126, wire_4117, wire_13235, wire_13205, wire_13175, wire_13145, wire_6304, wire_4138, wire_4132, wire_4123, wire_4117, wire_13233, wire_13203, wire_13173, wire_13143, wire_6302, wire_4138, wire_4132, wire_4123, wire_4117, wire_13231, wire_13201, wire_13171, wire_13141, wire_6300, wire_4138, wire_4132, wire_4123, wire_4117, wire_13649, wire_13619, wire_13589, wire_13559, wire_6479, wire_4180, wire_4138, wire_4129, wire_4123, wire_13647, wire_13617, wire_13587, wire_13557, wire_6477, wire_4180, wire_4138, wire_4129, wire_4123, wire_13645, wire_13615, wire_13585, wire_13555, wire_6475, wire_4180, wire_4138, wire_4129, wire_4123, wire_13643, wire_13613, wire_13583, wire_13553, wire_6473, wire_4180, wire_4135, wire_4129, wire_4120, wire_13641, wire_13611, wire_13581, wire_13551, wire_6471, wire_4180, wire_4135, wire_4129, wire_4120, wire_13639, wire_13609, wire_13579, wire_13549, wire_6469, wire_4180, wire_4135, wire_4129, wire_4120, wire_13637, wire_13607, wire_13577, wire_13547, wire_6467, wire_4176, wire_4135, wire_4126, wire_4120, wire_13635, wire_13605, wire_13575, wire_13545, wire_6465, wire_4176, wire_4135, wire_4126, wire_4120, wire_13633, wire_13603, wire_13573, wire_13543, wire_6463, wire_4176, wire_4135, wire_4126, wire_4120, wire_13631, wire_13601, wire_13571, wire_13541, wire_6461, wire_4176, wire_4132, wire_4126, wire_4117, wire_13629, wire_13599, wire_13569, wire_13539, wire_6459, wire_4176, wire_4132, wire_4126, wire_4117, wire_13627, wire_13597, wire_13567, wire_13537, wire_6457, wire_4176, wire_4132, wire_4126, wire_4117, wire_13625, wire_13595, wire_13565, wire_13535, wire_6455, wire_4138, wire_4132, wire_4123, wire_4117, wire_13623, wire_13593, wire_13563, wire_13533, wire_6453, wire_4138, wire_4132, wire_4123, wire_4117, wire_13621, wire_13591, wire_13561, wire_13531, wire_6451, wire_4138, wire_4132, wire_4123, wire_4117};
    // CHNAXY TOTAL: 30
    assign wire_6331 = io_tile_0_8_chanxy_out[0];
    assign wire_6333 = io_tile_0_8_chanxy_out[1];
    assign wire_6335 = io_tile_0_8_chanxy_out[2];
    assign wire_6337 = io_tile_0_8_chanxy_out[3];
    assign wire_6339 = io_tile_0_8_chanxy_out[4];
    assign wire_6341 = io_tile_0_8_chanxy_out[5];
    assign wire_6343 = io_tile_0_8_chanxy_out[6];
    assign wire_6345 = io_tile_0_8_chanxy_out[7];
    assign wire_6347 = io_tile_0_8_chanxy_out[8];
    assign wire_6349 = io_tile_0_8_chanxy_out[9];
    assign wire_6351 = io_tile_0_8_chanxy_out[10];
    assign wire_6353 = io_tile_0_8_chanxy_out[11];
    assign wire_6355 = io_tile_0_8_chanxy_out[12];
    assign wire_6357 = io_tile_0_8_chanxy_out[13];
    assign wire_6359 = io_tile_0_8_chanxy_out[14];
    assign wire_6420 = io_tile_0_8_chanxy_out[15];
    assign wire_6422 = io_tile_0_8_chanxy_out[16];
    assign wire_6424 = io_tile_0_8_chanxy_out[17];
    assign wire_6426 = io_tile_0_8_chanxy_out[18];
    assign wire_6428 = io_tile_0_8_chanxy_out[19];
    assign wire_6430 = io_tile_0_8_chanxy_out[20];
    assign wire_6432 = io_tile_0_8_chanxy_out[21];
    assign wire_6434 = io_tile_0_8_chanxy_out[22];
    assign wire_6436 = io_tile_0_8_chanxy_out[23];
    assign wire_6438 = io_tile_0_8_chanxy_out[24];
    assign wire_6440 = io_tile_0_8_chanxy_out[25];
    assign wire_6442 = io_tile_0_8_chanxy_out[26];
    assign wire_6444 = io_tile_0_8_chanxy_out[27];
    assign wire_6446 = io_tile_0_8_chanxy_out[28];
    assign wire_6448 = io_tile_0_8_chanxy_out[29];
    assign io_tile_0_9_chanxy_in = {wire_13649, wire_13619, wire_13589, wire_13559, wire_6358, wire_4696, wire_4654, wire_4645, wire_4639, wire_13647, wire_13617, wire_13587, wire_13557, wire_6356, wire_4696, wire_4654, wire_4645, wire_4639, wire_13645, wire_13615, wire_13585, wire_13555, wire_6354, wire_4696, wire_4654, wire_4645, wire_4639, wire_13643, wire_13613, wire_13583, wire_13553, wire_6352, wire_4696, wire_4651, wire_4645, wire_4636, wire_13641, wire_13611, wire_13581, wire_13551, wire_6350, wire_4696, wire_4651, wire_4645, wire_4636, wire_13639, wire_13609, wire_13579, wire_13549, wire_6348, wire_4696, wire_4651, wire_4645, wire_4636, wire_13637, wire_13607, wire_13577, wire_13547, wire_6346, wire_4692, wire_4651, wire_4642, wire_4636, wire_13635, wire_13605, wire_13575, wire_13545, wire_6344, wire_4692, wire_4651, wire_4642, wire_4636, wire_13633, wire_13603, wire_13573, wire_13543, wire_6342, wire_4692, wire_4651, wire_4642, wire_4636, wire_13631, wire_13601, wire_13571, wire_13541, wire_6340, wire_4692, wire_4648, wire_4642, wire_4633, wire_13629, wire_13599, wire_13569, wire_13539, wire_6338, wire_4692, wire_4648, wire_4642, wire_4633, wire_13627, wire_13597, wire_13567, wire_13537, wire_6336, wire_4692, wire_4648, wire_4642, wire_4633, wire_13625, wire_13595, wire_13565, wire_13535, wire_6334, wire_4654, wire_4648, wire_4639, wire_4633, wire_13623, wire_13593, wire_13563, wire_13533, wire_6332, wire_4654, wire_4648, wire_4639, wire_4633, wire_13621, wire_13591, wire_13561, wire_13531, wire_6330, wire_4654, wire_4648, wire_4639, wire_4633, wire_14039, wire_14009, wire_13979, wire_13949, wire_6509, wire_4696, wire_4654, wire_4645, wire_4639, wire_14037, wire_14007, wire_13977, wire_13947, wire_6507, wire_4696, wire_4654, wire_4645, wire_4639, wire_14035, wire_14005, wire_13975, wire_13945, wire_6505, wire_4696, wire_4654, wire_4645, wire_4639, wire_14033, wire_14003, wire_13973, wire_13943, wire_6503, wire_4696, wire_4651, wire_4645, wire_4636, wire_14031, wire_14001, wire_13971, wire_13941, wire_6501, wire_4696, wire_4651, wire_4645, wire_4636, wire_14029, wire_13999, wire_13969, wire_13939, wire_6499, wire_4696, wire_4651, wire_4645, wire_4636, wire_14027, wire_13997, wire_13967, wire_13937, wire_6497, wire_4692, wire_4651, wire_4642, wire_4636, wire_14025, wire_13995, wire_13965, wire_13935, wire_6495, wire_4692, wire_4651, wire_4642, wire_4636, wire_14023, wire_13993, wire_13963, wire_13933, wire_6493, wire_4692, wire_4651, wire_4642, wire_4636, wire_14021, wire_13991, wire_13961, wire_13931, wire_6491, wire_4692, wire_4648, wire_4642, wire_4633, wire_14019, wire_13989, wire_13959, wire_13929, wire_6489, wire_4692, wire_4648, wire_4642, wire_4633, wire_14017, wire_13987, wire_13957, wire_13927, wire_6487, wire_4692, wire_4648, wire_4642, wire_4633, wire_14015, wire_13985, wire_13955, wire_13925, wire_6485, wire_4654, wire_4648, wire_4639, wire_4633, wire_14013, wire_13983, wire_13953, wire_13923, wire_6483, wire_4654, wire_4648, wire_4639, wire_4633, wire_14011, wire_13981, wire_13951, wire_13921, wire_6481, wire_4654, wire_4648, wire_4639, wire_4633};
    // CHNAXY TOTAL: 30
    assign wire_6361 = io_tile_0_9_chanxy_out[0];
    assign wire_6363 = io_tile_0_9_chanxy_out[1];
    assign wire_6365 = io_tile_0_9_chanxy_out[2];
    assign wire_6367 = io_tile_0_9_chanxy_out[3];
    assign wire_6369 = io_tile_0_9_chanxy_out[4];
    assign wire_6371 = io_tile_0_9_chanxy_out[5];
    assign wire_6373 = io_tile_0_9_chanxy_out[6];
    assign wire_6375 = io_tile_0_9_chanxy_out[7];
    assign wire_6377 = io_tile_0_9_chanxy_out[8];
    assign wire_6379 = io_tile_0_9_chanxy_out[9];
    assign wire_6381 = io_tile_0_9_chanxy_out[10];
    assign wire_6383 = io_tile_0_9_chanxy_out[11];
    assign wire_6385 = io_tile_0_9_chanxy_out[12];
    assign wire_6387 = io_tile_0_9_chanxy_out[13];
    assign wire_6389 = io_tile_0_9_chanxy_out[14];
    assign wire_6450 = io_tile_0_9_chanxy_out[15];
    assign wire_6452 = io_tile_0_9_chanxy_out[16];
    assign wire_6454 = io_tile_0_9_chanxy_out[17];
    assign wire_6456 = io_tile_0_9_chanxy_out[18];
    assign wire_6458 = io_tile_0_9_chanxy_out[19];
    assign wire_6460 = io_tile_0_9_chanxy_out[20];
    assign wire_6462 = io_tile_0_9_chanxy_out[21];
    assign wire_6464 = io_tile_0_9_chanxy_out[22];
    assign wire_6466 = io_tile_0_9_chanxy_out[23];
    assign wire_6468 = io_tile_0_9_chanxy_out[24];
    assign wire_6470 = io_tile_0_9_chanxy_out[25];
    assign wire_6472 = io_tile_0_9_chanxy_out[26];
    assign wire_6474 = io_tile_0_9_chanxy_out[27];
    assign wire_6476 = io_tile_0_9_chanxy_out[28];
    assign wire_6478 = io_tile_0_9_chanxy_out[29];
    assign io_tile_0_10_chanxy_in = {wire_14317, wire_5212, wire_14039, wire_14009, wire_13979, wire_13949, wire_6388, wire_5212, wire_5170, wire_5161, wire_5155, wire_14325, wire_5208, wire_14037, wire_14007, wire_13977, wire_13947, wire_6386, wire_5212, wire_5170, wire_5161, wire_5155, wire_14333, wire_5208, wire_14035, wire_14005, wire_13975, wire_13945, wire_6384, wire_5212, wire_5170, wire_5161, wire_5155, wire_14341, wire_5170, wire_14033, wire_14003, wire_13973, wire_13943, wire_6382, wire_5212, wire_5167, wire_5161, wire_5152, wire_14349, wire_5167, wire_14031, wire_14001, wire_13971, wire_13941, wire_6380, wire_5212, wire_5167, wire_5161, wire_5152, wire_14357, wire_5167, wire_14029, wire_13999, wire_13969, wire_13939, wire_6378, wire_5212, wire_5167, wire_5161, wire_5152, wire_14365, wire_5164, wire_14027, wire_13997, wire_13967, wire_13937, wire_6376, wire_5208, wire_5167, wire_5158, wire_5152, wire_14373, wire_5161, wire_14025, wire_13995, wire_13965, wire_13935, wire_6374, wire_5208, wire_5167, wire_5158, wire_5152, wire_14381, wire_5161, wire_14023, wire_13993, wire_13963, wire_13933, wire_6372, wire_5208, wire_5167, wire_5158, wire_5152, wire_14389, wire_5158, wire_14021, wire_13991, wire_13961, wire_13931, wire_6370, wire_5208, wire_5164, wire_5158, wire_5149, wire_14397, wire_5155, wire_14019, wire_13989, wire_13959, wire_13929, wire_6368, wire_5208, wire_5164, wire_5158, wire_5149, wire_14405, wire_5155, wire_14017, wire_13987, wire_13957, wire_13927, wire_6366, wire_5208, wire_5164, wire_5158, wire_5149, wire_14413, wire_5152, wire_14015, wire_13985, wire_13955, wire_13925, wire_6364, wire_5170, wire_5164, wire_5155, wire_5149, wire_14421, wire_5149, wire_14013, wire_13983, wire_13953, wire_13923, wire_6362, wire_5170, wire_5164, wire_5155, wire_5149, wire_14429, wire_5149, wire_14011, wire_13981, wire_13951, wire_13921, wire_6360, wire_5170, wire_5164, wire_5155, wire_5149, wire_14319, wire_5212, wire_14327, wire_5208, wire_14335, wire_5208, wire_14343, wire_5170, wire_14351, wire_5167, wire_14359, wire_5167, wire_14367, wire_5164, wire_14375, wire_5161, wire_14383, wire_5161, wire_14391, wire_5158, wire_14399, wire_5155, wire_14407, wire_5155, wire_14415, wire_5152, wire_14423, wire_5149, wire_14311, wire_5149, wire_14313, wire_5212, wire_14321, wire_5212, wire_14329, wire_5208, wire_14337, wire_5170, wire_14345, wire_5170, wire_14353, wire_5167, wire_14361, wire_5164, wire_14369, wire_5164, wire_14377, wire_5161, wire_14385, wire_5158, wire_14393, wire_5158, wire_14401, wire_5155, wire_14409, wire_5152, wire_14417, wire_5152, wire_14425, wire_5149, wire_14315, wire_5212, wire_14323, wire_5212, wire_14331, wire_5208, wire_14339, wire_5170, wire_14347, wire_5170, wire_14355, wire_5167, wire_14363, wire_5164, wire_14371, wire_5164, wire_14379, wire_5161, wire_14387, wire_5158, wire_14395, wire_5158, wire_14403, wire_5155, wire_14411, wire_5152, wire_14419, wire_5152, wire_14427, wire_5149};
    // CHNAXY TOTAL: 75
    assign wire_6391 = io_tile_0_10_chanxy_out[0];
    assign wire_6393 = io_tile_0_10_chanxy_out[1];
    assign wire_6395 = io_tile_0_10_chanxy_out[2];
    assign wire_6397 = io_tile_0_10_chanxy_out[3];
    assign wire_6399 = io_tile_0_10_chanxy_out[4];
    assign wire_6401 = io_tile_0_10_chanxy_out[5];
    assign wire_6403 = io_tile_0_10_chanxy_out[6];
    assign wire_6405 = io_tile_0_10_chanxy_out[7];
    assign wire_6407 = io_tile_0_10_chanxy_out[8];
    assign wire_6409 = io_tile_0_10_chanxy_out[9];
    assign wire_6411 = io_tile_0_10_chanxy_out[10];
    assign wire_6413 = io_tile_0_10_chanxy_out[11];
    assign wire_6415 = io_tile_0_10_chanxy_out[12];
    assign wire_6417 = io_tile_0_10_chanxy_out[13];
    assign wire_6419 = io_tile_0_10_chanxy_out[14];
    assign wire_6421 = io_tile_0_10_chanxy_out[15];
    assign wire_6423 = io_tile_0_10_chanxy_out[16];
    assign wire_6425 = io_tile_0_10_chanxy_out[17];
    assign wire_6427 = io_tile_0_10_chanxy_out[18];
    assign wire_6429 = io_tile_0_10_chanxy_out[19];
    assign wire_6431 = io_tile_0_10_chanxy_out[20];
    assign wire_6433 = io_tile_0_10_chanxy_out[21];
    assign wire_6435 = io_tile_0_10_chanxy_out[22];
    assign wire_6437 = io_tile_0_10_chanxy_out[23];
    assign wire_6439 = io_tile_0_10_chanxy_out[24];
    assign wire_6441 = io_tile_0_10_chanxy_out[25];
    assign wire_6443 = io_tile_0_10_chanxy_out[26];
    assign wire_6445 = io_tile_0_10_chanxy_out[27];
    assign wire_6447 = io_tile_0_10_chanxy_out[28];
    assign wire_6449 = io_tile_0_10_chanxy_out[29];
    assign wire_6451 = io_tile_0_10_chanxy_out[30];
    assign wire_6453 = io_tile_0_10_chanxy_out[31];
    assign wire_6455 = io_tile_0_10_chanxy_out[32];
    assign wire_6457 = io_tile_0_10_chanxy_out[33];
    assign wire_6459 = io_tile_0_10_chanxy_out[34];
    assign wire_6461 = io_tile_0_10_chanxy_out[35];
    assign wire_6463 = io_tile_0_10_chanxy_out[36];
    assign wire_6465 = io_tile_0_10_chanxy_out[37];
    assign wire_6467 = io_tile_0_10_chanxy_out[38];
    assign wire_6469 = io_tile_0_10_chanxy_out[39];
    assign wire_6471 = io_tile_0_10_chanxy_out[40];
    assign wire_6473 = io_tile_0_10_chanxy_out[41];
    assign wire_6475 = io_tile_0_10_chanxy_out[42];
    assign wire_6477 = io_tile_0_10_chanxy_out[43];
    assign wire_6479 = io_tile_0_10_chanxy_out[44];
    assign wire_6480 = io_tile_0_10_chanxy_out[45];
    assign wire_6481 = io_tile_0_10_chanxy_out[46];
    assign wire_6482 = io_tile_0_10_chanxy_out[47];
    assign wire_6483 = io_tile_0_10_chanxy_out[48];
    assign wire_6484 = io_tile_0_10_chanxy_out[49];
    assign wire_6485 = io_tile_0_10_chanxy_out[50];
    assign wire_6486 = io_tile_0_10_chanxy_out[51];
    assign wire_6487 = io_tile_0_10_chanxy_out[52];
    assign wire_6488 = io_tile_0_10_chanxy_out[53];
    assign wire_6489 = io_tile_0_10_chanxy_out[54];
    assign wire_6490 = io_tile_0_10_chanxy_out[55];
    assign wire_6491 = io_tile_0_10_chanxy_out[56];
    assign wire_6492 = io_tile_0_10_chanxy_out[57];
    assign wire_6493 = io_tile_0_10_chanxy_out[58];
    assign wire_6494 = io_tile_0_10_chanxy_out[59];
    assign wire_6495 = io_tile_0_10_chanxy_out[60];
    assign wire_6496 = io_tile_0_10_chanxy_out[61];
    assign wire_6497 = io_tile_0_10_chanxy_out[62];
    assign wire_6498 = io_tile_0_10_chanxy_out[63];
    assign wire_6499 = io_tile_0_10_chanxy_out[64];
    assign wire_6500 = io_tile_0_10_chanxy_out[65];
    assign wire_6501 = io_tile_0_10_chanxy_out[66];
    assign wire_6502 = io_tile_0_10_chanxy_out[67];
    assign wire_6503 = io_tile_0_10_chanxy_out[68];
    assign wire_6504 = io_tile_0_10_chanxy_out[69];
    assign wire_6505 = io_tile_0_10_chanxy_out[70];
    assign wire_6506 = io_tile_0_10_chanxy_out[71];
    assign wire_6507 = io_tile_0_10_chanxy_out[72];
    assign wire_6508 = io_tile_0_10_chanxy_out[73];
    assign wire_6509 = io_tile_0_10_chanxy_out[74];
endmodule
