module io_sbcb_wc(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [339:0] io_chanxy_in,
    input [159:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[99:0] io_chanxy_out);

  wire[99:0] T0;
  wire[99:0] T1;
  wire[98:0] T2;
  wire[98:0] T3;
  wire[97:0] T4;
  wire[97:0] T5;
  wire[96:0] T6;
  wire[96:0] T7;
  wire[95:0] T8;
  wire[95:0] T9;
  wire[94:0] T10;
  wire[94:0] T11;
  wire[93:0] T12;
  wire[93:0] T13;
  wire[92:0] T14;
  wire[92:0] T15;
  wire[91:0] T16;
  wire[91:0] T17;
  wire[90:0] T18;
  wire[90:0] T19;
  wire[89:0] T20;
  wire[89:0] T21;
  wire[88:0] T22;
  wire[88:0] T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[86:0] T26;
  wire[86:0] T27;
  wire[85:0] T28;
  wire[85:0] T29;
  wire[84:0] T30;
  wire[84:0] T31;
  wire[83:0] T32;
  wire[83:0] T33;
  wire[82:0] T34;
  wire[82:0] T35;
  wire[81:0] T36;
  wire[81:0] T37;
  wire[80:0] T38;
  wire[80:0] T39;
  wire[79:0] T40;
  wire[79:0] T41;
  wire[78:0] T42;
  wire[78:0] T43;
  wire[77:0] T44;
  wire[77:0] T45;
  wire[76:0] T46;
  wire[76:0] T47;
  wire[75:0] T48;
  wire[75:0] T49;
  wire[74:0] T50;
  wire[74:0] T51;
  wire[73:0] T52;
  wire[73:0] T53;
  wire[72:0] T54;
  wire[72:0] T55;
  wire[71:0] T56;
  wire[71:0] T57;
  wire[70:0] T58;
  wire[70:0] T59;
  wire[69:0] T60;
  wire[69:0] T61;
  wire[68:0] T62;
  wire[68:0] T63;
  wire[67:0] T64;
  wire[67:0] T65;
  wire[66:0] T66;
  wire[66:0] T67;
  wire[65:0] T68;
  wire[65:0] T69;
  wire[64:0] T70;
  wire[64:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[62:0] T74;
  wire[62:0] T75;
  wire[61:0] T76;
  wire[61:0] T77;
  wire[60:0] T78;
  wire[60:0] T79;
  wire[59:0] T80;
  wire[59:0] T81;
  wire[58:0] T82;
  wire[58:0] T83;
  wire[57:0] T84;
  wire[57:0] T85;
  wire[56:0] T86;
  wire[56:0] T87;
  wire[55:0] T88;
  wire[55:0] T89;
  wire[54:0] T90;
  wire[54:0] T91;
  wire[53:0] T92;
  wire[53:0] T93;
  wire[52:0] T94;
  wire[52:0] T95;
  wire[51:0] T96;
  wire[51:0] T97;
  wire[50:0] T98;
  wire[50:0] T99;
  wire[49:0] T100;
  wire[49:0] T101;
  wire[48:0] T102;
  wire[48:0] T103;
  wire[47:0] T104;
  wire[47:0] T105;
  wire[46:0] T106;
  wire[46:0] T107;
  wire[45:0] T108;
  wire[45:0] T109;
  wire[44:0] T110;
  wire[44:0] T111;
  wire[43:0] T112;
  wire[43:0] T113;
  wire[42:0] T114;
  wire[42:0] T115;
  wire[41:0] T116;
  wire[41:0] T117;
  wire[40:0] T118;
  wire[40:0] T119;
  wire[39:0] T120;
  wire[39:0] T121;
  wire[38:0] T122;
  wire[38:0] T123;
  wire[37:0] T124;
  wire[37:0] T125;
  wire[36:0] T126;
  wire[36:0] T127;
  wire[35:0] T128;
  wire[35:0] T129;
  wire[34:0] T130;
  wire[34:0] T131;
  wire[33:0] T132;
  wire[33:0] T133;
  wire[32:0] T134;
  wire[32:0] T135;
  wire[31:0] T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire[30:0] T139;
  wire[29:0] T140;
  wire[29:0] T141;
  wire[28:0] T142;
  wire[28:0] T143;
  wire[27:0] T144;
  wire[27:0] T145;
  wire[26:0] T146;
  wire[26:0] T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire[24:0] T150;
  wire[24:0] T151;
  wire[23:0] T152;
  wire[23:0] T153;
  wire[22:0] T154;
  wire[22:0] T155;
  wire[21:0] T156;
  wire[21:0] T157;
  wire[20:0] T158;
  wire[20:0] T159;
  wire[19:0] T160;
  wire[19:0] T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[17:0] T164;
  wire[17:0] T165;
  wire[16:0] T166;
  wire[16:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire[14:0] T170;
  wire[14:0] T171;
  wire[13:0] T172;
  wire[13:0] T173;
  wire[12:0] T174;
  wire[12:0] T175;
  wire[11:0] T176;
  wire[11:0] T177;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[9:0] T180;
  wire[9:0] T181;
  wire[8:0] T182;
  wire[8:0] T183;
  wire[7:0] T184;
  wire[7:0] T185;
  wire[6:0] T186;
  wire[6:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] T219;
  wire[8:0] T220;
  wire[8:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[8:0] T260;
  wire[8:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[8:0] T300;
  wire[8:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[8:0] T340;
  wire[8:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[8:0] T380;
  wire[8:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[8:0] T420;
  wire[8:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[8:0] T460;
  wire[8:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[8:0] T500;
  wire[8:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[8:0] T540;
  wire[8:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[8:0] T580;
  wire[8:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[3:0] T617;
  wire[3:0] T618;
  wire[3:0] T619;
  wire[8:0] T620;
  wire[8:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[3:0] T657;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[8:0] T660;
  wire[8:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[8:0] T700;
  wire[8:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[3:0] T737;
  wire[3:0] T738;
  wire[3:0] T739;
  wire[8:0] T740;
  wire[8:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[8:0] T780;
  wire[8:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[3:0] T817;
  wire[3:0] T818;
  wire[3:0] T819;
  wire[8:0] T820;
  wire[8:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[8:0] T860;
  wire[8:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[8:0] T900;
  wire[8:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[8:0] T940;
  wire[8:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[8:0] T980;
  wire[8:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire[7:0] T998;
  wire[7:0] T999;
  wire[6:0] T1000;
  wire[6:0] T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[4:0] T1004;
  wire[4:0] T1005;
  wire[3:0] T1006;
  wire[3:0] T1007;
  wire[2:0] T1008;
  wire[2:0] T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire[15:0] T1015;
  wire[15:0] T1016;
  wire[15:0] T1017;
  wire[3:0] T1018;
  wire[15:0] T1019;
  wire[15:0] T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[15:0] T1024;
  wire[15:0] T1025;
  wire[15:0] T1026;
  wire[3:0] T1027;
  wire[15:0] T1028;
  wire[15:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[15:0] T1033;
  wire[15:0] T1034;
  wire[15:0] T1035;
  wire[3:0] T1036;
  wire[15:0] T1037;
  wire[15:0] T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire[15:0] T1042;
  wire[15:0] T1043;
  wire[15:0] T1044;
  wire[3:0] T1045;
  wire[15:0] T1046;
  wire[15:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire[15:0] T1051;
  wire[15:0] T1052;
  wire[15:0] T1053;
  wire[3:0] T1054;
  wire[15:0] T1055;
  wire[15:0] T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[15:0] T1060;
  wire[15:0] T1061;
  wire[15:0] T1062;
  wire[3:0] T1063;
  wire[15:0] T1064;
  wire[15:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[15:0] T1069;
  wire[15:0] T1070;
  wire[15:0] T1071;
  wire[3:0] T1072;
  wire[15:0] T1073;
  wire[15:0] T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire[15:0] T1078;
  wire[15:0] T1079;
  wire[15:0] T1080;
  wire[3:0] T1081;
  wire[15:0] T1082;
  wire[15:0] T1083;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T990, T2};
  assign T2 = T3;
  assign T3 = {T982, T4};
  assign T4 = T5;
  assign T5 = {T974, T6};
  assign T6 = T7;
  assign T7 = {T966, T8};
  assign T8 = T9;
  assign T9 = {T958, T10};
  assign T10 = T11;
  assign T11 = {T950, T12};
  assign T12 = T13;
  assign T13 = {T942, T14};
  assign T14 = T15;
  assign T15 = {T934, T16};
  assign T16 = T17;
  assign T17 = {T926, T18};
  assign T18 = T19;
  assign T19 = {T918, T20};
  assign T20 = T21;
  assign T21 = {T910, T22};
  assign T22 = T23;
  assign T23 = {T902, T24};
  assign T24 = T25;
  assign T25 = {T894, T26};
  assign T26 = T27;
  assign T27 = {T886, T28};
  assign T28 = T29;
  assign T29 = {T878, T30};
  assign T30 = T31;
  assign T31 = {T870, T32};
  assign T32 = T33;
  assign T33 = {T862, T34};
  assign T34 = T35;
  assign T35 = {T854, T36};
  assign T36 = T37;
  assign T37 = {T846, T38};
  assign T38 = T39;
  assign T39 = {T838, T40};
  assign T40 = T41;
  assign T41 = {T830, T42};
  assign T42 = T43;
  assign T43 = {T822, T44};
  assign T44 = T45;
  assign T45 = {T814, T46};
  assign T46 = T47;
  assign T47 = {T806, T48};
  assign T48 = T49;
  assign T49 = {T798, T50};
  assign T50 = T51;
  assign T51 = {T790, T52};
  assign T52 = T53;
  assign T53 = {T782, T54};
  assign T54 = T55;
  assign T55 = {T774, T56};
  assign T56 = T57;
  assign T57 = {T766, T58};
  assign T58 = T59;
  assign T59 = {T758, T60};
  assign T60 = T61;
  assign T61 = {T750, T62};
  assign T62 = T63;
  assign T63 = {T742, T64};
  assign T64 = T65;
  assign T65 = {T734, T66};
  assign T66 = T67;
  assign T67 = {T726, T68};
  assign T68 = T69;
  assign T69 = {T718, T70};
  assign T70 = T71;
  assign T71 = {T710, T72};
  assign T72 = T73;
  assign T73 = {T702, T74};
  assign T74 = T75;
  assign T75 = {T694, T76};
  assign T76 = T77;
  assign T77 = {T686, T78};
  assign T78 = T79;
  assign T79 = {T678, T80};
  assign T80 = T81;
  assign T81 = {T670, T82};
  assign T82 = T83;
  assign T83 = {T662, T84};
  assign T84 = T85;
  assign T85 = {T654, T86};
  assign T86 = T87;
  assign T87 = {T646, T88};
  assign T88 = T89;
  assign T89 = {T638, T90};
  assign T90 = T91;
  assign T91 = {T630, T92};
  assign T92 = T93;
  assign T93 = {T622, T94};
  assign T94 = T95;
  assign T95 = {T614, T96};
  assign T96 = T97;
  assign T97 = {T606, T98};
  assign T98 = T99;
  assign T99 = {T598, T100};
  assign T100 = T101;
  assign T101 = {T590, T102};
  assign T102 = T103;
  assign T103 = {T582, T104};
  assign T104 = T105;
  assign T105 = {T574, T106};
  assign T106 = T107;
  assign T107 = {T566, T108};
  assign T108 = T109;
  assign T109 = {T558, T110};
  assign T110 = T111;
  assign T111 = {T550, T112};
  assign T112 = T113;
  assign T113 = {T542, T114};
  assign T114 = T115;
  assign T115 = {T534, T116};
  assign T116 = T117;
  assign T117 = {T526, T118};
  assign T118 = T119;
  assign T119 = {T518, T120};
  assign T120 = T121;
  assign T121 = {T510, T122};
  assign T122 = T123;
  assign T123 = {T502, T124};
  assign T124 = T125;
  assign T125 = {T494, T126};
  assign T126 = T127;
  assign T127 = {T486, T128};
  assign T128 = T129;
  assign T129 = {T478, T130};
  assign T130 = T131;
  assign T131 = {T470, T132};
  assign T132 = T133;
  assign T133 = {T462, T134};
  assign T134 = T135;
  assign T135 = {T454, T136};
  assign T136 = T137;
  assign T137 = {T446, T138};
  assign T138 = T139;
  assign T139 = {T438, T140};
  assign T140 = T141;
  assign T141 = {T430, T142};
  assign T142 = T143;
  assign T143 = {T422, T144};
  assign T144 = T145;
  assign T145 = {T414, T146};
  assign T146 = T147;
  assign T147 = {T406, T148};
  assign T148 = T149;
  assign T149 = {T398, T150};
  assign T150 = T151;
  assign T151 = {T390, T152};
  assign T152 = T153;
  assign T153 = {T382, T154};
  assign T154 = T155;
  assign T155 = {T374, T156};
  assign T156 = T157;
  assign T157 = {T366, T158};
  assign T158 = T159;
  assign T159 = {T358, T160};
  assign T160 = T161;
  assign T161 = {T350, T162};
  assign T162 = T163;
  assign T163 = {T342, T164};
  assign T164 = T165;
  assign T165 = {T334, T166};
  assign T166 = T167;
  assign T167 = {T326, T168};
  assign T168 = T169;
  assign T169 = {T318, T170};
  assign T170 = T171;
  assign T171 = {T310, T172};
  assign T172 = T173;
  assign T173 = {T302, T174};
  assign T174 = T175;
  assign T175 = {T294, T176};
  assign T176 = T177;
  assign T177 = {T286, T178};
  assign T178 = T179;
  assign T179 = {T278, T180};
  assign T180 = T181;
  assign T181 = {T270, T182};
  assign T182 = T183;
  assign T183 = {T262, T184};
  assign T184 = T185;
  assign T185 = {T254, T186};
  assign T186 = T187;
  assign T187 = {T246, T188};
  assign T188 = T189;
  assign T189 = {T238, T190};
  assign T190 = T191;
  assign T191 = {T230, T192};
  assign T192 = T193;
  assign T193 = {T222, T194};
  assign T194 = T195;
  assign T195 = {T214, T196};
  assign T196 = T197;
  assign T197 = {T206, T198};
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[3'h5/* 5*/:2'h2/* 2*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[4'hc/* 12*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[3'h6/* 6*/:3'h6/* 6*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[4'he/* 14*/:4'hd/* 13*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[5'h10/* 16*/:4'hf/* 15*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[5'h12/* 18*/:5'h11/* 17*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[5'h14/* 20*/:5'h13/* 19*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[4'hd/* 13*/:4'ha/* 10*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[5'h1d/* 29*/:5'h15/* 21*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[5'h15/* 21*/:5'h12/* 18*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[6'h2e/* 46*/:6'h26/* 38*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h30/* 48*/:6'h2f/* 47*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h32/* 50*/:6'h31/* 49*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[6'h34/* 52*/:6'h33/* 51*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[6'h36/* 54*/:6'h35/* 53*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h1d/* 29*/:5'h1a/* 26*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[6'h3f/* 63*/:6'h37/* 55*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h25/* 37*/:6'h22/* 34*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[7'h50/* 80*/:7'h48/* 72*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[7'h52/* 82*/:7'h51/* 81*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[7'h54/* 84*/:7'h53/* 83*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[7'h56/* 86*/:7'h55/* 85*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[7'h58/* 88*/:7'h57/* 87*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[6'h2d/* 45*/:6'h2a/* 42*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[7'h61/* 97*/:7'h59/* 89*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h2e/* 46*/:6'h2e/* 46*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h2f/* 47*/:6'h2f/* 47*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h35/* 53*/:6'h32/* 50*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h72/* 114*/:7'h6a/* 106*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h74/* 116*/:7'h73/* 115*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h76/* 118*/:7'h75/* 117*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h78/* 120*/:7'h77/* 119*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h7a/* 122*/:7'h79/* 121*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[6'h3d/* 61*/:6'h3a/* 58*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[8'h83/* 131*/:7'h7b/* 123*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[6'h3e/* 62*/:6'h3e/* 62*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[8'h85/* 133*/:8'h84/* 132*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[6'h3f/* 63*/:6'h3f/* 63*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[8'h87/* 135*/:8'h86/* 134*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h41/* 65*/:7'h41/* 65*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[8'h94/* 148*/:8'h8c/* 140*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[7'h46/* 70*/:7'h46/* 70*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[8'h96/* 150*/:8'h95/* 149*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[7'h47/* 71*/:7'h47/* 71*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[8'h98/* 152*/:8'h97/* 151*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[8'h9a/* 154*/:8'h99/* 153*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[7'h4d/* 77*/:7'h4a/* 74*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[8'ha5/* 165*/:8'h9d/* 157*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[7'h4e/* 78*/:7'h4e/* 78*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[8'hab/* 171*/:8'haa/* 170*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[8'had/* 173*/:8'hac/* 172*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h55/* 85*/:7'h52/* 82*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[8'hb6/* 182*/:8'hae/* 174*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'hb8/* 184*/:8'hb7/* 183*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'hba/* 186*/:8'hb9/* 185*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'hbe/* 190*/:8'hbd/* 189*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'hc7/* 199*/:8'hbf/* 191*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'hcb/* 203*/:8'hca/* 202*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'hcf/* 207*/:8'hce/* 206*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h65/* 101*/:7'h62/* 98*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'hd8/* 216*/:8'hd0/* 208*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h66/* 102*/:7'h66/* 102*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hdc/* 220*/:8'hdb/* 219*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hde/* 222*/:8'hdd/* 221*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'he0/* 224*/:8'hdf/* 223*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h6d/* 109*/:7'h6a/* 106*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'he9/* 233*/:8'he1/* 225*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h6e/* 110*/:7'h6e/* 110*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'heb/* 235*/:8'hea/* 234*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'hed/* 237*/:8'hec/* 236*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'hef/* 239*/:8'hee/* 238*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'hfa/* 250*/:8'hf2/* 242*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h102/* 258*/:9'h101/* 257*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h7d/* 125*/:7'h7a/* 122*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h10b/* 267*/:9'h103/* 259*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h113/* 275*/:9'h112/* 274*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h11c/* 284*/:9'h114/* 276*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h12d/* 301*/:9'h125/* 293*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h135/* 309*/:9'h134/* 308*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h95/* 149*/:8'h92/* 146*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h13e/* 318*/:9'h136/* 310*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h96/* 150*/:8'h96/* 150*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h140/* 320*/:9'h13f/* 319*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'h9d/* 157*/:8'h9a/* 154*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h14f/* 335*/:9'h147/* 327*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h151/* 337*/:9'h150/* 336*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign io_ipin_out = T998;
  assign T998 = T999;
  assign T999 = {T1075, T1000};
  assign T1000 = T1001;
  assign T1001 = {T1066, T1002};
  assign T1002 = T1003;
  assign T1003 = {T1057, T1004};
  assign T1004 = T1005;
  assign T1005 = {T1048, T1006};
  assign T1006 = T1007;
  assign T1007 = {T1039, T1008};
  assign T1008 = T1009;
  assign T1009 = {T1030, T1010};
  assign T1010 = T1011;
  assign T1011 = {T1021, T1012};
  assign T1012 = T1013;
  assign T1013 = T1014;
  assign T1014 = T1019[T1015];
  assign T1015 = T1016;
  assign T1016 = T1017;
  assign T1017 = {12'h0/* 0*/, T1018};
  assign T1018 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1019 = T1020;
  assign T1020 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = T1028[T1024];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = {12'h0/* 0*/, T1027};
  assign T1027 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1028 = T1029;
  assign T1029 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1037[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = {12'h0/* 0*/, T1036};
  assign T1036 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1037 = T1038;
  assign T1038 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1039 = T1040;
  assign T1040 = T1041;
  assign T1041 = T1046[T1042];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = {12'h0/* 0*/, T1045};
  assign T1045 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1046 = T1047;
  assign T1047 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1048 = T1049;
  assign T1049 = T1050;
  assign T1050 = T1055[T1051];
  assign T1051 = T1052;
  assign T1052 = T1053;
  assign T1053 = {12'h0/* 0*/, T1054};
  assign T1054 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1055 = T1056;
  assign T1056 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = T1064[T1060];
  assign T1060 = T1061;
  assign T1061 = T1062;
  assign T1062 = {12'h0/* 0*/, T1063};
  assign T1063 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1064 = T1065;
  assign T1065 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1073[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = {12'h0/* 0*/, T1072};
  assign T1072 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1073 = T1074;
  assign T1074 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1075 = T1076;
  assign T1076 = T1077;
  assign T1077 = T1082[T1078];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = {12'h0/* 0*/, T1081};
  assign T1081 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1082 = T1083;
  assign T1083 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule


module io_tile_sp_0(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [339:0] io_chanxy_in,
    output[99:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[99:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_wc_1(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [359:0] io_chanxy_in,
    input [159:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[39:0] io_chanxy_out);

  wire[39:0] T0;
  wire[39:0] T1;
  wire[38:0] T2;
  wire[38:0] T3;
  wire[37:0] T4;
  wire[37:0] T5;
  wire[36:0] T6;
  wire[36:0] T7;
  wire[35:0] T8;
  wire[35:0] T9;
  wire[34:0] T10;
  wire[34:0] T11;
  wire[33:0] T12;
  wire[33:0] T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[31:0] T16;
  wire[31:0] T17;
  wire[30:0] T18;
  wire[30:0] T19;
  wire[29:0] T20;
  wire[29:0] T21;
  wire[28:0] T22;
  wire[28:0] T23;
  wire[27:0] T24;
  wire[27:0] T25;
  wire[26:0] T26;
  wire[26:0] T27;
  wire[25:0] T28;
  wire[25:0] T29;
  wire[24:0] T30;
  wire[24:0] T31;
  wire[23:0] T32;
  wire[23:0] T33;
  wire[22:0] T34;
  wire[22:0] T35;
  wire[21:0] T36;
  wire[21:0] T37;
  wire[20:0] T38;
  wire[20:0] T39;
  wire[19:0] T40;
  wire[19:0] T41;
  wire[18:0] T42;
  wire[18:0] T43;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[16:0] T46;
  wire[16:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[14:0] T50;
  wire[14:0] T51;
  wire[13:0] T52;
  wire[13:0] T53;
  wire[12:0] T54;
  wire[12:0] T55;
  wire[11:0] T56;
  wire[11:0] T57;
  wire[10:0] T58;
  wire[10:0] T59;
  wire[9:0] T60;
  wire[9:0] T61;
  wire[8:0] T62;
  wire[8:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire[4:0] T70;
  wire[4:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire[8:0] T84;
  wire[8:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire[8:0] T92;
  wire[8:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire[3:0] T99;
  wire[8:0] T100;
  wire[8:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[8:0] T108;
  wire[8:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire[8:0] T116;
  wire[8:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[8:0] T124;
  wire[8:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[8:0] T132;
  wire[8:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire[8:0] T140;
  wire[8:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[3:0] T146;
  wire[3:0] T147;
  wire[8:0] T148;
  wire[8:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] T154;
  wire[3:0] T155;
  wire[8:0] T156;
  wire[8:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[3:0] T161;
  wire[3:0] T162;
  wire[3:0] T163;
  wire[8:0] T164;
  wire[8:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire[8:0] T172;
  wire[8:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire[3:0] T177;
  wire[3:0] T178;
  wire[3:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire[3:0] T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[8:0] T188;
  wire[8:0] T189;
  wire T190;
  wire T191;
  wire T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire[8:0] T196;
  wire[8:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire[3:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[8:0] T204;
  wire[8:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire[3:0] T209;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[8:0] T212;
  wire[8:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] T219;
  wire[8:0] T220;
  wire[8:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire[3:0] T225;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[8:0] T228;
  wire[8:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[8:0] T236;
  wire[8:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[8:0] T244;
  wire[8:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[3:0] T249;
  wire[3:0] T250;
  wire[3:0] T251;
  wire[8:0] T252;
  wire[8:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[8:0] T260;
  wire[8:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] T265;
  wire[3:0] T266;
  wire[3:0] T267;
  wire[8:0] T268;
  wire[8:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire[3:0] T273;
  wire[3:0] T274;
  wire[3:0] T275;
  wire[8:0] T276;
  wire[8:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[8:0] T284;
  wire[8:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[8:0] T292;
  wire[8:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[8:0] T300;
  wire[8:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[8:0] T308;
  wire[8:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[8:0] T316;
  wire[8:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[8:0] T324;
  wire[8:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[8:0] T332;
  wire[8:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[8:0] T340;
  wire[8:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[8:0] T348;
  wire[8:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[8:0] T356;
  wire[8:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[8:0] T364;
  wire[8:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[8:0] T372;
  wire[8:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[8:0] T380;
  wire[8:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[8:0] T388;
  wire[8:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[8:0] T396;
  wire[8:0] T397;
  wire[7:0] T398;
  wire[7:0] T399;
  wire[6:0] T400;
  wire[6:0] T401;
  wire[5:0] T402;
  wire[5:0] T403;
  wire[4:0] T404;
  wire[4:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire[2:0] T408;
  wire[2:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire T412;
  wire T413;
  wire T414;
  wire[15:0] T415;
  wire[15:0] T416;
  wire[15:0] T417;
  wire[3:0] T418;
  wire[15:0] T419;
  wire[15:0] T420;
  wire T421;
  wire T422;
  wire T423;
  wire[15:0] T424;
  wire[15:0] T425;
  wire[15:0] T426;
  wire[3:0] T427;
  wire[15:0] T428;
  wire[15:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[15:0] T433;
  wire[15:0] T434;
  wire[15:0] T435;
  wire[3:0] T436;
  wire[15:0] T437;
  wire[15:0] T438;
  wire T439;
  wire T440;
  wire T441;
  wire[15:0] T442;
  wire[15:0] T443;
  wire[15:0] T444;
  wire[3:0] T445;
  wire[15:0] T446;
  wire[15:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[15:0] T451;
  wire[15:0] T452;
  wire[15:0] T453;
  wire[3:0] T454;
  wire[15:0] T455;
  wire[15:0] T456;
  wire T457;
  wire T458;
  wire T459;
  wire[15:0] T460;
  wire[15:0] T461;
  wire[15:0] T462;
  wire[3:0] T463;
  wire[15:0] T464;
  wire[15:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire[15:0] T469;
  wire[15:0] T470;
  wire[15:0] T471;
  wire[3:0] T472;
  wire[15:0] T473;
  wire[15:0] T474;
  wire T475;
  wire T476;
  wire T477;
  wire[15:0] T478;
  wire[15:0] T479;
  wire[15:0] T480;
  wire[3:0] T481;
  wire[15:0] T482;
  wire[15:0] T483;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T390, T2};
  assign T2 = T3;
  assign T3 = {T382, T4};
  assign T4 = T5;
  assign T5 = {T374, T6};
  assign T6 = T7;
  assign T7 = {T366, T8};
  assign T8 = T9;
  assign T9 = {T358, T10};
  assign T10 = T11;
  assign T11 = {T350, T12};
  assign T12 = T13;
  assign T13 = {T342, T14};
  assign T14 = T15;
  assign T15 = {T334, T16};
  assign T16 = T17;
  assign T17 = {T326, T18};
  assign T18 = T19;
  assign T19 = {T318, T20};
  assign T20 = T21;
  assign T21 = {T310, T22};
  assign T22 = T23;
  assign T23 = {T302, T24};
  assign T24 = T25;
  assign T25 = {T294, T26};
  assign T26 = T27;
  assign T27 = {T286, T28};
  assign T28 = T29;
  assign T29 = {T278, T30};
  assign T30 = T31;
  assign T31 = {T270, T32};
  assign T32 = T33;
  assign T33 = {T262, T34};
  assign T34 = T35;
  assign T35 = {T254, T36};
  assign T36 = T37;
  assign T37 = {T246, T38};
  assign T38 = T39;
  assign T39 = {T238, T40};
  assign T40 = T41;
  assign T41 = {T230, T42};
  assign T42 = T43;
  assign T43 = {T222, T44};
  assign T44 = T45;
  assign T45 = {T214, T46};
  assign T46 = T47;
  assign T47 = {T206, T48};
  assign T48 = T49;
  assign T49 = {T198, T50};
  assign T50 = T51;
  assign T51 = {T190, T52};
  assign T52 = T53;
  assign T53 = {T182, T54};
  assign T54 = T55;
  assign T55 = {T174, T56};
  assign T56 = T57;
  assign T57 = {T166, T58};
  assign T58 = T59;
  assign T59 = {T158, T60};
  assign T60 = T61;
  assign T61 = {T150, T62};
  assign T62 = T63;
  assign T63 = {T142, T64};
  assign T64 = T65;
  assign T65 = {T134, T66};
  assign T66 = T67;
  assign T67 = {T126, T68};
  assign T68 = T69;
  assign T69 = {T118, T70};
  assign T70 = T71;
  assign T71 = {T110, T72};
  assign T72 = T73;
  assign T73 = {T102, T74};
  assign T74 = T75;
  assign T75 = {T94, T76};
  assign T76 = T77;
  assign T77 = {T86, T78};
  assign T78 = T79;
  assign T79 = T80;
  assign T80 = T84[T81];
  assign T81 = T82;
  assign T82 = T83;
  assign T83 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T84 = T85;
  assign T85 = io_chanxy_in[4'h8/* 8*/:1'h0/* 0*/];
  assign T86 = T87;
  assign T87 = T88;
  assign T88 = T92[T89];
  assign T89 = T90;
  assign T90 = T91;
  assign T91 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T92 = T93;
  assign T93 = io_chanxy_in[5'h11/* 17*/:4'h9/* 9*/];
  assign T94 = T95;
  assign T95 = T96;
  assign T96 = T100[T97];
  assign T97 = T98;
  assign T98 = T99;
  assign T99 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T100 = T101;
  assign T101 = io_chanxy_in[5'h1a/* 26*/:5'h12/* 18*/];
  assign T102 = T103;
  assign T103 = T104;
  assign T104 = T108[T105];
  assign T105 = T106;
  assign T106 = T107;
  assign T107 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T108 = T109;
  assign T109 = io_chanxy_in[6'h23/* 35*/:5'h1b/* 27*/];
  assign T110 = T111;
  assign T111 = T112;
  assign T112 = T116[T113];
  assign T113 = T114;
  assign T114 = T115;
  assign T115 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T116 = T117;
  assign T117 = io_chanxy_in[6'h2c/* 44*/:6'h24/* 36*/];
  assign T118 = T119;
  assign T119 = T120;
  assign T120 = T124[T121];
  assign T121 = T122;
  assign T122 = T123;
  assign T123 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T124 = T125;
  assign T125 = io_chanxy_in[6'h35/* 53*/:6'h2d/* 45*/];
  assign T126 = T127;
  assign T127 = T128;
  assign T128 = T132[T129];
  assign T129 = T130;
  assign T130 = T131;
  assign T131 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T132 = T133;
  assign T133 = io_chanxy_in[6'h3e/* 62*/:6'h36/* 54*/];
  assign T134 = T135;
  assign T135 = T136;
  assign T136 = T140[T137];
  assign T137 = T138;
  assign T138 = T139;
  assign T139 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T140 = T141;
  assign T141 = io_chanxy_in[7'h47/* 71*/:6'h3f/* 63*/];
  assign T142 = T143;
  assign T143 = T144;
  assign T144 = T148[T145];
  assign T145 = T146;
  assign T146 = T147;
  assign T147 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T148 = T149;
  assign T149 = io_chanxy_in[7'h50/* 80*/:7'h48/* 72*/];
  assign T150 = T151;
  assign T151 = T152;
  assign T152 = T156[T153];
  assign T153 = T154;
  assign T154 = T155;
  assign T155 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T156 = T157;
  assign T157 = io_chanxy_in[7'h59/* 89*/:7'h51/* 81*/];
  assign T158 = T159;
  assign T159 = T160;
  assign T160 = T164[T161];
  assign T161 = T162;
  assign T162 = T163;
  assign T163 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T164 = T165;
  assign T165 = io_chanxy_in[7'h62/* 98*/:7'h5a/* 90*/];
  assign T166 = T167;
  assign T167 = T168;
  assign T168 = T172[T169];
  assign T169 = T170;
  assign T170 = T171;
  assign T171 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T172 = T173;
  assign T173 = io_chanxy_in[7'h6b/* 107*/:7'h63/* 99*/];
  assign T174 = T175;
  assign T175 = T176;
  assign T176 = T180[T177];
  assign T177 = T178;
  assign T178 = T179;
  assign T179 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T180 = T181;
  assign T181 = io_chanxy_in[7'h74/* 116*/:7'h6c/* 108*/];
  assign T182 = T183;
  assign T183 = T184;
  assign T184 = T188[T185];
  assign T185 = T186;
  assign T186 = T187;
  assign T187 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T188 = T189;
  assign T189 = io_chanxy_in[7'h7d/* 125*/:7'h75/* 117*/];
  assign T190 = T191;
  assign T191 = T192;
  assign T192 = T196[T193];
  assign T193 = T194;
  assign T194 = T195;
  assign T195 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T196 = T197;
  assign T197 = io_chanxy_in[8'h86/* 134*/:7'h7e/* 126*/];
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[8'h8f/* 143*/:8'h87/* 135*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[8'h98/* 152*/:8'h90/* 144*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[8'ha1/* 161*/:8'h99/* 153*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[8'haa/* 170*/:8'ha2/* 162*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[8'hb3/* 179*/:8'hab/* 171*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[8'hbc/* 188*/:8'hb4/* 180*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[8'hc5/* 197*/:8'hbd/* 189*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[8'hce/* 206*/:8'hc6/* 198*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[8'hd7/* 215*/:8'hcf/* 207*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[8'he0/* 224*/:8'hd8/* 216*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[8'he9/* 233*/:8'he1/* 225*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[8'hf2/* 242*/:8'hea/* 234*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[8'hfb/* 251*/:8'hf3/* 243*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[9'h104/* 260*/:8'hfc/* 252*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[9'h10d/* 269*/:9'h105/* 261*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[9'h116/* 278*/:9'h10e/* 270*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[9'h11f/* 287*/:9'h117/* 279*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[9'h128/* 296*/:9'h120/* 288*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[9'h131/* 305*/:9'h129/* 297*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[9'h13a/* 314*/:9'h132/* 306*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[9'h143/* 323*/:9'h13b/* 315*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[9'h14c/* 332*/:9'h144/* 324*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[9'h155/* 341*/:9'h14d/* 333*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[9'h15e/* 350*/:9'h156/* 342*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[9'h167/* 359*/:9'h15f/* 351*/];
  assign io_ipin_out = T398;
  assign T398 = T399;
  assign T399 = {T475, T400};
  assign T400 = T401;
  assign T401 = {T466, T402};
  assign T402 = T403;
  assign T403 = {T457, T404};
  assign T404 = T405;
  assign T405 = {T448, T406};
  assign T406 = T407;
  assign T407 = {T439, T408};
  assign T408 = T409;
  assign T409 = {T430, T410};
  assign T410 = T411;
  assign T411 = {T421, T412};
  assign T412 = T413;
  assign T413 = T414;
  assign T414 = T419[T415];
  assign T415 = T416;
  assign T416 = T417;
  assign T417 = {12'h0/* 0*/, T418};
  assign T418 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T419 = T420;
  assign T420 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = T428[T424];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = {12'h0/* 0*/, T427};
  assign T427 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T428 = T429;
  assign T429 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T437[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = {12'h0/* 0*/, T436};
  assign T436 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T437 = T438;
  assign T438 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T439 = T440;
  assign T440 = T441;
  assign T441 = T446[T442];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = {12'h0/* 0*/, T445};
  assign T445 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T446 = T447;
  assign T447 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T455[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = {12'h0/* 0*/, T454};
  assign T454 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T455 = T456;
  assign T456 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = T464[T460];
  assign T460 = T461;
  assign T461 = T462;
  assign T462 = {12'h0/* 0*/, T463};
  assign T463 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T464 = T465;
  assign T465 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T473[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = {12'h0/* 0*/, T472};
  assign T472 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T473 = T474;
  assign T474 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = T482[T478];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = {12'h0/* 0*/, T481};
  assign T481 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T482 = T483;
  assign T483 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule

module io_tile_sp_1(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [359:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_2(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [359:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_3(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [359:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_wc_2(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [339:0] io_chanxy_in,
    input [159:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[99:0] io_chanxy_out);

  wire[99:0] T0;
  wire[99:0] T1;
  wire[98:0] T2;
  wire[98:0] T3;
  wire[97:0] T4;
  wire[97:0] T5;
  wire[96:0] T6;
  wire[96:0] T7;
  wire[95:0] T8;
  wire[95:0] T9;
  wire[94:0] T10;
  wire[94:0] T11;
  wire[93:0] T12;
  wire[93:0] T13;
  wire[92:0] T14;
  wire[92:0] T15;
  wire[91:0] T16;
  wire[91:0] T17;
  wire[90:0] T18;
  wire[90:0] T19;
  wire[89:0] T20;
  wire[89:0] T21;
  wire[88:0] T22;
  wire[88:0] T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[86:0] T26;
  wire[86:0] T27;
  wire[85:0] T28;
  wire[85:0] T29;
  wire[84:0] T30;
  wire[84:0] T31;
  wire[83:0] T32;
  wire[83:0] T33;
  wire[82:0] T34;
  wire[82:0] T35;
  wire[81:0] T36;
  wire[81:0] T37;
  wire[80:0] T38;
  wire[80:0] T39;
  wire[79:0] T40;
  wire[79:0] T41;
  wire[78:0] T42;
  wire[78:0] T43;
  wire[77:0] T44;
  wire[77:0] T45;
  wire[76:0] T46;
  wire[76:0] T47;
  wire[75:0] T48;
  wire[75:0] T49;
  wire[74:0] T50;
  wire[74:0] T51;
  wire[73:0] T52;
  wire[73:0] T53;
  wire[72:0] T54;
  wire[72:0] T55;
  wire[71:0] T56;
  wire[71:0] T57;
  wire[70:0] T58;
  wire[70:0] T59;
  wire[69:0] T60;
  wire[69:0] T61;
  wire[68:0] T62;
  wire[68:0] T63;
  wire[67:0] T64;
  wire[67:0] T65;
  wire[66:0] T66;
  wire[66:0] T67;
  wire[65:0] T68;
  wire[65:0] T69;
  wire[64:0] T70;
  wire[64:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[62:0] T74;
  wire[62:0] T75;
  wire[61:0] T76;
  wire[61:0] T77;
  wire[60:0] T78;
  wire[60:0] T79;
  wire[59:0] T80;
  wire[59:0] T81;
  wire[58:0] T82;
  wire[58:0] T83;
  wire[57:0] T84;
  wire[57:0] T85;
  wire[56:0] T86;
  wire[56:0] T87;
  wire[55:0] T88;
  wire[55:0] T89;
  wire[54:0] T90;
  wire[54:0] T91;
  wire[53:0] T92;
  wire[53:0] T93;
  wire[52:0] T94;
  wire[52:0] T95;
  wire[51:0] T96;
  wire[51:0] T97;
  wire[50:0] T98;
  wire[50:0] T99;
  wire[49:0] T100;
  wire[49:0] T101;
  wire[48:0] T102;
  wire[48:0] T103;
  wire[47:0] T104;
  wire[47:0] T105;
  wire[46:0] T106;
  wire[46:0] T107;
  wire[45:0] T108;
  wire[45:0] T109;
  wire[44:0] T110;
  wire[44:0] T111;
  wire[43:0] T112;
  wire[43:0] T113;
  wire[42:0] T114;
  wire[42:0] T115;
  wire[41:0] T116;
  wire[41:0] T117;
  wire[40:0] T118;
  wire[40:0] T119;
  wire[39:0] T120;
  wire[39:0] T121;
  wire[38:0] T122;
  wire[38:0] T123;
  wire[37:0] T124;
  wire[37:0] T125;
  wire[36:0] T126;
  wire[36:0] T127;
  wire[35:0] T128;
  wire[35:0] T129;
  wire[34:0] T130;
  wire[34:0] T131;
  wire[33:0] T132;
  wire[33:0] T133;
  wire[32:0] T134;
  wire[32:0] T135;
  wire[31:0] T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire[30:0] T139;
  wire[29:0] T140;
  wire[29:0] T141;
  wire[28:0] T142;
  wire[28:0] T143;
  wire[27:0] T144;
  wire[27:0] T145;
  wire[26:0] T146;
  wire[26:0] T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire[24:0] T150;
  wire[24:0] T151;
  wire[23:0] T152;
  wire[23:0] T153;
  wire[22:0] T154;
  wire[22:0] T155;
  wire[21:0] T156;
  wire[21:0] T157;
  wire[20:0] T158;
  wire[20:0] T159;
  wire[19:0] T160;
  wire[19:0] T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[17:0] T164;
  wire[17:0] T165;
  wire[16:0] T166;
  wire[16:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire[14:0] T170;
  wire[14:0] T171;
  wire[13:0] T172;
  wire[13:0] T173;
  wire[12:0] T174;
  wire[12:0] T175;
  wire[11:0] T176;
  wire[11:0] T177;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[9:0] T180;
  wire[9:0] T181;
  wire[8:0] T182;
  wire[8:0] T183;
  wire[7:0] T184;
  wire[7:0] T185;
  wire[6:0] T186;
  wire[6:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[1:0] T260;
  wire[1:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[3:0] T681;
  wire[3:0] T682;
  wire[3:0] T683;
  wire[8:0] T684;
  wire[8:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[8:0] T700;
  wire[8:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[3:0] T713;
  wire[3:0] T714;
  wire[3:0] T715;
  wire[8:0] T716;
  wire[8:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[3:0] T729;
  wire[3:0] T730;
  wire[3:0] T731;
  wire[8:0] T732;
  wire[8:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[3:0] T745;
  wire[3:0] T746;
  wire[3:0] T747;
  wire[8:0] T748;
  wire[8:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire[8:0] T764;
  wire[8:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[8:0] T780;
  wire[8:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[3:0] T793;
  wire[3:0] T794;
  wire[3:0] T795;
  wire[8:0] T796;
  wire[8:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[3:0] T809;
  wire[3:0] T810;
  wire[3:0] T811;
  wire[8:0] T812;
  wire[8:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[8:0] T828;
  wire[8:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[3:0] T841;
  wire[3:0] T842;
  wire[3:0] T843;
  wire[8:0] T844;
  wire[8:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[8:0] T860;
  wire[8:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T875;
  wire[8:0] T876;
  wire[8:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[3:0] T890;
  wire[3:0] T891;
  wire[8:0] T892;
  wire[8:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[3:0] T905;
  wire[3:0] T906;
  wire[3:0] T907;
  wire[8:0] T908;
  wire[8:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[3:0] T921;
  wire[3:0] T922;
  wire[3:0] T923;
  wire[8:0] T924;
  wire[8:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[8:0] T940;
  wire[8:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[3:0] T953;
  wire[3:0] T954;
  wire[3:0] T955;
  wire[8:0] T956;
  wire[8:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[3:0] T969;
  wire[3:0] T970;
  wire[3:0] T971;
  wire[8:0] T972;
  wire[8:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[3:0] T985;
  wire[3:0] T986;
  wire[3:0] T987;
  wire[8:0] T988;
  wire[8:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire[7:0] T998;
  wire[7:0] T999;
  wire[6:0] T1000;
  wire[6:0] T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[4:0] T1004;
  wire[4:0] T1005;
  wire[3:0] T1006;
  wire[3:0] T1007;
  wire[2:0] T1008;
  wire[2:0] T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire[15:0] T1015;
  wire[15:0] T1016;
  wire[15:0] T1017;
  wire[3:0] T1018;
  wire[15:0] T1019;
  wire[15:0] T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[15:0] T1024;
  wire[15:0] T1025;
  wire[15:0] T1026;
  wire[3:0] T1027;
  wire[15:0] T1028;
  wire[15:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[15:0] T1033;
  wire[15:0] T1034;
  wire[15:0] T1035;
  wire[3:0] T1036;
  wire[15:0] T1037;
  wire[15:0] T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire[15:0] T1042;
  wire[15:0] T1043;
  wire[15:0] T1044;
  wire[3:0] T1045;
  wire[15:0] T1046;
  wire[15:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire[15:0] T1051;
  wire[15:0] T1052;
  wire[15:0] T1053;
  wire[3:0] T1054;
  wire[15:0] T1055;
  wire[15:0] T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[15:0] T1060;
  wire[15:0] T1061;
  wire[15:0] T1062;
  wire[3:0] T1063;
  wire[15:0] T1064;
  wire[15:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[15:0] T1069;
  wire[15:0] T1070;
  wire[15:0] T1071;
  wire[3:0] T1072;
  wire[15:0] T1073;
  wire[15:0] T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire[15:0] T1078;
  wire[15:0] T1079;
  wire[15:0] T1080;
  wire[3:0] T1081;
  wire[15:0] T1082;
  wire[15:0] T1083;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T990, T2};
  assign T2 = T3;
  assign T3 = {T982, T4};
  assign T4 = T5;
  assign T5 = {T974, T6};
  assign T6 = T7;
  assign T7 = {T966, T8};
  assign T8 = T9;
  assign T9 = {T958, T10};
  assign T10 = T11;
  assign T11 = {T950, T12};
  assign T12 = T13;
  assign T13 = {T942, T14};
  assign T14 = T15;
  assign T15 = {T934, T16};
  assign T16 = T17;
  assign T17 = {T926, T18};
  assign T18 = T19;
  assign T19 = {T918, T20};
  assign T20 = T21;
  assign T21 = {T910, T22};
  assign T22 = T23;
  assign T23 = {T902, T24};
  assign T24 = T25;
  assign T25 = {T894, T26};
  assign T26 = T27;
  assign T27 = {T886, T28};
  assign T28 = T29;
  assign T29 = {T878, T30};
  assign T30 = T31;
  assign T31 = {T870, T32};
  assign T32 = T33;
  assign T33 = {T862, T34};
  assign T34 = T35;
  assign T35 = {T854, T36};
  assign T36 = T37;
  assign T37 = {T846, T38};
  assign T38 = T39;
  assign T39 = {T838, T40};
  assign T40 = T41;
  assign T41 = {T830, T42};
  assign T42 = T43;
  assign T43 = {T822, T44};
  assign T44 = T45;
  assign T45 = {T814, T46};
  assign T46 = T47;
  assign T47 = {T806, T48};
  assign T48 = T49;
  assign T49 = {T798, T50};
  assign T50 = T51;
  assign T51 = {T790, T52};
  assign T52 = T53;
  assign T53 = {T782, T54};
  assign T54 = T55;
  assign T55 = {T774, T56};
  assign T56 = T57;
  assign T57 = {T766, T58};
  assign T58 = T59;
  assign T59 = {T758, T60};
  assign T60 = T61;
  assign T61 = {T750, T62};
  assign T62 = T63;
  assign T63 = {T742, T64};
  assign T64 = T65;
  assign T65 = {T734, T66};
  assign T66 = T67;
  assign T67 = {T726, T68};
  assign T68 = T69;
  assign T69 = {T718, T70};
  assign T70 = T71;
  assign T71 = {T710, T72};
  assign T72 = T73;
  assign T73 = {T702, T74};
  assign T74 = T75;
  assign T75 = {T694, T76};
  assign T76 = T77;
  assign T77 = {T686, T78};
  assign T78 = T79;
  assign T79 = {T678, T80};
  assign T80 = T81;
  assign T81 = {T670, T82};
  assign T82 = T83;
  assign T83 = {T662, T84};
  assign T84 = T85;
  assign T85 = {T654, T86};
  assign T86 = T87;
  assign T87 = {T646, T88};
  assign T88 = T89;
  assign T89 = {T638, T90};
  assign T90 = T91;
  assign T91 = {T630, T92};
  assign T92 = T93;
  assign T93 = {T622, T94};
  assign T94 = T95;
  assign T95 = {T614, T96};
  assign T96 = T97;
  assign T97 = {T606, T98};
  assign T98 = T99;
  assign T99 = {T598, T100};
  assign T100 = T101;
  assign T101 = {T590, T102};
  assign T102 = T103;
  assign T103 = {T582, T104};
  assign T104 = T105;
  assign T105 = {T574, T106};
  assign T106 = T107;
  assign T107 = {T566, T108};
  assign T108 = T109;
  assign T109 = {T558, T110};
  assign T110 = T111;
  assign T111 = {T550, T112};
  assign T112 = T113;
  assign T113 = {T542, T114};
  assign T114 = T115;
  assign T115 = {T534, T116};
  assign T116 = T117;
  assign T117 = {T526, T118};
  assign T118 = T119;
  assign T119 = {T518, T120};
  assign T120 = T121;
  assign T121 = {T510, T122};
  assign T122 = T123;
  assign T123 = {T502, T124};
  assign T124 = T125;
  assign T125 = {T494, T126};
  assign T126 = T127;
  assign T127 = {T486, T128};
  assign T128 = T129;
  assign T129 = {T478, T130};
  assign T130 = T131;
  assign T131 = {T470, T132};
  assign T132 = T133;
  assign T133 = {T462, T134};
  assign T134 = T135;
  assign T135 = {T454, T136};
  assign T136 = T137;
  assign T137 = {T446, T138};
  assign T138 = T139;
  assign T139 = {T438, T140};
  assign T140 = T141;
  assign T141 = {T430, T142};
  assign T142 = T143;
  assign T143 = {T422, T144};
  assign T144 = T145;
  assign T145 = {T414, T146};
  assign T146 = T147;
  assign T147 = {T406, T148};
  assign T148 = T149;
  assign T149 = {T398, T150};
  assign T150 = T151;
  assign T151 = {T390, T152};
  assign T152 = T153;
  assign T153 = {T382, T154};
  assign T154 = T155;
  assign T155 = {T374, T156};
  assign T156 = T157;
  assign T157 = {T366, T158};
  assign T158 = T159;
  assign T159 = {T358, T160};
  assign T160 = T161;
  assign T161 = {T350, T162};
  assign T162 = T163;
  assign T163 = {T342, T164};
  assign T164 = T165;
  assign T165 = {T334, T166};
  assign T166 = T167;
  assign T167 = {T326, T168};
  assign T168 = T169;
  assign T169 = {T318, T170};
  assign T170 = T171;
  assign T171 = {T310, T172};
  assign T172 = T173;
  assign T173 = {T302, T174};
  assign T174 = T175;
  assign T175 = {T294, T176};
  assign T176 = T177;
  assign T177 = {T286, T178};
  assign T178 = T179;
  assign T179 = {T278, T180};
  assign T180 = T181;
  assign T181 = {T270, T182};
  assign T182 = T183;
  assign T183 = {T262, T184};
  assign T184 = T185;
  assign T185 = {T254, T186};
  assign T186 = T187;
  assign T187 = {T246, T188};
  assign T188 = T189;
  assign T189 = {T238, T190};
  assign T190 = T191;
  assign T191 = {T230, T192};
  assign T192 = T193;
  assign T193 = {T222, T194};
  assign T194 = T195;
  assign T195 = {T214, T196};
  assign T196 = T197;
  assign T197 = {T206, T198};
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[2'h2/* 2*/:2'h2/* 2*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[3'h5/* 5*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[2'h3/* 3*/:2'h3/* 3*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[3'h7/* 7*/:3'h6/* 6*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[3'h4/* 4*/:3'h4/* 4*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[4'h9/* 9*/:4'h8/* 8*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[3'h5/* 5*/:3'h5/* 5*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[4'hb/* 11*/:4'ha/* 10*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[3'h6/* 6*/:3'h6/* 6*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[4'hd/* 13*/:4'hc/* 12*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[4'hf/* 15*/:4'he/* 14*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[5'h11/* 17*/:5'h10/* 16*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[4'hb/* 11*/:4'hb/* 11*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[6'h33/* 51*/:6'h32/* 50*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[6'h35/* 53*/:6'h34/* 52*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[7'h55/* 85*/:7'h54/* 84*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[6'h2b/* 43*/:6'h2b/* 43*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[7'h57/* 87*/:7'h56/* 86*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[6'h2c/* 44*/:6'h2c/* 44*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[7'h59/* 89*/:7'h58/* 88*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[6'h2d/* 45*/:6'h2d/* 45*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h2e/* 46*/:6'h2e/* 46*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h2f/* 47*/:6'h2f/* 47*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[6'h34/* 52*/:6'h34/* 52*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[6'h35/* 53*/:6'h35/* 53*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[7'h71/* 113*/:7'h70/* 112*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h73/* 115*/:7'h72/* 114*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h75/* 117*/:7'h74/* 116*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[7'h77/* 119*/:7'h76/* 118*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'h80/* 128*/:7'h78/* 120*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'h82/* 130*/:8'h81/* 129*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h44/* 68*/:7'h41/* 65*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'h8b/* 139*/:8'h83/* 131*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h45/* 69*/:7'h45/* 69*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h49/* 73*/:7'h46/* 70*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'h96/* 150*/:8'h8e/* 142*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'h98/* 152*/:8'h97/* 151*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'ha1/* 161*/:8'h99/* 153*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'hac/* 172*/:8'ha4/* 164*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h54/* 84*/:7'h54/* 84*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'hae/* 174*/:8'had/* 173*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h58/* 88*/:7'h55/* 85*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'hb7/* 183*/:8'haf/* 175*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'hc2/* 194*/:8'hba/* 186*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h62/* 98*/:7'h5f/* 95*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'hcd/* 205*/:8'hc5/* 197*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h63/* 99*/:7'h63/* 99*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'hcf/* 207*/:8'hce/* 206*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'hd8/* 216*/:8'hd0/* 208*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h6c/* 108*/:7'h69/* 105*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'he3/* 227*/:8'hdb/* 219*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h6d/* 109*/:7'h6d/* 109*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'he5/* 229*/:8'he4/* 228*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[7'h71/* 113*/:7'h6e/* 110*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'hee/* 238*/:8'he6/* 230*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[8'hf0/* 240*/:8'hef/* 239*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[8'hf9/* 249*/:8'hf1/* 241*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h104/* 260*/:8'hfc/* 252*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[7'h7c/* 124*/:7'h7c/* 124*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h106/* 262*/:9'h105/* 261*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h80/* 128*/:7'h7d/* 125*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h10f/* 271*/:9'h107/* 263*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h11a/* 282*/:9'h112/* 274*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h8a/* 138*/:8'h87/* 135*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h125/* 293*/:9'h11d/* 285*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h127/* 295*/:9'h126/* 294*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h130/* 304*/:9'h128/* 296*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h132/* 306*/:9'h131/* 305*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'h94/* 148*/:8'h91/* 145*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h13b/* 315*/:9'h133/* 307*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'h95/* 149*/:8'h95/* 149*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h13d/* 317*/:9'h13c/* 316*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h146/* 326*/:9'h13e/* 318*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h151/* 337*/:9'h149/* 329*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign io_ipin_out = T998;
  assign T998 = T999;
  assign T999 = {T1075, T1000};
  assign T1000 = T1001;
  assign T1001 = {T1066, T1002};
  assign T1002 = T1003;
  assign T1003 = {T1057, T1004};
  assign T1004 = T1005;
  assign T1005 = {T1048, T1006};
  assign T1006 = T1007;
  assign T1007 = {T1039, T1008};
  assign T1008 = T1009;
  assign T1009 = {T1030, T1010};
  assign T1010 = T1011;
  assign T1011 = {T1021, T1012};
  assign T1012 = T1013;
  assign T1013 = T1014;
  assign T1014 = T1019[T1015];
  assign T1015 = T1016;
  assign T1016 = T1017;
  assign T1017 = {12'h0/* 0*/, T1018};
  assign T1018 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1019 = T1020;
  assign T1020 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = T1028[T1024];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = {12'h0/* 0*/, T1027};
  assign T1027 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1028 = T1029;
  assign T1029 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1037[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = {12'h0/* 0*/, T1036};
  assign T1036 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1037 = T1038;
  assign T1038 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1039 = T1040;
  assign T1040 = T1041;
  assign T1041 = T1046[T1042];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = {12'h0/* 0*/, T1045};
  assign T1045 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1046 = T1047;
  assign T1047 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1048 = T1049;
  assign T1049 = T1050;
  assign T1050 = T1055[T1051];
  assign T1051 = T1052;
  assign T1052 = T1053;
  assign T1053 = {12'h0/* 0*/, T1054};
  assign T1054 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1055 = T1056;
  assign T1056 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = T1064[T1060];
  assign T1060 = T1061;
  assign T1061 = T1062;
  assign T1062 = {12'h0/* 0*/, T1063};
  assign T1063 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1064 = T1065;
  assign T1065 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1073[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = {12'h0/* 0*/, T1072};
  assign T1072 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1073 = T1074;
  assign T1074 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1075 = T1076;
  assign T1076 = T1077;
  assign T1077 = T1082[T1078];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = {12'h0/* 0*/, T1081};
  assign T1081 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1082 = T1083;
  assign T1083 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule

module io_tile_sp_4(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [339:0] io_chanxy_in,
    output[99:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[99:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_2 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_woc(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    output[7:0] io_ipin_out);

  wire[7:0] T0;
  wire[7:0] T1;
  wire[6:0] T2;
  wire[6:0] T3;
  wire[5:0] T4;
  wire[5:0] T5;
  wire[4:0] T6;
  wire[4:0] T7;
  wire[3:0] T8;
  wire[3:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[1:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire[15:0] T17;
  wire[15:0] T18;
  wire[15:0] T19;
  wire[3:0] T20;
  wire[15:0] T21;
  wire[15:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire[15:0] T26;
  wire[15:0] T27;
  wire[15:0] T28;
  wire[3:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire T32;
  wire T33;
  wire T34;
  wire[15:0] T35;
  wire[15:0] T36;
  wire[15:0] T37;
  wire[3:0] T38;
  wire[15:0] T39;
  wire[15:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire[15:0] T44;
  wire[15:0] T45;
  wire[15:0] T46;
  wire[3:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire T50;
  wire T51;
  wire T52;
  wire[15:0] T53;
  wire[15:0] T54;
  wire[15:0] T55;
  wire[3:0] T56;
  wire[15:0] T57;
  wire[15:0] T58;
  wire T59;
  wire T60;
  wire T61;
  wire[15:0] T62;
  wire[15:0] T63;
  wire[15:0] T64;
  wire[3:0] T65;
  wire[15:0] T66;
  wire[15:0] T67;
  wire T68;
  wire T69;
  wire T70;
  wire[15:0] T71;
  wire[15:0] T72;
  wire[15:0] T73;
  wire[3:0] T74;
  wire[15:0] T75;
  wire[15:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire[15:0] T82;
  wire[3:0] T83;
  wire[15:0] T84;
  wire[15:0] T85;

  assign io_ipin_out = T0;
  assign T0 = T1;
  assign T1 = {T77, T2};
  assign T2 = T3;
  assign T3 = {T68, T4};
  assign T4 = T5;
  assign T5 = {T59, T6};
  assign T6 = T7;
  assign T7 = {T50, T8};
  assign T8 = T9;
  assign T9 = {T41, T10};
  assign T10 = T11;
  assign T11 = {T32, T12};
  assign T12 = T13;
  assign T13 = {T23, T14};
  assign T14 = T15;
  assign T15 = T16;
  assign T16 = T21[T17];
  assign T17 = T18;
  assign T18 = T19;
  assign T19 = {12'h0/* 0*/, T20};
  assign T20 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T21 = T22;
  assign T22 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T23 = T24;
  assign T24 = T25;
  assign T25 = T30[T26];
  assign T26 = T27;
  assign T27 = T28;
  assign T28 = {12'h0/* 0*/, T29};
  assign T29 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T30 = T31;
  assign T31 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T32 = T33;
  assign T33 = T34;
  assign T34 = T39[T35];
  assign T35 = T36;
  assign T36 = T37;
  assign T37 = {12'h0/* 0*/, T38};
  assign T38 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T39 = T40;
  assign T40 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T41 = T42;
  assign T42 = T43;
  assign T43 = T48[T44];
  assign T44 = T45;
  assign T45 = T46;
  assign T46 = {12'h0/* 0*/, T47};
  assign T47 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T48 = T49;
  assign T49 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T50 = T51;
  assign T51 = T52;
  assign T52 = T57[T53];
  assign T53 = T54;
  assign T54 = T55;
  assign T55 = {12'h0/* 0*/, T56};
  assign T56 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T57 = T58;
  assign T58 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T59 = T60;
  assign T60 = T61;
  assign T61 = T66[T62];
  assign T62 = T63;
  assign T63 = T64;
  assign T64 = {12'h0/* 0*/, T65};
  assign T65 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T66 = T67;
  assign T67 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T68 = T69;
  assign T69 = T70;
  assign T70 = T75[T71];
  assign T71 = T72;
  assign T72 = T73;
  assign T73 = {12'h0/* 0*/, T74};
  assign T74 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T75 = T76;
  assign T76 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T77 = T78;
  assign T78 = T79;
  assign T79 = T84[T80];
  assign T80 = T81;
  assign T81 = T82;
  assign T82 = {12'h0/* 0*/, T83};
  assign T83 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T84 = T85;
  assign T85 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule


module io_tile_sp_5(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_6(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_7(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_8(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_9(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_wc_3(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [355:0] io_chanxy_in,
    input [167:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[99:0] io_chanxy_out);

  wire[99:0] T0;
  wire[99:0] T1;
  wire[98:0] T2;
  wire[98:0] T3;
  wire[97:0] T4;
  wire[97:0] T5;
  wire[96:0] T6;
  wire[96:0] T7;
  wire[95:0] T8;
  wire[95:0] T9;
  wire[94:0] T10;
  wire[94:0] T11;
  wire[93:0] T12;
  wire[93:0] T13;
  wire[92:0] T14;
  wire[92:0] T15;
  wire[91:0] T16;
  wire[91:0] T17;
  wire[90:0] T18;
  wire[90:0] T19;
  wire[89:0] T20;
  wire[89:0] T21;
  wire[88:0] T22;
  wire[88:0] T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[86:0] T26;
  wire[86:0] T27;
  wire[85:0] T28;
  wire[85:0] T29;
  wire[84:0] T30;
  wire[84:0] T31;
  wire[83:0] T32;
  wire[83:0] T33;
  wire[82:0] T34;
  wire[82:0] T35;
  wire[81:0] T36;
  wire[81:0] T37;
  wire[80:0] T38;
  wire[80:0] T39;
  wire[79:0] T40;
  wire[79:0] T41;
  wire[78:0] T42;
  wire[78:0] T43;
  wire[77:0] T44;
  wire[77:0] T45;
  wire[76:0] T46;
  wire[76:0] T47;
  wire[75:0] T48;
  wire[75:0] T49;
  wire[74:0] T50;
  wire[74:0] T51;
  wire[73:0] T52;
  wire[73:0] T53;
  wire[72:0] T54;
  wire[72:0] T55;
  wire[71:0] T56;
  wire[71:0] T57;
  wire[70:0] T58;
  wire[70:0] T59;
  wire[69:0] T60;
  wire[69:0] T61;
  wire[68:0] T62;
  wire[68:0] T63;
  wire[67:0] T64;
  wire[67:0] T65;
  wire[66:0] T66;
  wire[66:0] T67;
  wire[65:0] T68;
  wire[65:0] T69;
  wire[64:0] T70;
  wire[64:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[62:0] T74;
  wire[62:0] T75;
  wire[61:0] T76;
  wire[61:0] T77;
  wire[60:0] T78;
  wire[60:0] T79;
  wire[59:0] T80;
  wire[59:0] T81;
  wire[58:0] T82;
  wire[58:0] T83;
  wire[57:0] T84;
  wire[57:0] T85;
  wire[56:0] T86;
  wire[56:0] T87;
  wire[55:0] T88;
  wire[55:0] T89;
  wire[54:0] T90;
  wire[54:0] T91;
  wire[53:0] T92;
  wire[53:0] T93;
  wire[52:0] T94;
  wire[52:0] T95;
  wire[51:0] T96;
  wire[51:0] T97;
  wire[50:0] T98;
  wire[50:0] T99;
  wire[49:0] T100;
  wire[49:0] T101;
  wire[48:0] T102;
  wire[48:0] T103;
  wire[47:0] T104;
  wire[47:0] T105;
  wire[46:0] T106;
  wire[46:0] T107;
  wire[45:0] T108;
  wire[45:0] T109;
  wire[44:0] T110;
  wire[44:0] T111;
  wire[43:0] T112;
  wire[43:0] T113;
  wire[42:0] T114;
  wire[42:0] T115;
  wire[41:0] T116;
  wire[41:0] T117;
  wire[40:0] T118;
  wire[40:0] T119;
  wire[39:0] T120;
  wire[39:0] T121;
  wire[38:0] T122;
  wire[38:0] T123;
  wire[37:0] T124;
  wire[37:0] T125;
  wire[36:0] T126;
  wire[36:0] T127;
  wire[35:0] T128;
  wire[35:0] T129;
  wire[34:0] T130;
  wire[34:0] T131;
  wire[33:0] T132;
  wire[33:0] T133;
  wire[32:0] T134;
  wire[32:0] T135;
  wire[31:0] T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire[30:0] T139;
  wire[29:0] T140;
  wire[29:0] T141;
  wire[28:0] T142;
  wire[28:0] T143;
  wire[27:0] T144;
  wire[27:0] T145;
  wire[26:0] T146;
  wire[26:0] T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire[24:0] T150;
  wire[24:0] T151;
  wire[23:0] T152;
  wire[23:0] T153;
  wire[22:0] T154;
  wire[22:0] T155;
  wire[21:0] T156;
  wire[21:0] T157;
  wire[20:0] T158;
  wire[20:0] T159;
  wire[19:0] T160;
  wire[19:0] T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[17:0] T164;
  wire[17:0] T165;
  wire[16:0] T166;
  wire[16:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire[14:0] T170;
  wire[14:0] T171;
  wire[13:0] T172;
  wire[13:0] T173;
  wire[12:0] T174;
  wire[12:0] T175;
  wire[11:0] T176;
  wire[11:0] T177;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[9:0] T180;
  wire[9:0] T181;
  wire[8:0] T182;
  wire[8:0] T183;
  wire[7:0] T184;
  wire[7:0] T185;
  wire[6:0] T186;
  wire[6:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire[1:0] T201;
  wire[1:0] T202;
  wire[1:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire[1:0] T209;
  wire[1:0] T210;
  wire[1:0] T211;
  wire[2:0] T212;
  wire[2:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] T219;
  wire[9:0] T220;
  wire[9:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire[1:0] T225;
  wire[1:0] T226;
  wire[1:0] T227;
  wire[2:0] T228;
  wire[2:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire[1:0] T233;
  wire[1:0] T234;
  wire[1:0] T235;
  wire[2:0] T236;
  wire[2:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire[1:0] T241;
  wire[1:0] T242;
  wire[1:0] T243;
  wire[2:0] T244;
  wire[2:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[1:0] T249;
  wire[1:0] T250;
  wire[1:0] T251;
  wire[2:0] T252;
  wire[2:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire[1:0] T265;
  wire[1:0] T266;
  wire[1:0] T267;
  wire[2:0] T268;
  wire[2:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire[1:0] T273;
  wire[1:0] T274;
  wire[1:0] T275;
  wire[2:0] T276;
  wire[2:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[9:0] T300;
  wire[9:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[9:0] T340;
  wire[9:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[9:0] T420;
  wire[9:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[9:0] T460;
  wire[9:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[9:0] T500;
  wire[9:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[8:0] T540;
  wire[8:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[8:0] T580;
  wire[8:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[3:0] T617;
  wire[3:0] T618;
  wire[3:0] T619;
  wire[8:0] T620;
  wire[8:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[3:0] T657;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[8:0] T660;
  wire[8:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[8:0] T700;
  wire[8:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[3:0] T737;
  wire[3:0] T738;
  wire[3:0] T739;
  wire[8:0] T740;
  wire[8:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[8:0] T780;
  wire[8:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[3:0] T817;
  wire[3:0] T818;
  wire[3:0] T819;
  wire[8:0] T820;
  wire[8:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[8:0] T860;
  wire[8:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[8:0] T900;
  wire[8:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[8:0] T940;
  wire[8:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[8:0] T980;
  wire[8:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire[7:0] T998;
  wire[7:0] T999;
  wire[6:0] T1000;
  wire[6:0] T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[4:0] T1004;
  wire[4:0] T1005;
  wire[3:0] T1006;
  wire[3:0] T1007;
  wire[2:0] T1008;
  wire[2:0] T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire[15:0] T1015;
  wire[15:0] T1016;
  wire[15:0] T1017;
  wire[3:0] T1018;
  wire[15:0] T1019;
  wire[15:0] T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[15:0] T1024;
  wire[15:0] T1025;
  wire[15:0] T1026;
  wire[3:0] T1027;
  wire[15:0] T1028;
  wire[15:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[15:0] T1033;
  wire[15:0] T1034;
  wire[15:0] T1035;
  wire[3:0] T1036;
  wire[15:0] T1037;
  wire[15:0] T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire[15:0] T1042;
  wire[15:0] T1043;
  wire[15:0] T1044;
  wire[3:0] T1045;
  wire[15:0] T1046;
  wire[15:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire[15:0] T1051;
  wire[15:0] T1052;
  wire[15:0] T1053;
  wire[3:0] T1054;
  wire[15:0] T1055;
  wire[15:0] T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[15:0] T1060;
  wire[15:0] T1061;
  wire[15:0] T1062;
  wire[3:0] T1063;
  wire[15:0] T1064;
  wire[15:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[15:0] T1069;
  wire[15:0] T1070;
  wire[15:0] T1071;
  wire[3:0] T1072;
  wire[15:0] T1073;
  wire[15:0] T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire[15:0] T1078;
  wire[15:0] T1079;
  wire[15:0] T1080;
  wire[3:0] T1081;
  wire[15:0] T1082;
  wire[15:0] T1083;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T990, T2};
  assign T2 = T3;
  assign T3 = {T982, T4};
  assign T4 = T5;
  assign T5 = {T974, T6};
  assign T6 = T7;
  assign T7 = {T966, T8};
  assign T8 = T9;
  assign T9 = {T958, T10};
  assign T10 = T11;
  assign T11 = {T950, T12};
  assign T12 = T13;
  assign T13 = {T942, T14};
  assign T14 = T15;
  assign T15 = {T934, T16};
  assign T16 = T17;
  assign T17 = {T926, T18};
  assign T18 = T19;
  assign T19 = {T918, T20};
  assign T20 = T21;
  assign T21 = {T910, T22};
  assign T22 = T23;
  assign T23 = {T902, T24};
  assign T24 = T25;
  assign T25 = {T894, T26};
  assign T26 = T27;
  assign T27 = {T886, T28};
  assign T28 = T29;
  assign T29 = {T878, T30};
  assign T30 = T31;
  assign T31 = {T870, T32};
  assign T32 = T33;
  assign T33 = {T862, T34};
  assign T34 = T35;
  assign T35 = {T854, T36};
  assign T36 = T37;
  assign T37 = {T846, T38};
  assign T38 = T39;
  assign T39 = {T838, T40};
  assign T40 = T41;
  assign T41 = {T830, T42};
  assign T42 = T43;
  assign T43 = {T822, T44};
  assign T44 = T45;
  assign T45 = {T814, T46};
  assign T46 = T47;
  assign T47 = {T806, T48};
  assign T48 = T49;
  assign T49 = {T798, T50};
  assign T50 = T51;
  assign T51 = {T790, T52};
  assign T52 = T53;
  assign T53 = {T782, T54};
  assign T54 = T55;
  assign T55 = {T774, T56};
  assign T56 = T57;
  assign T57 = {T766, T58};
  assign T58 = T59;
  assign T59 = {T758, T60};
  assign T60 = T61;
  assign T61 = {T750, T62};
  assign T62 = T63;
  assign T63 = {T742, T64};
  assign T64 = T65;
  assign T65 = {T734, T66};
  assign T66 = T67;
  assign T67 = {T726, T68};
  assign T68 = T69;
  assign T69 = {T718, T70};
  assign T70 = T71;
  assign T71 = {T710, T72};
  assign T72 = T73;
  assign T73 = {T702, T74};
  assign T74 = T75;
  assign T75 = {T694, T76};
  assign T76 = T77;
  assign T77 = {T686, T78};
  assign T78 = T79;
  assign T79 = {T678, T80};
  assign T80 = T81;
  assign T81 = {T670, T82};
  assign T82 = T83;
  assign T83 = {T662, T84};
  assign T84 = T85;
  assign T85 = {T654, T86};
  assign T86 = T87;
  assign T87 = {T646, T88};
  assign T88 = T89;
  assign T89 = {T638, T90};
  assign T90 = T91;
  assign T91 = {T630, T92};
  assign T92 = T93;
  assign T93 = {T622, T94};
  assign T94 = T95;
  assign T95 = {T614, T96};
  assign T96 = T97;
  assign T97 = {T606, T98};
  assign T98 = T99;
  assign T99 = {T598, T100};
  assign T100 = T101;
  assign T101 = {T590, T102};
  assign T102 = T103;
  assign T103 = {T582, T104};
  assign T104 = T105;
  assign T105 = {T574, T106};
  assign T106 = T107;
  assign T107 = {T566, T108};
  assign T108 = T109;
  assign T109 = {T558, T110};
  assign T110 = T111;
  assign T111 = {T550, T112};
  assign T112 = T113;
  assign T113 = {T542, T114};
  assign T114 = T115;
  assign T115 = {T534, T116};
  assign T116 = T117;
  assign T117 = {T526, T118};
  assign T118 = T119;
  assign T119 = {T518, T120};
  assign T120 = T121;
  assign T121 = {T510, T122};
  assign T122 = T123;
  assign T123 = {T502, T124};
  assign T124 = T125;
  assign T125 = {T494, T126};
  assign T126 = T127;
  assign T127 = {T486, T128};
  assign T128 = T129;
  assign T129 = {T478, T130};
  assign T130 = T131;
  assign T131 = {T470, T132};
  assign T132 = T133;
  assign T133 = {T462, T134};
  assign T134 = T135;
  assign T135 = {T454, T136};
  assign T136 = T137;
  assign T137 = {T446, T138};
  assign T138 = T139;
  assign T139 = {T438, T140};
  assign T140 = T141;
  assign T141 = {T430, T142};
  assign T142 = T143;
  assign T143 = {T422, T144};
  assign T144 = T145;
  assign T145 = {T414, T146};
  assign T146 = T147;
  assign T147 = {T406, T148};
  assign T148 = T149;
  assign T149 = {T398, T150};
  assign T150 = T151;
  assign T151 = {T390, T152};
  assign T152 = T153;
  assign T153 = {T382, T154};
  assign T154 = T155;
  assign T155 = {T374, T156};
  assign T156 = T157;
  assign T157 = {T366, T158};
  assign T158 = T159;
  assign T159 = {T358, T160};
  assign T160 = T161;
  assign T161 = {T350, T162};
  assign T162 = T163;
  assign T163 = {T342, T164};
  assign T164 = T165;
  assign T165 = {T334, T166};
  assign T166 = T167;
  assign T167 = {T326, T168};
  assign T168 = T169;
  assign T169 = {T318, T170};
  assign T170 = T171;
  assign T171 = {T310, T172};
  assign T172 = T173;
  assign T173 = {T302, T174};
  assign T174 = T175;
  assign T175 = {T294, T176};
  assign T176 = T177;
  assign T177 = {T286, T178};
  assign T178 = T179;
  assign T179 = {T278, T180};
  assign T180 = T181;
  assign T181 = {T270, T182};
  assign T182 = T183;
  assign T183 = {T262, T184};
  assign T184 = T185;
  assign T185 = {T254, T186};
  assign T186 = T187;
  assign T187 = {T246, T188};
  assign T188 = T189;
  assign T189 = {T238, T190};
  assign T190 = T191;
  assign T191 = {T230, T192};
  assign T192 = T193;
  assign T193 = {T222, T194};
  assign T194 = T195;
  assign T195 = {T214, T196};
  assign T196 = T197;
  assign T197 = {T206, T198};
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[4'hf/* 15*/:3'h6/* 6*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[5'h12/* 18*/:5'h10/* 16*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[5'h15/* 21*/:5'h13/* 19*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[5'h18/* 24*/:5'h16/* 22*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[5'h1b/* 27*/:5'h19/* 25*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[6'h25/* 37*/:5'h1c/* 28*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[5'h15/* 21*/:5'h14/* 20*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[6'h28/* 40*/:6'h26/* 38*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[6'h2b/* 43*/:6'h29/* 41*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[5'h1d/* 29*/:5'h1a/* 26*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[6'h39/* 57*/:6'h30/* 48*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[6'h25/* 37*/:6'h22/* 34*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[7'h4b/* 75*/:7'h42/* 66*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h2d/* 45*/:6'h2a/* 42*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[7'h5d/* 93*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h2e/* 46*/:6'h2e/* 46*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h2f/* 47*/:6'h2f/* 47*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[6'h35/* 53*/:6'h32/* 50*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[7'h6f/* 111*/:7'h66/* 102*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[7'h71/* 113*/:7'h70/* 112*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[7'h73/* 115*/:7'h72/* 114*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h75/* 117*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h77/* 119*/:7'h76/* 118*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h3d/* 61*/:6'h3a/* 58*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[8'h81/* 129*/:7'h78/* 120*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h3e/* 62*/:6'h3e/* 62*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[8'h83/* 131*/:8'h82/* 130*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h3f/* 63*/:6'h3f/* 63*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[8'h85/* 133*/:8'h84/* 132*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[8'h87/* 135*/:8'h86/* 134*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h41/* 65*/:7'h41/* 65*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[8'h93/* 147*/:8'h8a/* 138*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h46/* 70*/:7'h46/* 70*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[8'h95/* 149*/:8'h94/* 148*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h47/* 71*/:7'h47/* 71*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[8'h97/* 151*/:8'h96/* 150*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[8'h99/* 153*/:8'h98/* 152*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[7'h4d/* 77*/:7'h4a/* 74*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[8'ha4/* 164*/:8'h9c/* 156*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[7'h4e/* 78*/:7'h4e/* 78*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[8'ha6/* 166*/:8'ha5/* 165*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[8'ha8/* 168*/:8'ha7/* 167*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[8'haa/* 170*/:8'ha9/* 169*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[8'hac/* 172*/:8'hab/* 171*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[7'h55/* 85*/:7'h52/* 82*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[8'hb5/* 181*/:8'had/* 173*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[8'hbb/* 187*/:8'hba/* 186*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[8'hbd/* 189*/:8'hbc/* 188*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[8'hc6/* 198*/:8'hbe/* 190*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'hca/* 202*/:8'hc9/* 201*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'hcc/* 204*/:8'hcb/* 203*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'hce/* 206*/:8'hcd/* 205*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h65/* 101*/:7'h62/* 98*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'hd7/* 215*/:8'hcf/* 207*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h66/* 102*/:7'h66/* 102*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'hdb/* 219*/:8'hda/* 218*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'hdf/* 223*/:8'hde/* 222*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h6d/* 109*/:7'h6a/* 106*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'he8/* 232*/:8'he0/* 224*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h6e/* 110*/:7'h6e/* 110*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hec/* 236*/:8'heb/* 235*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hee/* 238*/:8'hed/* 237*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'hf0/* 240*/:8'hef/* 239*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'hf9/* 249*/:8'hf1/* 241*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'hfd/* 253*/:8'hfc/* 252*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'hff/* 255*/:8'hfe/* 254*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[9'h101/* 257*/:9'h100/* 256*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h7d/* 125*/:7'h7a/* 122*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[9'h10a/* 266*/:9'h102/* 258*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h110/* 272*/:9'h10f/* 271*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h112/* 274*/:9'h111/* 273*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h11b/* 283*/:9'h113/* 275*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h11d/* 285*/:9'h11c/* 284*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h11f/* 287*/:9'h11e/* 286*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h121/* 289*/:9'h120/* 288*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h123/* 291*/:9'h122/* 290*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h12c/* 300*/:9'h124/* 292*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h130/* 304*/:9'h12f/* 303*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h132/* 306*/:9'h131/* 305*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h134/* 308*/:9'h133/* 307*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h95/* 149*/:8'h92/* 146*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h13d/* 317*/:9'h135/* 309*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h96/* 150*/:8'h96/* 150*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h13f/* 319*/:9'h13e/* 318*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h141/* 321*/:9'h140/* 320*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h143/* 323*/:9'h142/* 322*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h145/* 325*/:9'h144/* 324*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h9d/* 157*/:8'h9a/* 154*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h14e/* 334*/:9'h146/* 326*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h150/* 336*/:9'h14f/* 335*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h152/* 338*/:9'h151/* 337*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h154/* 340*/:9'h153/* 339*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h156/* 342*/:9'h155/* 341*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'ha5/* 165*/:8'ha2/* 162*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h15f/* 351*/:9'h157/* 343*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'ha6/* 166*/:8'ha6/* 166*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h161/* 353*/:9'h160/* 352*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h163/* 355*/:9'h162/* 354*/];
  assign io_ipin_out = T998;
  assign T998 = T999;
  assign T999 = {T1075, T1000};
  assign T1000 = T1001;
  assign T1001 = {T1066, T1002};
  assign T1002 = T1003;
  assign T1003 = {T1057, T1004};
  assign T1004 = T1005;
  assign T1005 = {T1048, T1006};
  assign T1006 = T1007;
  assign T1007 = {T1039, T1008};
  assign T1008 = T1009;
  assign T1009 = {T1030, T1010};
  assign T1010 = T1011;
  assign T1011 = {T1021, T1012};
  assign T1012 = T1013;
  assign T1013 = T1014;
  assign T1014 = T1019[T1015];
  assign T1015 = T1016;
  assign T1016 = T1017;
  assign T1017 = {12'h0/* 0*/, T1018};
  assign T1018 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1019 = T1020;
  assign T1020 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = T1028[T1024];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = {12'h0/* 0*/, T1027};
  assign T1027 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1028 = T1029;
  assign T1029 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1037[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = {12'h0/* 0*/, T1036};
  assign T1036 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1037 = T1038;
  assign T1038 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1039 = T1040;
  assign T1040 = T1041;
  assign T1041 = T1046[T1042];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = {12'h0/* 0*/, T1045};
  assign T1045 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1046 = T1047;
  assign T1047 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1048 = T1049;
  assign T1049 = T1050;
  assign T1050 = T1055[T1051];
  assign T1051 = T1052;
  assign T1052 = T1053;
  assign T1053 = {12'h0/* 0*/, T1054};
  assign T1054 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1055 = T1056;
  assign T1056 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = T1064[T1060];
  assign T1060 = T1061;
  assign T1061 = T1062;
  assign T1062 = {12'h0/* 0*/, T1063};
  assign T1063 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1064 = T1065;
  assign T1065 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1073[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = {12'h0/* 0*/, T1072};
  assign T1072 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1073 = T1074;
  assign T1074 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1075 = T1076;
  assign T1076 = T1077;
  assign T1077 = T1082[T1078];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = {12'h0/* 0*/, T1081};
  assign T1081 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1082 = T1083;
  assign T1083 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule


module io_tile_sp_10(input clk, input reset,
    input [31:0] io_configs_in,
    input [6:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [355:0] io_chanxy_in,
    output[99:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[167:0] T0;
  wire[223:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[99:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hc7/* 199*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_x_loc = T3;
  assign T3 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_3 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_7 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_wc_4(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [375:0] io_chanxy_in,
    input [159:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[39:0] io_chanxy_out);

  wire[39:0] T0;
  wire[39:0] T1;
  wire[38:0] T2;
  wire[38:0] T3;
  wire[37:0] T4;
  wire[37:0] T5;
  wire[36:0] T6;
  wire[36:0] T7;
  wire[35:0] T8;
  wire[35:0] T9;
  wire[34:0] T10;
  wire[34:0] T11;
  wire[33:0] T12;
  wire[33:0] T13;
  wire[32:0] T14;
  wire[32:0] T15;
  wire[31:0] T16;
  wire[31:0] T17;
  wire[30:0] T18;
  wire[30:0] T19;
  wire[29:0] T20;
  wire[29:0] T21;
  wire[28:0] T22;
  wire[28:0] T23;
  wire[27:0] T24;
  wire[27:0] T25;
  wire[26:0] T26;
  wire[26:0] T27;
  wire[25:0] T28;
  wire[25:0] T29;
  wire[24:0] T30;
  wire[24:0] T31;
  wire[23:0] T32;
  wire[23:0] T33;
  wire[22:0] T34;
  wire[22:0] T35;
  wire[21:0] T36;
  wire[21:0] T37;
  wire[20:0] T38;
  wire[20:0] T39;
  wire[19:0] T40;
  wire[19:0] T41;
  wire[18:0] T42;
  wire[18:0] T43;
  wire[17:0] T44;
  wire[17:0] T45;
  wire[16:0] T46;
  wire[16:0] T47;
  wire[15:0] T48;
  wire[15:0] T49;
  wire[14:0] T50;
  wire[14:0] T51;
  wire[13:0] T52;
  wire[13:0] T53;
  wire[12:0] T54;
  wire[12:0] T55;
  wire[11:0] T56;
  wire[11:0] T57;
  wire[10:0] T58;
  wire[10:0] T59;
  wire[9:0] T60;
  wire[9:0] T61;
  wire[8:0] T62;
  wire[8:0] T63;
  wire[7:0] T64;
  wire[7:0] T65;
  wire[6:0] T66;
  wire[6:0] T67;
  wire[5:0] T68;
  wire[5:0] T69;
  wire[4:0] T70;
  wire[4:0] T71;
  wire[3:0] T72;
  wire[3:0] T73;
  wire[2:0] T74;
  wire[2:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire T80;
  wire[3:0] T81;
  wire[3:0] T82;
  wire[3:0] T83;
  wire[9:0] T84;
  wire[9:0] T85;
  wire T86;
  wire T87;
  wire T88;
  wire[3:0] T89;
  wire[3:0] T90;
  wire[3:0] T91;
  wire[9:0] T92;
  wire[9:0] T93;
  wire T94;
  wire T95;
  wire T96;
  wire[3:0] T97;
  wire[3:0] T98;
  wire[3:0] T99;
  wire[9:0] T100;
  wire[9:0] T101;
  wire T102;
  wire T103;
  wire T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[9:0] T108;
  wire[9:0] T109;
  wire T110;
  wire T111;
  wire T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire[9:0] T116;
  wire[9:0] T117;
  wire T118;
  wire T119;
  wire T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[9:0] T124;
  wire[9:0] T125;
  wire T126;
  wire T127;
  wire T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[9:0] T132;
  wire[9:0] T133;
  wire T134;
  wire T135;
  wire T136;
  wire[3:0] T137;
  wire[3:0] T138;
  wire[3:0] T139;
  wire[9:0] T140;
  wire[9:0] T141;
  wire T142;
  wire T143;
  wire T144;
  wire[3:0] T145;
  wire[3:0] T146;
  wire[3:0] T147;
  wire[8:0] T148;
  wire[8:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire[3:0] T153;
  wire[3:0] T154;
  wire[3:0] T155;
  wire[8:0] T156;
  wire[8:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire[3:0] T161;
  wire[3:0] T162;
  wire[3:0] T163;
  wire[8:0] T164;
  wire[8:0] T165;
  wire T166;
  wire T167;
  wire T168;
  wire[3:0] T169;
  wire[3:0] T170;
  wire[3:0] T171;
  wire[8:0] T172;
  wire[8:0] T173;
  wire T174;
  wire T175;
  wire T176;
  wire[3:0] T177;
  wire[3:0] T178;
  wire[3:0] T179;
  wire[8:0] T180;
  wire[8:0] T181;
  wire T182;
  wire T183;
  wire T184;
  wire[3:0] T185;
  wire[3:0] T186;
  wire[3:0] T187;
  wire[8:0] T188;
  wire[8:0] T189;
  wire T190;
  wire T191;
  wire T192;
  wire[3:0] T193;
  wire[3:0] T194;
  wire[3:0] T195;
  wire[8:0] T196;
  wire[8:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire[3:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[8:0] T204;
  wire[8:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire[3:0] T209;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[8:0] T212;
  wire[8:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire[3:0] T219;
  wire[8:0] T220;
  wire[8:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire[3:0] T225;
  wire[3:0] T226;
  wire[3:0] T227;
  wire[8:0] T228;
  wire[8:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire[3:0] T233;
  wire[3:0] T234;
  wire[3:0] T235;
  wire[8:0] T236;
  wire[8:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire[3:0] T241;
  wire[3:0] T242;
  wire[3:0] T243;
  wire[9:0] T244;
  wire[9:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire[3:0] T249;
  wire[3:0] T250;
  wire[3:0] T251;
  wire[9:0] T252;
  wire[9:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire[3:0] T257;
  wire[3:0] T258;
  wire[3:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire[3:0] T265;
  wire[3:0] T266;
  wire[3:0] T267;
  wire[9:0] T268;
  wire[9:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire[3:0] T273;
  wire[3:0] T274;
  wire[3:0] T275;
  wire[9:0] T276;
  wire[9:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[9:0] T284;
  wire[9:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[9:0] T292;
  wire[9:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[9:0] T300;
  wire[9:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[8:0] T308;
  wire[8:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[8:0] T316;
  wire[8:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[8:0] T324;
  wire[8:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[8:0] T332;
  wire[8:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[8:0] T340;
  wire[8:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[8:0] T348;
  wire[8:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[8:0] T356;
  wire[8:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[8:0] T364;
  wire[8:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[8:0] T372;
  wire[8:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[8:0] T380;
  wire[8:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[8:0] T388;
  wire[8:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[8:0] T396;
  wire[8:0] T397;
  wire[7:0] T398;
  wire[7:0] T399;
  wire[6:0] T400;
  wire[6:0] T401;
  wire[5:0] T402;
  wire[5:0] T403;
  wire[4:0] T404;
  wire[4:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire[2:0] T408;
  wire[2:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire T412;
  wire T413;
  wire T414;
  wire[15:0] T415;
  wire[15:0] T416;
  wire[15:0] T417;
  wire[3:0] T418;
  wire[15:0] T419;
  wire[15:0] T420;
  wire T421;
  wire T422;
  wire T423;
  wire[15:0] T424;
  wire[15:0] T425;
  wire[15:0] T426;
  wire[3:0] T427;
  wire[15:0] T428;
  wire[15:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[15:0] T433;
  wire[15:0] T434;
  wire[15:0] T435;
  wire[3:0] T436;
  wire[15:0] T437;
  wire[15:0] T438;
  wire T439;
  wire T440;
  wire T441;
  wire[15:0] T442;
  wire[15:0] T443;
  wire[15:0] T444;
  wire[3:0] T445;
  wire[15:0] T446;
  wire[15:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[15:0] T451;
  wire[15:0] T452;
  wire[15:0] T453;
  wire[3:0] T454;
  wire[15:0] T455;
  wire[15:0] T456;
  wire T457;
  wire T458;
  wire T459;
  wire[15:0] T460;
  wire[15:0] T461;
  wire[15:0] T462;
  wire[3:0] T463;
  wire[15:0] T464;
  wire[15:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire[15:0] T469;
  wire[15:0] T470;
  wire[15:0] T471;
  wire[3:0] T472;
  wire[15:0] T473;
  wire[15:0] T474;
  wire T475;
  wire T476;
  wire T477;
  wire[15:0] T478;
  wire[15:0] T479;
  wire[15:0] T480;
  wire[3:0] T481;
  wire[15:0] T482;
  wire[15:0] T483;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T390, T2};
  assign T2 = T3;
  assign T3 = {T382, T4};
  assign T4 = T5;
  assign T5 = {T374, T6};
  assign T6 = T7;
  assign T7 = {T366, T8};
  assign T8 = T9;
  assign T9 = {T358, T10};
  assign T10 = T11;
  assign T11 = {T350, T12};
  assign T12 = T13;
  assign T13 = {T342, T14};
  assign T14 = T15;
  assign T15 = {T334, T16};
  assign T16 = T17;
  assign T17 = {T326, T18};
  assign T18 = T19;
  assign T19 = {T318, T20};
  assign T20 = T21;
  assign T21 = {T310, T22};
  assign T22 = T23;
  assign T23 = {T302, T24};
  assign T24 = T25;
  assign T25 = {T294, T26};
  assign T26 = T27;
  assign T27 = {T286, T28};
  assign T28 = T29;
  assign T29 = {T278, T30};
  assign T30 = T31;
  assign T31 = {T270, T32};
  assign T32 = T33;
  assign T33 = {T262, T34};
  assign T34 = T35;
  assign T35 = {T254, T36};
  assign T36 = T37;
  assign T37 = {T246, T38};
  assign T38 = T39;
  assign T39 = {T238, T40};
  assign T40 = T41;
  assign T41 = {T230, T42};
  assign T42 = T43;
  assign T43 = {T222, T44};
  assign T44 = T45;
  assign T45 = {T214, T46};
  assign T46 = T47;
  assign T47 = {T206, T48};
  assign T48 = T49;
  assign T49 = {T198, T50};
  assign T50 = T51;
  assign T51 = {T190, T52};
  assign T52 = T53;
  assign T53 = {T182, T54};
  assign T54 = T55;
  assign T55 = {T174, T56};
  assign T56 = T57;
  assign T57 = {T166, T58};
  assign T58 = T59;
  assign T59 = {T158, T60};
  assign T60 = T61;
  assign T61 = {T150, T62};
  assign T62 = T63;
  assign T63 = {T142, T64};
  assign T64 = T65;
  assign T65 = {T134, T66};
  assign T66 = T67;
  assign T67 = {T126, T68};
  assign T68 = T69;
  assign T69 = {T118, T70};
  assign T70 = T71;
  assign T71 = {T110, T72};
  assign T72 = T73;
  assign T73 = {T102, T74};
  assign T74 = T75;
  assign T75 = {T94, T76};
  assign T76 = T77;
  assign T77 = {T86, T78};
  assign T78 = T79;
  assign T79 = T80;
  assign T80 = T84[T81];
  assign T81 = T82;
  assign T82 = T83;
  assign T83 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T84 = T85;
  assign T85 = io_chanxy_in[4'h9/* 9*/:1'h0/* 0*/];
  assign T86 = T87;
  assign T87 = T88;
  assign T88 = T92[T89];
  assign T89 = T90;
  assign T90 = T91;
  assign T91 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T92 = T93;
  assign T93 = io_chanxy_in[5'h13/* 19*/:4'ha/* 10*/];
  assign T94 = T95;
  assign T95 = T96;
  assign T96 = T100[T97];
  assign T97 = T98;
  assign T98 = T99;
  assign T99 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T100 = T101;
  assign T101 = io_chanxy_in[5'h1d/* 29*/:5'h14/* 20*/];
  assign T102 = T103;
  assign T103 = T104;
  assign T104 = T108[T105];
  assign T105 = T106;
  assign T106 = T107;
  assign T107 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T108 = T109;
  assign T109 = io_chanxy_in[6'h27/* 39*/:5'h1e/* 30*/];
  assign T110 = T111;
  assign T111 = T112;
  assign T112 = T116[T113];
  assign T113 = T114;
  assign T114 = T115;
  assign T115 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T116 = T117;
  assign T117 = io_chanxy_in[6'h31/* 49*/:6'h28/* 40*/];
  assign T118 = T119;
  assign T119 = T120;
  assign T120 = T124[T121];
  assign T121 = T122;
  assign T122 = T123;
  assign T123 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T124 = T125;
  assign T125 = io_chanxy_in[6'h3b/* 59*/:6'h32/* 50*/];
  assign T126 = T127;
  assign T127 = T128;
  assign T128 = T132[T129];
  assign T129 = T130;
  assign T130 = T131;
  assign T131 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T132 = T133;
  assign T133 = io_chanxy_in[7'h45/* 69*/:6'h3c/* 60*/];
  assign T134 = T135;
  assign T135 = T136;
  assign T136 = T140[T137];
  assign T137 = T138;
  assign T138 = T139;
  assign T139 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T140 = T141;
  assign T141 = io_chanxy_in[7'h4f/* 79*/:7'h46/* 70*/];
  assign T142 = T143;
  assign T143 = T144;
  assign T144 = T148[T145];
  assign T145 = T146;
  assign T146 = T147;
  assign T147 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T148 = T149;
  assign T149 = io_chanxy_in[7'h58/* 88*/:7'h50/* 80*/];
  assign T150 = T151;
  assign T151 = T152;
  assign T152 = T156[T153];
  assign T153 = T154;
  assign T154 = T155;
  assign T155 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T156 = T157;
  assign T157 = io_chanxy_in[7'h61/* 97*/:7'h59/* 89*/];
  assign T158 = T159;
  assign T159 = T160;
  assign T160 = T164[T161];
  assign T161 = T162;
  assign T162 = T163;
  assign T163 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T164 = T165;
  assign T165 = io_chanxy_in[7'h6a/* 106*/:7'h62/* 98*/];
  assign T166 = T167;
  assign T167 = T168;
  assign T168 = T172[T169];
  assign T169 = T170;
  assign T170 = T171;
  assign T171 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T172 = T173;
  assign T173 = io_chanxy_in[7'h73/* 115*/:7'h6b/* 107*/];
  assign T174 = T175;
  assign T175 = T176;
  assign T176 = T180[T177];
  assign T177 = T178;
  assign T178 = T179;
  assign T179 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T180 = T181;
  assign T181 = io_chanxy_in[7'h7c/* 124*/:7'h74/* 116*/];
  assign T182 = T183;
  assign T183 = T184;
  assign T184 = T188[T185];
  assign T185 = T186;
  assign T186 = T187;
  assign T187 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T188 = T189;
  assign T189 = io_chanxy_in[8'h85/* 133*/:7'h7d/* 125*/];
  assign T190 = T191;
  assign T191 = T192;
  assign T192 = T196[T193];
  assign T193 = T194;
  assign T194 = T195;
  assign T195 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T196 = T197;
  assign T197 = io_chanxy_in[8'h8e/* 142*/:8'h86/* 134*/];
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[8'h97/* 151*/:8'h8f/* 143*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[8'ha0/* 160*/:8'h98/* 152*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[8'ha9/* 169*/:8'ha1/* 161*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[8'hb2/* 178*/:8'haa/* 170*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[8'hbb/* 187*/:8'hb3/* 179*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[8'hc5/* 197*/:8'hbc/* 188*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[8'hcf/* 207*/:8'hc6/* 198*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[8'hd9/* 217*/:8'hd0/* 208*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[8'he3/* 227*/:8'hda/* 218*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[8'hed/* 237*/:8'he4/* 228*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[8'hf7/* 247*/:8'hee/* 238*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[9'h101/* 257*/:8'hf8/* 248*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[9'h10b/* 267*/:9'h102/* 258*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[9'h114/* 276*/:9'h10c/* 268*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[9'h11d/* 285*/:9'h115/* 277*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[9'h126/* 294*/:9'h11e/* 286*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[9'h12f/* 303*/:9'h127/* 295*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[9'h138/* 312*/:9'h130/* 304*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[9'h141/* 321*/:9'h139/* 313*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[9'h14a/* 330*/:9'h142/* 322*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[9'h153/* 339*/:9'h14b/* 331*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[9'h15c/* 348*/:9'h154/* 340*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[9'h165/* 357*/:9'h15d/* 349*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[9'h16e/* 366*/:9'h166/* 358*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[9'h177/* 375*/:9'h16f/* 367*/];
  assign io_ipin_out = T398;
  assign T398 = T399;
  assign T399 = {T475, T400};
  assign T400 = T401;
  assign T401 = {T466, T402};
  assign T402 = T403;
  assign T403 = {T457, T404};
  assign T404 = T405;
  assign T405 = {T448, T406};
  assign T406 = T407;
  assign T407 = {T439, T408};
  assign T408 = T409;
  assign T409 = {T430, T410};
  assign T410 = T411;
  assign T411 = {T421, T412};
  assign T412 = T413;
  assign T413 = T414;
  assign T414 = T419[T415];
  assign T415 = T416;
  assign T416 = T417;
  assign T417 = {12'h0/* 0*/, T418};
  assign T418 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T419 = T420;
  assign T420 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = T428[T424];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = {12'h0/* 0*/, T427};
  assign T427 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T428 = T429;
  assign T429 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T437[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = {12'h0/* 0*/, T436};
  assign T436 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T437 = T438;
  assign T438 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T439 = T440;
  assign T440 = T441;
  assign T441 = T446[T442];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = {12'h0/* 0*/, T445};
  assign T445 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T446 = T447;
  assign T447 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T455[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = {12'h0/* 0*/, T454};
  assign T454 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T455 = T456;
  assign T456 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = T464[T460];
  assign T460 = T461;
  assign T461 = T462;
  assign T462 = {12'h0/* 0*/, T463};
  assign T463 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T464 = T465;
  assign T465 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T473[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = {12'h0/* 0*/, T472};
  assign T472 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T473 = T474;
  assign T474 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = T482[T478];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = {12'h0/* 0*/, T481};
  assign T481 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T482 = T483;
  assign T483 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule

module io_tile_sp_11(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [375:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_x_loc = T3;
  assign T3 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_12(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [375:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_x_loc = T3;
  assign T3 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_13(input clk, input reset,
    input [31:0] io_configs_in,
    input [5:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [375:0] io_chanxy_in,
    output[39:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[159:0] T0;
  wire[191:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[39:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hbf/* 191*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_x_loc = T3;
  assign T3 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_6 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_sbcb_wc_5(
    input [127:0] io_ipin_in,
    input [31:0] io_ipin_config,
    input [355:0] io_chanxy_in,
    input [167:0] io_chanxy_config,
    output[7:0] io_ipin_out,
    output[99:0] io_chanxy_out);

  wire[99:0] T0;
  wire[99:0] T1;
  wire[98:0] T2;
  wire[98:0] T3;
  wire[97:0] T4;
  wire[97:0] T5;
  wire[96:0] T6;
  wire[96:0] T7;
  wire[95:0] T8;
  wire[95:0] T9;
  wire[94:0] T10;
  wire[94:0] T11;
  wire[93:0] T12;
  wire[93:0] T13;
  wire[92:0] T14;
  wire[92:0] T15;
  wire[91:0] T16;
  wire[91:0] T17;
  wire[90:0] T18;
  wire[90:0] T19;
  wire[89:0] T20;
  wire[89:0] T21;
  wire[88:0] T22;
  wire[88:0] T23;
  wire[87:0] T24;
  wire[87:0] T25;
  wire[86:0] T26;
  wire[86:0] T27;
  wire[85:0] T28;
  wire[85:0] T29;
  wire[84:0] T30;
  wire[84:0] T31;
  wire[83:0] T32;
  wire[83:0] T33;
  wire[82:0] T34;
  wire[82:0] T35;
  wire[81:0] T36;
  wire[81:0] T37;
  wire[80:0] T38;
  wire[80:0] T39;
  wire[79:0] T40;
  wire[79:0] T41;
  wire[78:0] T42;
  wire[78:0] T43;
  wire[77:0] T44;
  wire[77:0] T45;
  wire[76:0] T46;
  wire[76:0] T47;
  wire[75:0] T48;
  wire[75:0] T49;
  wire[74:0] T50;
  wire[74:0] T51;
  wire[73:0] T52;
  wire[73:0] T53;
  wire[72:0] T54;
  wire[72:0] T55;
  wire[71:0] T56;
  wire[71:0] T57;
  wire[70:0] T58;
  wire[70:0] T59;
  wire[69:0] T60;
  wire[69:0] T61;
  wire[68:0] T62;
  wire[68:0] T63;
  wire[67:0] T64;
  wire[67:0] T65;
  wire[66:0] T66;
  wire[66:0] T67;
  wire[65:0] T68;
  wire[65:0] T69;
  wire[64:0] T70;
  wire[64:0] T71;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[62:0] T74;
  wire[62:0] T75;
  wire[61:0] T76;
  wire[61:0] T77;
  wire[60:0] T78;
  wire[60:0] T79;
  wire[59:0] T80;
  wire[59:0] T81;
  wire[58:0] T82;
  wire[58:0] T83;
  wire[57:0] T84;
  wire[57:0] T85;
  wire[56:0] T86;
  wire[56:0] T87;
  wire[55:0] T88;
  wire[55:0] T89;
  wire[54:0] T90;
  wire[54:0] T91;
  wire[53:0] T92;
  wire[53:0] T93;
  wire[52:0] T94;
  wire[52:0] T95;
  wire[51:0] T96;
  wire[51:0] T97;
  wire[50:0] T98;
  wire[50:0] T99;
  wire[49:0] T100;
  wire[49:0] T101;
  wire[48:0] T102;
  wire[48:0] T103;
  wire[47:0] T104;
  wire[47:0] T105;
  wire[46:0] T106;
  wire[46:0] T107;
  wire[45:0] T108;
  wire[45:0] T109;
  wire[44:0] T110;
  wire[44:0] T111;
  wire[43:0] T112;
  wire[43:0] T113;
  wire[42:0] T114;
  wire[42:0] T115;
  wire[41:0] T116;
  wire[41:0] T117;
  wire[40:0] T118;
  wire[40:0] T119;
  wire[39:0] T120;
  wire[39:0] T121;
  wire[38:0] T122;
  wire[38:0] T123;
  wire[37:0] T124;
  wire[37:0] T125;
  wire[36:0] T126;
  wire[36:0] T127;
  wire[35:0] T128;
  wire[35:0] T129;
  wire[34:0] T130;
  wire[34:0] T131;
  wire[33:0] T132;
  wire[33:0] T133;
  wire[32:0] T134;
  wire[32:0] T135;
  wire[31:0] T136;
  wire[31:0] T137;
  wire[30:0] T138;
  wire[30:0] T139;
  wire[29:0] T140;
  wire[29:0] T141;
  wire[28:0] T142;
  wire[28:0] T143;
  wire[27:0] T144;
  wire[27:0] T145;
  wire[26:0] T146;
  wire[26:0] T147;
  wire[25:0] T148;
  wire[25:0] T149;
  wire[24:0] T150;
  wire[24:0] T151;
  wire[23:0] T152;
  wire[23:0] T153;
  wire[22:0] T154;
  wire[22:0] T155;
  wire[21:0] T156;
  wire[21:0] T157;
  wire[20:0] T158;
  wire[20:0] T159;
  wire[19:0] T160;
  wire[19:0] T161;
  wire[18:0] T162;
  wire[18:0] T163;
  wire[17:0] T164;
  wire[17:0] T165;
  wire[16:0] T166;
  wire[16:0] T167;
  wire[15:0] T168;
  wire[15:0] T169;
  wire[14:0] T170;
  wire[14:0] T171;
  wire[13:0] T172;
  wire[13:0] T173;
  wire[12:0] T174;
  wire[12:0] T175;
  wire[11:0] T176;
  wire[11:0] T177;
  wire[10:0] T178;
  wire[10:0] T179;
  wire[9:0] T180;
  wire[9:0] T181;
  wire[8:0] T182;
  wire[8:0] T183;
  wire[7:0] T184;
  wire[7:0] T185;
  wire[6:0] T186;
  wire[6:0] T187;
  wire[5:0] T188;
  wire[5:0] T189;
  wire[4:0] T190;
  wire[4:0] T191;
  wire[3:0] T192;
  wire[3:0] T193;
  wire[2:0] T194;
  wire[2:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire[1:0] T201;
  wire[1:0] T202;
  wire[1:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire T206;
  wire T207;
  wire T208;
  wire[1:0] T209;
  wire[1:0] T210;
  wire[1:0] T211;
  wire[2:0] T212;
  wire[2:0] T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire[1:0] T260;
  wire[1:0] T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[1:0] T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[2:0] T364;
  wire[2:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[2:0] T372;
  wire[2:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire[1:0] T523;
  wire[2:0] T524;
  wire[2:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[1:0] T529;
  wire[1:0] T530;
  wire[1:0] T531;
  wire[2:0] T532;
  wire[2:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[3:0] T681;
  wire[3:0] T682;
  wire[3:0] T683;
  wire[9:0] T684;
  wire[9:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[1:0] T689;
  wire[1:0] T690;
  wire[1:0] T691;
  wire[2:0] T692;
  wire[2:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[9:0] T700;
  wire[9:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[1:0] T705;
  wire[1:0] T706;
  wire[1:0] T707;
  wire[2:0] T708;
  wire[2:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[3:0] T713;
  wire[3:0] T714;
  wire[3:0] T715;
  wire[9:0] T716;
  wire[9:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[3:0] T729;
  wire[3:0] T730;
  wire[3:0] T731;
  wire[9:0] T732;
  wire[9:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[3:0] T745;
  wire[3:0] T746;
  wire[3:0] T747;
  wire[9:0] T748;
  wire[9:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire[9:0] T764;
  wire[9:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[9:0] T780;
  wire[9:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[3:0] T793;
  wire[3:0] T794;
  wire[3:0] T795;
  wire[9:0] T796;
  wire[9:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[3:0] T809;
  wire[3:0] T810;
  wire[3:0] T811;
  wire[8:0] T812;
  wire[8:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[8:0] T828;
  wire[8:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[3:0] T841;
  wire[3:0] T842;
  wire[3:0] T843;
  wire[8:0] T844;
  wire[8:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[8:0] T860;
  wire[8:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T875;
  wire[8:0] T876;
  wire[8:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[3:0] T890;
  wire[3:0] T891;
  wire[8:0] T892;
  wire[8:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[3:0] T905;
  wire[3:0] T906;
  wire[3:0] T907;
  wire[8:0] T908;
  wire[8:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[3:0] T921;
  wire[3:0] T922;
  wire[3:0] T923;
  wire[8:0] T924;
  wire[8:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[8:0] T940;
  wire[8:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[3:0] T953;
  wire[3:0] T954;
  wire[3:0] T955;
  wire[8:0] T956;
  wire[8:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[3:0] T969;
  wire[3:0] T970;
  wire[3:0] T971;
  wire[8:0] T972;
  wire[8:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[3:0] T985;
  wire[3:0] T986;
  wire[3:0] T987;
  wire[8:0] T988;
  wire[8:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire[7:0] T998;
  wire[7:0] T999;
  wire[6:0] T1000;
  wire[6:0] T1001;
  wire[5:0] T1002;
  wire[5:0] T1003;
  wire[4:0] T1004;
  wire[4:0] T1005;
  wire[3:0] T1006;
  wire[3:0] T1007;
  wire[2:0] T1008;
  wire[2:0] T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire[15:0] T1015;
  wire[15:0] T1016;
  wire[15:0] T1017;
  wire[3:0] T1018;
  wire[15:0] T1019;
  wire[15:0] T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[15:0] T1024;
  wire[15:0] T1025;
  wire[15:0] T1026;
  wire[3:0] T1027;
  wire[15:0] T1028;
  wire[15:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[15:0] T1033;
  wire[15:0] T1034;
  wire[15:0] T1035;
  wire[3:0] T1036;
  wire[15:0] T1037;
  wire[15:0] T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire[15:0] T1042;
  wire[15:0] T1043;
  wire[15:0] T1044;
  wire[3:0] T1045;
  wire[15:0] T1046;
  wire[15:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire[15:0] T1051;
  wire[15:0] T1052;
  wire[15:0] T1053;
  wire[3:0] T1054;
  wire[15:0] T1055;
  wire[15:0] T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[15:0] T1060;
  wire[15:0] T1061;
  wire[15:0] T1062;
  wire[3:0] T1063;
  wire[15:0] T1064;
  wire[15:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[15:0] T1069;
  wire[15:0] T1070;
  wire[15:0] T1071;
  wire[3:0] T1072;
  wire[15:0] T1073;
  wire[15:0] T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire[15:0] T1078;
  wire[15:0] T1079;
  wire[15:0] T1080;
  wire[3:0] T1081;
  wire[15:0] T1082;
  wire[15:0] T1083;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T990, T2};
  assign T2 = T3;
  assign T3 = {T982, T4};
  assign T4 = T5;
  assign T5 = {T974, T6};
  assign T6 = T7;
  assign T7 = {T966, T8};
  assign T8 = T9;
  assign T9 = {T958, T10};
  assign T10 = T11;
  assign T11 = {T950, T12};
  assign T12 = T13;
  assign T13 = {T942, T14};
  assign T14 = T15;
  assign T15 = {T934, T16};
  assign T16 = T17;
  assign T17 = {T926, T18};
  assign T18 = T19;
  assign T19 = {T918, T20};
  assign T20 = T21;
  assign T21 = {T910, T22};
  assign T22 = T23;
  assign T23 = {T902, T24};
  assign T24 = T25;
  assign T25 = {T894, T26};
  assign T26 = T27;
  assign T27 = {T886, T28};
  assign T28 = T29;
  assign T29 = {T878, T30};
  assign T30 = T31;
  assign T31 = {T870, T32};
  assign T32 = T33;
  assign T33 = {T862, T34};
  assign T34 = T35;
  assign T35 = {T854, T36};
  assign T36 = T37;
  assign T37 = {T846, T38};
  assign T38 = T39;
  assign T39 = {T838, T40};
  assign T40 = T41;
  assign T41 = {T830, T42};
  assign T42 = T43;
  assign T43 = {T822, T44};
  assign T44 = T45;
  assign T45 = {T814, T46};
  assign T46 = T47;
  assign T47 = {T806, T48};
  assign T48 = T49;
  assign T49 = {T798, T50};
  assign T50 = T51;
  assign T51 = {T790, T52};
  assign T52 = T53;
  assign T53 = {T782, T54};
  assign T54 = T55;
  assign T55 = {T774, T56};
  assign T56 = T57;
  assign T57 = {T766, T58};
  assign T58 = T59;
  assign T59 = {T758, T60};
  assign T60 = T61;
  assign T61 = {T750, T62};
  assign T62 = T63;
  assign T63 = {T742, T64};
  assign T64 = T65;
  assign T65 = {T734, T66};
  assign T66 = T67;
  assign T67 = {T726, T68};
  assign T68 = T69;
  assign T69 = {T718, T70};
  assign T70 = T71;
  assign T71 = {T710, T72};
  assign T72 = T73;
  assign T73 = {T702, T74};
  assign T74 = T75;
  assign T75 = {T694, T76};
  assign T76 = T77;
  assign T77 = {T686, T78};
  assign T78 = T79;
  assign T79 = {T678, T80};
  assign T80 = T81;
  assign T81 = {T670, T82};
  assign T82 = T83;
  assign T83 = {T662, T84};
  assign T84 = T85;
  assign T85 = {T654, T86};
  assign T86 = T87;
  assign T87 = {T646, T88};
  assign T88 = T89;
  assign T89 = {T638, T90};
  assign T90 = T91;
  assign T91 = {T630, T92};
  assign T92 = T93;
  assign T93 = {T622, T94};
  assign T94 = T95;
  assign T95 = {T614, T96};
  assign T96 = T97;
  assign T97 = {T606, T98};
  assign T98 = T99;
  assign T99 = {T598, T100};
  assign T100 = T101;
  assign T101 = {T590, T102};
  assign T102 = T103;
  assign T103 = {T582, T104};
  assign T104 = T105;
  assign T105 = {T574, T106};
  assign T106 = T107;
  assign T107 = {T566, T108};
  assign T108 = T109;
  assign T109 = {T558, T110};
  assign T110 = T111;
  assign T111 = {T550, T112};
  assign T112 = T113;
  assign T113 = {T542, T114};
  assign T114 = T115;
  assign T115 = {T534, T116};
  assign T116 = T117;
  assign T117 = {T526, T118};
  assign T118 = T119;
  assign T119 = {T518, T120};
  assign T120 = T121;
  assign T121 = {T510, T122};
  assign T122 = T123;
  assign T123 = {T502, T124};
  assign T124 = T125;
  assign T125 = {T494, T126};
  assign T126 = T127;
  assign T127 = {T486, T128};
  assign T128 = T129;
  assign T129 = {T478, T130};
  assign T130 = T131;
  assign T131 = {T470, T132};
  assign T132 = T133;
  assign T133 = {T462, T134};
  assign T134 = T135;
  assign T135 = {T454, T136};
  assign T136 = T137;
  assign T137 = {T446, T138};
  assign T138 = T139;
  assign T139 = {T438, T140};
  assign T140 = T141;
  assign T141 = {T430, T142};
  assign T142 = T143;
  assign T143 = {T422, T144};
  assign T144 = T145;
  assign T145 = {T414, T146};
  assign T146 = T147;
  assign T147 = {T406, T148};
  assign T148 = T149;
  assign T149 = {T398, T150};
  assign T150 = T151;
  assign T151 = {T390, T152};
  assign T152 = T153;
  assign T153 = {T382, T154};
  assign T154 = T155;
  assign T155 = {T374, T156};
  assign T156 = T157;
  assign T157 = {T366, T158};
  assign T158 = T159;
  assign T159 = {T358, T160};
  assign T160 = T161;
  assign T161 = {T350, T162};
  assign T162 = T163;
  assign T163 = {T342, T164};
  assign T164 = T165;
  assign T165 = {T334, T166};
  assign T166 = T167;
  assign T167 = {T326, T168};
  assign T168 = T169;
  assign T169 = {T318, T170};
  assign T170 = T171;
  assign T171 = {T310, T172};
  assign T172 = T173;
  assign T173 = {T302, T174};
  assign T174 = T175;
  assign T175 = {T294, T176};
  assign T176 = T177;
  assign T177 = {T286, T178};
  assign T178 = T179;
  assign T179 = {T278, T180};
  assign T180 = T181;
  assign T181 = {T270, T182};
  assign T182 = T183;
  assign T183 = {T262, T184};
  assign T184 = T185;
  assign T185 = {T254, T186};
  assign T186 = T187;
  assign T187 = {T246, T188};
  assign T188 = T189;
  assign T189 = {T238, T190};
  assign T190 = T191;
  assign T191 = {T230, T192};
  assign T192 = T193;
  assign T193 = {T222, T194};
  assign T194 = T195;
  assign T195 = {T214, T196};
  assign T196 = T197;
  assign T197 = {T206, T198};
  assign T198 = T199;
  assign T199 = T200;
  assign T200 = T204[T201];
  assign T201 = T202;
  assign T202 = T203;
  assign T203 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T204 = T205;
  assign T205 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T206 = T207;
  assign T207 = T208;
  assign T208 = T212[T209];
  assign T209 = T210;
  assign T210 = T211;
  assign T211 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T212 = T213;
  assign T213 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T214 = T215;
  assign T215 = T216;
  assign T216 = T220[T217];
  assign T217 = T218;
  assign T218 = T219;
  assign T219 = io_chanxy_config[3'h4/* 4*/:3'h4/* 4*/];
  assign T220 = T221;
  assign T221 = io_chanxy_in[3'h7/* 7*/:3'h6/* 6*/];
  assign T222 = T223;
  assign T223 = T224;
  assign T224 = T228[T225];
  assign T225 = T226;
  assign T226 = T227;
  assign T227 = io_chanxy_config[3'h5/* 5*/:3'h5/* 5*/];
  assign T228 = T229;
  assign T229 = io_chanxy_in[4'h9/* 9*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = T232;
  assign T232 = T236[T233];
  assign T233 = T234;
  assign T234 = T235;
  assign T235 = io_chanxy_config[3'h6/* 6*/:3'h6/* 6*/];
  assign T236 = T237;
  assign T237 = io_chanxy_in[4'hb/* 11*/:4'ha/* 10*/];
  assign T238 = T239;
  assign T239 = T240;
  assign T240 = T244[T241];
  assign T241 = T242;
  assign T242 = T243;
  assign T243 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T244 = T245;
  assign T245 = io_chanxy_in[4'hd/* 13*/:4'hc/* 12*/];
  assign T246 = T247;
  assign T247 = T248;
  assign T248 = T252[T249];
  assign T249 = T250;
  assign T250 = T251;
  assign T251 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T252 = T253;
  assign T253 = io_chanxy_in[4'hf/* 15*/:4'he/* 14*/];
  assign T254 = T255;
  assign T255 = T256;
  assign T256 = T260[T257];
  assign T257 = T258;
  assign T258 = T259;
  assign T259 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T260 = T261;
  assign T261 = io_chanxy_in[5'h11/* 17*/:5'h10/* 16*/];
  assign T262 = T263;
  assign T263 = T264;
  assign T264 = T268[T265];
  assign T265 = T266;
  assign T266 = T267;
  assign T267 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T268 = T269;
  assign T269 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T270 = T271;
  assign T271 = T272;
  assign T272 = T276[T273];
  assign T273 = T274;
  assign T274 = T275;
  assign T275 = io_chanxy_config[4'hb/* 11*/:4'hb/* 11*/];
  assign T276 = T277;
  assign T277 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[6'h2c/* 44*/:6'h2a/* 42*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h2f/* 47*/:6'h2d/* 45*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[6'h33/* 51*/:6'h32/* 50*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[6'h35/* 53*/:6'h34/* 52*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[6'h2b/* 43*/:6'h2b/* 43*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[7'h56/* 86*/:7'h54/* 84*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[7'h59/* 89*/:7'h57/* 87*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h34/* 52*/:6'h34/* 52*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h35/* 53*/:6'h35/* 53*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[7'h71/* 113*/:7'h70/* 112*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[6'h3c/* 60*/:6'h3c/* 60*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[7'h73/* 115*/:7'h72/* 114*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[6'h3d/* 61*/:6'h3d/* 61*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[7'h75/* 117*/:7'h74/* 116*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[6'h3e/* 62*/:6'h3e/* 62*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[7'h77/* 119*/:7'h76/* 118*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[6'h3f/* 63*/:6'h3f/* 63*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h79/* 121*/:7'h78/* 120*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h41/* 65*/:7'h41/* 65*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'h87/* 135*/:7'h7e/* 126*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'h8a/* 138*/:8'h88/* 136*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'h94/* 148*/:8'h8b/* 139*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'h97/* 151*/:8'h95/* 149*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h51/* 81*/:7'h4e/* 78*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'ha1/* 161*/:8'h98/* 152*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h56/* 86*/:7'h53/* 83*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'had/* 173*/:8'ha4/* 164*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'hb9/* 185*/:8'hb0/* 176*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h5c/* 92*/:7'h5c/* 92*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'hbb/* 187*/:8'hba/* 186*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h60/* 96*/:7'h5d/* 93*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'hc5/* 197*/:8'hbc/* 188*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h65/* 101*/:7'h62/* 98*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'hd1/* 209*/:8'hc8/* 200*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h66/* 102*/:7'h66/* 102*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h6a/* 106*/:7'h67/* 103*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'hdd/* 221*/:8'hd4/* 212*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h6b/* 107*/:7'h6b/* 107*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'hdf/* 223*/:8'hde/* 222*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'he8/* 232*/:8'he0/* 224*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h74/* 116*/:7'h71/* 113*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'hf3/* 243*/:8'heb/* 235*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h75/* 117*/:7'h75/* 117*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'hf5/* 245*/:8'hf4/* 244*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[7'h79/* 121*/:7'h76/* 118*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'hfe/* 254*/:8'hf6/* 246*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[7'h7e/* 126*/:7'h7b/* 123*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h109/* 265*/:9'h101/* 257*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h114/* 276*/:9'h10c/* 268*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'h84/* 132*/:8'h84/* 132*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h116/* 278*/:9'h115/* 277*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h88/* 136*/:8'h85/* 133*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h11f/* 287*/:9'h117/* 279*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h121/* 289*/:9'h120/* 288*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h12a/* 298*/:9'h122/* 290*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h12c/* 300*/:9'h12b/* 299*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h92/* 146*/:8'h8f/* 143*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h135/* 309*/:9'h12d/* 301*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h93/* 147*/:8'h93/* 147*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h137/* 311*/:9'h136/* 310*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h140/* 320*/:9'h138/* 312*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'h9c/* 156*/:8'h99/* 153*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h14b/* 331*/:9'h143/* 323*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'h9d/* 157*/:8'h9d/* 157*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h14d/* 333*/:9'h14c/* 332*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'ha1/* 161*/:8'h9e/* 158*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h156/* 342*/:9'h14e/* 334*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'ha2/* 162*/:8'ha2/* 162*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h158/* 344*/:9'h157/* 343*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'ha6/* 166*/:8'ha3/* 163*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h161/* 353*/:9'h159/* 345*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h163/* 355*/:9'h162/* 354*/];
  assign io_ipin_out = T998;
  assign T998 = T999;
  assign T999 = {T1075, T1000};
  assign T1000 = T1001;
  assign T1001 = {T1066, T1002};
  assign T1002 = T1003;
  assign T1003 = {T1057, T1004};
  assign T1004 = T1005;
  assign T1005 = {T1048, T1006};
  assign T1006 = T1007;
  assign T1007 = {T1039, T1008};
  assign T1008 = T1009;
  assign T1009 = {T1030, T1010};
  assign T1010 = T1011;
  assign T1011 = {T1021, T1012};
  assign T1012 = T1013;
  assign T1013 = T1014;
  assign T1014 = T1019[T1015];
  assign T1015 = T1016;
  assign T1016 = T1017;
  assign T1017 = {12'h0/* 0*/, T1018};
  assign T1018 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1019 = T1020;
  assign T1020 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = T1028[T1024];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = {12'h0/* 0*/, T1027};
  assign T1027 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1028 = T1029;
  assign T1029 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1037[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = {12'h0/* 0*/, T1036};
  assign T1036 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1037 = T1038;
  assign T1038 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1039 = T1040;
  assign T1040 = T1041;
  assign T1041 = T1046[T1042];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = {12'h0/* 0*/, T1045};
  assign T1045 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1046 = T1047;
  assign T1047 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1048 = T1049;
  assign T1049 = T1050;
  assign T1050 = T1055[T1051];
  assign T1051 = T1052;
  assign T1052 = T1053;
  assign T1053 = {12'h0/* 0*/, T1054};
  assign T1054 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1055 = T1056;
  assign T1056 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = T1064[T1060];
  assign T1060 = T1061;
  assign T1061 = T1062;
  assign T1062 = {12'h0/* 0*/, T1063};
  assign T1063 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1064 = T1065;
  assign T1065 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1073[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = {12'h0/* 0*/, T1072};
  assign T1072 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1073 = T1074;
  assign T1074 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1075 = T1076;
  assign T1076 = T1077;
  assign T1077 = T1082[T1078];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = {12'h0/* 0*/, T1081};
  assign T1081 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1082 = T1083;
  assign T1083 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
endmodule

module io_tile_sp_14(input clk, input reset,
    input [31:0] io_configs_in,
    input [6:0] io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    input [355:0] io_chanxy_in,
    output[99:0] io_chanxy_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[167:0] T0;
  wire[223:0] this_config_io_configs_out;
  wire[31:0] T1;
  wire[7:0] T2;
  wire[7:0] T3;
  wire[99:0] this_sbcb_io_chanxy_out;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[8'hc7/* 199*/:6'h20/* 32*/];
  assign T1 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h0/* 0*/};
  assign io_x_loc = T3;
  assign T3 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_wc_5 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
    configs_latches_7 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_15(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T2;
  assign T2 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_16(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T2;
  assign T2 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_17(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T2;
  assign T2 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_18(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule

module io_tile_sp_19(input clk, input reset,
    input [31:0] io_configs_in,
    input  io_configs_en,
    input [7:0] io_io_input,
    output[7:0] io_io_output,
    output[7:0] io_opin_out,
    input [127:0] io_ipin_in,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[31:0] T0;
  wire[31:0] this_config_io_configs_out;
  wire[7:0] T1;
  wire[7:0] T2;
  wire[7:0] this_sbcb_io_ipin_out;

  assign T0 = this_config_io_configs_out[5'h1f/* 31*/:1'h0/* 0*/];
  assign io_y_loc = T1;
  assign T1 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T2;
  assign T2 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = io_io_input;
  assign io_io_output = this_sbcb_io_ipin_out;
  io_sbcb_woc this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ));
    configs_latches_1 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
endmodule


