



module sbcb_sp(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [605:0] io_chanxy_in,
    input [287:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[149:0] io_chanxy_out);

  wire[149:0] T0;
  wire[149:0] T1;
  wire[148:0] T2;
  wire[148:0] T3;
  wire[147:0] T4;
  wire[147:0] T5;
  wire[146:0] T6;
  wire[146:0] T7;
  wire[145:0] T8;
  wire[145:0] T9;
  wire[144:0] T10;
  wire[144:0] T11;
  wire[143:0] T12;
  wire[143:0] T13;
  wire[142:0] T14;
  wire[142:0] T15;
  wire[141:0] T16;
  wire[141:0] T17;
  wire[140:0] T18;
  wire[140:0] T19;
  wire[139:0] T20;
  wire[139:0] T21;
  wire[138:0] T22;
  wire[138:0] T23;
  wire[137:0] T24;
  wire[137:0] T25;
  wire[136:0] T26;
  wire[136:0] T27;
  wire[135:0] T28;
  wire[135:0] T29;
  wire[134:0] T30;
  wire[134:0] T31;
  wire[133:0] T32;
  wire[133:0] T33;
  wire[132:0] T34;
  wire[132:0] T35;
  wire[131:0] T36;
  wire[131:0] T37;
  wire[130:0] T38;
  wire[130:0] T39;
  wire[129:0] T40;
  wire[129:0] T41;
  wire[128:0] T42;
  wire[128:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[126:0] T46;
  wire[126:0] T47;
  wire[125:0] T48;
  wire[125:0] T49;
  wire[124:0] T50;
  wire[124:0] T51;
  wire[123:0] T52;
  wire[123:0] T53;
  wire[122:0] T54;
  wire[122:0] T55;
  wire[121:0] T56;
  wire[121:0] T57;
  wire[120:0] T58;
  wire[120:0] T59;
  wire[119:0] T60;
  wire[119:0] T61;
  wire[118:0] T62;
  wire[118:0] T63;
  wire[117:0] T64;
  wire[117:0] T65;
  wire[116:0] T66;
  wire[116:0] T67;
  wire[115:0] T68;
  wire[115:0] T69;
  wire[114:0] T70;
  wire[114:0] T71;
  wire[113:0] T72;
  wire[113:0] T73;
  wire[112:0] T74;
  wire[112:0] T75;
  wire[111:0] T76;
  wire[111:0] T77;
  wire[110:0] T78;
  wire[110:0] T79;
  wire[109:0] T80;
  wire[109:0] T81;
  wire[108:0] T82;
  wire[108:0] T83;
  wire[107:0] T84;
  wire[107:0] T85;
  wire[106:0] T86;
  wire[106:0] T87;
  wire[105:0] T88;
  wire[105:0] T89;
  wire[104:0] T90;
  wire[104:0] T91;
  wire[103:0] T92;
  wire[103:0] T93;
  wire[102:0] T94;
  wire[102:0] T95;
  wire[101:0] T96;
  wire[101:0] T97;
  wire[100:0] T98;
  wire[100:0] T99;
  wire[99:0] T100;
  wire[99:0] T101;
  wire[98:0] T102;
  wire[98:0] T103;
  wire[97:0] T104;
  wire[97:0] T105;
  wire[96:0] T106;
  wire[96:0] T107;
  wire[95:0] T108;
  wire[95:0] T109;
  wire[94:0] T110;
  wire[94:0] T111;
  wire[93:0] T112;
  wire[93:0] T113;
  wire[92:0] T114;
  wire[92:0] T115;
  wire[91:0] T116;
  wire[91:0] T117;
  wire[90:0] T118;
  wire[90:0] T119;
  wire[89:0] T120;
  wire[89:0] T121;
  wire[88:0] T122;
  wire[88:0] T123;
  wire[87:0] T124;
  wire[87:0] T125;
  wire[86:0] T126;
  wire[86:0] T127;
  wire[85:0] T128;
  wire[85:0] T129;
  wire[84:0] T130;
  wire[84:0] T131;
  wire[83:0] T132;
  wire[83:0] T133;
  wire[82:0] T134;
  wire[82:0] T135;
  wire[81:0] T136;
  wire[81:0] T137;
  wire[80:0] T138;
  wire[80:0] T139;
  wire[79:0] T140;
  wire[79:0] T141;
  wire[78:0] T142;
  wire[78:0] T143;
  wire[77:0] T144;
  wire[77:0] T145;
  wire[76:0] T146;
  wire[76:0] T147;
  wire[75:0] T148;
  wire[75:0] T149;
  wire[74:0] T150;
  wire[74:0] T151;
  wire[73:0] T152;
  wire[73:0] T153;
  wire[72:0] T154;
  wire[72:0] T155;
  wire[71:0] T156;
  wire[71:0] T157;
  wire[70:0] T158;
  wire[70:0] T159;
  wire[69:0] T160;
  wire[69:0] T161;
  wire[68:0] T162;
  wire[68:0] T163;
  wire[67:0] T164;
  wire[67:0] T165;
  wire[66:0] T166;
  wire[66:0] T167;
  wire[65:0] T168;
  wire[65:0] T169;
  wire[64:0] T170;
  wire[64:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[62:0] T174;
  wire[62:0] T175;
  wire[61:0] T176;
  wire[61:0] T177;
  wire[60:0] T178;
  wire[60:0] T179;
  wire[59:0] T180;
  wire[59:0] T181;
  wire[58:0] T182;
  wire[58:0] T183;
  wire[57:0] T184;
  wire[57:0] T185;
  wire[56:0] T186;
  wire[56:0] T187;
  wire[55:0] T188;
  wire[55:0] T189;
  wire[54:0] T190;
  wire[54:0] T191;
  wire[53:0] T192;
  wire[53:0] T193;
  wire[52:0] T194;
  wire[52:0] T195;
  wire[51:0] T196;
  wire[51:0] T197;
  wire[50:0] T198;
  wire[50:0] T199;
  wire[49:0] T200;
  wire[49:0] T201;
  wire[48:0] T202;
  wire[48:0] T203;
  wire[47:0] T204;
  wire[47:0] T205;
  wire[46:0] T206;
  wire[46:0] T207;
  wire[45:0] T208;
  wire[45:0] T209;
  wire[44:0] T210;
  wire[44:0] T211;
  wire[43:0] T212;
  wire[43:0] T213;
  wire[42:0] T214;
  wire[42:0] T215;
  wire[41:0] T216;
  wire[41:0] T217;
  wire[40:0] T218;
  wire[40:0] T219;
  wire[39:0] T220;
  wire[39:0] T221;
  wire[38:0] T222;
  wire[38:0] T223;
  wire[37:0] T224;
  wire[37:0] T225;
  wire[36:0] T226;
  wire[36:0] T227;
  wire[35:0] T228;
  wire[35:0] T229;
  wire[34:0] T230;
  wire[34:0] T231;
  wire[33:0] T232;
  wire[33:0] T233;
  wire[32:0] T234;
  wire[32:0] T235;
  wire[31:0] T236;
  wire[31:0] T237;
  wire[30:0] T238;
  wire[30:0] T239;
  wire[29:0] T240;
  wire[29:0] T241;
  wire[28:0] T242;
  wire[28:0] T243;
  wire[27:0] T244;
  wire[27:0] T245;
  wire[26:0] T246;
  wire[26:0] T247;
  wire[25:0] T248;
  wire[25:0] T249;
  wire[24:0] T250;
  wire[24:0] T251;
  wire[23:0] T252;
  wire[23:0] T253;
  wire[22:0] T254;
  wire[22:0] T255;
  wire[21:0] T256;
  wire[21:0] T257;
  wire[20:0] T258;
  wire[20:0] T259;
  wire[19:0] T260;
  wire[19:0] T261;
  wire[18:0] T262;
  wire[18:0] T263;
  wire[17:0] T264;
  wire[17:0] T265;
  wire[16:0] T266;
  wire[16:0] T267;
  wire[15:0] T268;
  wire[15:0] T269;
  wire[14:0] T270;
  wire[14:0] T271;
  wire[13:0] T272;
  wire[13:0] T273;
  wire[12:0] T274;
  wire[12:0] T275;
  wire[11:0] T276;
  wire[11:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire[9:0] T280;
  wire[9:0] T281;
  wire[8:0] T282;
  wire[8:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[6:0] T286;
  wire[6:0] T287;
  wire[5:0] T288;
  wire[5:0] T289;
  wire[4:0] T290;
  wire[4:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire[1:0] T296;
  wire[1:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] T303;
  wire[2:0] T304;
  wire[2:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire[1:0] T309;
  wire[1:0] T310;
  wire[1:0] T311;
  wire[2:0] T312;
  wire[2:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[2:0] T320;
  wire[2:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire[3:0] T325;
  wire[3:0] T326;
  wire[3:0] T327;
  wire[10:0] T328;
  wire[10:0] T329;
  wire T330;
  wire T331;
  wire T332;
  wire[1:0] T333;
  wire[1:0] T334;
  wire[1:0] T335;
  wire[2:0] T336;
  wire[2:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire[1:0] T341;
  wire[1:0] T342;
  wire[1:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire[1:0] T349;
  wire[1:0] T350;
  wire[1:0] T351;
  wire[2:0] T352;
  wire[2:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire[1:0] T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire[2:0] T360;
  wire[2:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire[3:0] T365;
  wire[3:0] T366;
  wire[3:0] T367;
  wire[10:0] T368;
  wire[10:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire[1:0] T373;
  wire[1:0] T374;
  wire[1:0] T375;
  wire[2:0] T376;
  wire[2:0] T377;
  wire T378;
  wire T379;
  wire T380;
  wire[1:0] T381;
  wire[1:0] T382;
  wire[1:0] T383;
  wire[2:0] T384;
  wire[2:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire[1:0] T389;
  wire[1:0] T390;
  wire[1:0] T391;
  wire[2:0] T392;
  wire[2:0] T393;
  wire T394;
  wire T395;
  wire T396;
  wire[1:0] T397;
  wire[1:0] T398;
  wire[1:0] T399;
  wire[2:0] T400;
  wire[2:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire[3:0] T405;
  wire[3:0] T406;
  wire[3:0] T407;
  wire[10:0] T408;
  wire[10:0] T409;
  wire T410;
  wire T411;
  wire T412;
  wire[1:0] T413;
  wire[1:0] T414;
  wire[1:0] T415;
  wire[2:0] T416;
  wire[2:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire[1:0] T421;
  wire[1:0] T422;
  wire[1:0] T423;
  wire[2:0] T424;
  wire[2:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire[1:0] T431;
  wire[2:0] T432;
  wire[2:0] T433;
  wire T434;
  wire T435;
  wire T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[2:0] T440;
  wire[2:0] T441;
  wire T442;
  wire T443;
  wire T444;
  wire[3:0] T445;
  wire[3:0] T446;
  wire[3:0] T447;
  wire[10:0] T448;
  wire[10:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire[1:0] T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire T458;
  wire T459;
  wire T460;
  wire[1:0] T461;
  wire[1:0] T462;
  wire[1:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire[1:0] T469;
  wire[1:0] T470;
  wire[1:0] T471;
  wire[2:0] T472;
  wire[2:0] T473;
  wire T474;
  wire T475;
  wire T476;
  wire[1:0] T477;
  wire[1:0] T478;
  wire[1:0] T479;
  wire[2:0] T480;
  wire[2:0] T481;
  wire T482;
  wire T483;
  wire T484;
  wire[3:0] T485;
  wire[3:0] T486;
  wire[3:0] T487;
  wire[10:0] T488;
  wire[10:0] T489;
  wire T490;
  wire T491;
  wire T492;
  wire[1:0] T493;
  wire[1:0] T494;
  wire[1:0] T495;
  wire[2:0] T496;
  wire[2:0] T497;
  wire T498;
  wire T499;
  wire T500;
  wire[1:0] T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire[2:0] T504;
  wire[2:0] T505;
  wire T506;
  wire T507;
  wire T508;
  wire[1:0] T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire[2:0] T512;
  wire[2:0] T513;
  wire T514;
  wire T515;
  wire T516;
  wire[1:0] T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire[2:0] T520;
  wire[2:0] T521;
  wire T522;
  wire T523;
  wire T524;
  wire[3:0] T525;
  wire[3:0] T526;
  wire[3:0] T527;
  wire[10:0] T528;
  wire[10:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire[1:0] T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire[2:0] T536;
  wire[2:0] T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire[1:0] T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[1:0] T552;
  wire[1:0] T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire[1:0] T560;
  wire[1:0] T561;
  wire T562;
  wire T563;
  wire T564;
  wire[3:0] T565;
  wire[3:0] T566;
  wire[3:0] T567;
  wire[10:0] T568;
  wire[10:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire[1:0] T576;
  wire[1:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire[1:0] T584;
  wire[1:0] T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[1:0] T592;
  wire[1:0] T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire[1:0] T600;
  wire[1:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire[3:0] T605;
  wire[3:0] T606;
  wire[3:0] T607;
  wire[10:0] T608;
  wire[10:0] T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire[1:0] T616;
  wire[1:0] T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[1:0] T624;
  wire[1:0] T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[1:0] T632;
  wire[1:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire[1:0] T640;
  wire[1:0] T641;
  wire T642;
  wire T643;
  wire T644;
  wire[3:0] T645;
  wire[3:0] T646;
  wire[3:0] T647;
  wire[10:0] T648;
  wire[10:0] T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire[1:0] T656;
  wire[1:0] T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire[1:0] T664;
  wire[1:0] T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire[1:0] T672;
  wire[1:0] T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire[1:0] T680;
  wire[1:0] T681;
  wire T682;
  wire T683;
  wire T684;
  wire[3:0] T685;
  wire[3:0] T686;
  wire[3:0] T687;
  wire[9:0] T688;
  wire[9:0] T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire T694;
  wire T695;
  wire[1:0] T696;
  wire[1:0] T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire[1:0] T704;
  wire[1:0] T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire[1:0] T712;
  wire[1:0] T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[1:0] T720;
  wire[1:0] T721;
  wire T722;
  wire T723;
  wire T724;
  wire[3:0] T725;
  wire[3:0] T726;
  wire[3:0] T727;
  wire[9:0] T728;
  wire[9:0] T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire[1:0] T736;
  wire[1:0] T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire[1:0] T744;
  wire[1:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire[1:0] T752;
  wire[1:0] T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire[1:0] T760;
  wire[1:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire[3:0] T765;
  wire[3:0] T766;
  wire[3:0] T767;
  wire[9:0] T768;
  wire[9:0] T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire[1:0] T776;
  wire[1:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[1:0] T784;
  wire[1:0] T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire[1:0] T792;
  wire[1:0] T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire[1:0] T800;
  wire[1:0] T801;
  wire T802;
  wire T803;
  wire T804;
  wire[3:0] T805;
  wire[3:0] T806;
  wire[3:0] T807;
  wire[9:0] T808;
  wire[9:0] T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire[1:0] T816;
  wire[1:0] T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire[1:0] T824;
  wire[1:0] T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire[1:0] T832;
  wire[1:0] T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire[1:0] T840;
  wire[1:0] T841;
  wire T842;
  wire T843;
  wire T844;
  wire[3:0] T845;
  wire[3:0] T846;
  wire[3:0] T847;
  wire[9:0] T848;
  wire[9:0] T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire[1:0] T856;
  wire[1:0] T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire[1:0] T864;
  wire[1:0] T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire[1:0] T872;
  wire[1:0] T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire[1:0] T880;
  wire[1:0] T881;
  wire T882;
  wire T883;
  wire T884;
  wire[3:0] T885;
  wire[3:0] T886;
  wire[3:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire[1:0] T896;
  wire[1:0] T897;
  wire T898;
  wire T899;
  wire T900;
  wire[1:0] T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire[2:0] T904;
  wire[2:0] T905;
  wire T906;
  wire T907;
  wire T908;
  wire[1:0] T909;
  wire[1:0] T910;
  wire[1:0] T911;
  wire[2:0] T912;
  wire[2:0] T913;
  wire T914;
  wire T915;
  wire T916;
  wire[1:0] T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire[2:0] T920;
  wire[2:0] T921;
  wire T922;
  wire T923;
  wire T924;
  wire[3:0] T925;
  wire[3:0] T926;
  wire[3:0] T927;
  wire[10:0] T928;
  wire[10:0] T929;
  wire T930;
  wire T931;
  wire T932;
  wire[1:0] T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire[2:0] T936;
  wire[2:0] T937;
  wire T938;
  wire T939;
  wire T940;
  wire[1:0] T941;
  wire[1:0] T942;
  wire[1:0] T943;
  wire[2:0] T944;
  wire[2:0] T945;
  wire T946;
  wire T947;
  wire T948;
  wire[1:0] T949;
  wire[1:0] T950;
  wire[1:0] T951;
  wire[2:0] T952;
  wire[2:0] T953;
  wire T954;
  wire T955;
  wire T956;
  wire[1:0] T957;
  wire[1:0] T958;
  wire[1:0] T959;
  wire[2:0] T960;
  wire[2:0] T961;
  wire T962;
  wire T963;
  wire T964;
  wire[3:0] T965;
  wire[3:0] T966;
  wire[3:0] T967;
  wire[10:0] T968;
  wire[10:0] T969;
  wire T970;
  wire T971;
  wire T972;
  wire[1:0] T973;
  wire[1:0] T974;
  wire[1:0] T975;
  wire[2:0] T976;
  wire[2:0] T977;
  wire T978;
  wire T979;
  wire T980;
  wire[1:0] T981;
  wire[1:0] T982;
  wire[1:0] T983;
  wire[2:0] T984;
  wire[2:0] T985;
  wire T986;
  wire T987;
  wire T988;
  wire[1:0] T989;
  wire[1:0] T990;
  wire[1:0] T991;
  wire[2:0] T992;
  wire[2:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire[1:0] T997;
  wire[1:0] T998;
  wire[1:0] T999;
  wire[2:0] T1000;
  wire[2:0] T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire[3:0] T1005;
  wire[3:0] T1006;
  wire[3:0] T1007;
  wire[10:0] T1008;
  wire[10:0] T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire[1:0] T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire[2:0] T1016;
  wire[2:0] T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire[1:0] T1021;
  wire[1:0] T1022;
  wire[1:0] T1023;
  wire[2:0] T1024;
  wire[2:0] T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire[1:0] T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire[2:0] T1032;
  wire[2:0] T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire[1:0] T1037;
  wire[1:0] T1038;
  wire[1:0] T1039;
  wire[2:0] T1040;
  wire[2:0] T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire[3:0] T1045;
  wire[3:0] T1046;
  wire[3:0] T1047;
  wire[10:0] T1048;
  wire[10:0] T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire[1:0] T1053;
  wire[1:0] T1054;
  wire[1:0] T1055;
  wire[2:0] T1056;
  wire[2:0] T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire[1:0] T1061;
  wire[1:0] T1062;
  wire[1:0] T1063;
  wire[2:0] T1064;
  wire[2:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire[1:0] T1069;
  wire[1:0] T1070;
  wire[1:0] T1071;
  wire[2:0] T1072;
  wire[2:0] T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire[1:0] T1077;
  wire[1:0] T1078;
  wire[1:0] T1079;
  wire[2:0] T1080;
  wire[2:0] T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire[3:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[10:0] T1088;
  wire[10:0] T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire[1:0] T1093;
  wire[1:0] T1094;
  wire[1:0] T1095;
  wire[2:0] T1096;
  wire[2:0] T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire[1:0] T1101;
  wire[1:0] T1102;
  wire[1:0] T1103;
  wire[2:0] T1104;
  wire[2:0] T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire[1:0] T1109;
  wire[1:0] T1110;
  wire[1:0] T1111;
  wire[2:0] T1112;
  wire[2:0] T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire[1:0] T1117;
  wire[1:0] T1118;
  wire[1:0] T1119;
  wire[2:0] T1120;
  wire[2:0] T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire[3:0] T1125;
  wire[3:0] T1126;
  wire[3:0] T1127;
  wire[10:0] T1128;
  wire[10:0] T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire[1:0] T1133;
  wire[1:0] T1134;
  wire[1:0] T1135;
  wire[2:0] T1136;
  wire[2:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[1:0] T1144;
  wire[1:0] T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire[1:0] T1152;
  wire[1:0] T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire[1:0] T1160;
  wire[1:0] T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire[3:0] T1165;
  wire[3:0] T1166;
  wire[3:0] T1167;
  wire[10:0] T1168;
  wire[10:0] T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire[1:0] T1176;
  wire[1:0] T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire[1:0] T1184;
  wire[1:0] T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire[1:0] T1192;
  wire[1:0] T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire[1:0] T1200;
  wire[1:0] T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire[3:0] T1205;
  wire[3:0] T1206;
  wire[3:0] T1207;
  wire[10:0] T1208;
  wire[10:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire[1:0] T1216;
  wire[1:0] T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire[1:0] T1224;
  wire[1:0] T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire[1:0] T1232;
  wire[1:0] T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire[1:0] T1240;
  wire[1:0] T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire[3:0] T1245;
  wire[3:0] T1246;
  wire[3:0] T1247;
  wire[10:0] T1248;
  wire[10:0] T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire[1:0] T1256;
  wire[1:0] T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire[1:0] T1264;
  wire[1:0] T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire[1:0] T1272;
  wire[1:0] T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire[1:0] T1280;
  wire[1:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire[3:0] T1285;
  wire[3:0] T1286;
  wire[3:0] T1287;
  wire[9:0] T1288;
  wire[9:0] T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire T1293;
  wire T1294;
  wire T1295;
  wire[1:0] T1296;
  wire[1:0] T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire[1:0] T1304;
  wire[1:0] T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire[1:0] T1312;
  wire[1:0] T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire[1:0] T1320;
  wire[1:0] T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire[3:0] T1325;
  wire[3:0] T1326;
  wire[3:0] T1327;
  wire[9:0] T1328;
  wire[9:0] T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire[1:0] T1336;
  wire[1:0] T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire T1343;
  wire[1:0] T1344;
  wire[1:0] T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[1:0] T1352;
  wire[1:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire[1:0] T1360;
  wire[1:0] T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire[3:0] T1365;
  wire[3:0] T1366;
  wire[3:0] T1367;
  wire[9:0] T1368;
  wire[9:0] T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire[1:0] T1376;
  wire[1:0] T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire[1:0] T1384;
  wire[1:0] T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire[1:0] T1392;
  wire[1:0] T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[1:0] T1400;
  wire[1:0] T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire[3:0] T1405;
  wire[3:0] T1406;
  wire[3:0] T1407;
  wire[9:0] T1408;
  wire[9:0] T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire T1414;
  wire T1415;
  wire[1:0] T1416;
  wire[1:0] T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire T1421;
  wire T1422;
  wire T1423;
  wire[1:0] T1424;
  wire[1:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[1:0] T1432;
  wire[1:0] T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire T1437;
  wire T1438;
  wire T1439;
  wire[1:0] T1440;
  wire[1:0] T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire[3:0] T1445;
  wire[3:0] T1446;
  wire[3:0] T1447;
  wire[9:0] T1448;
  wire[9:0] T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire[1:0] T1456;
  wire[1:0] T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire[1:0] T1464;
  wire[1:0] T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire[1:0] T1472;
  wire[1:0] T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire T1478;
  wire T1479;
  wire[1:0] T1480;
  wire[1:0] T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire[3:0] T1485;
  wire[3:0] T1486;
  wire[3:0] T1487;
  wire[9:0] T1488;
  wire[9:0] T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[1:0] T1496;
  wire[1:0] T1497;
  wire[22:0] T1498;
  wire[22:0] T1499;
  wire[21:0] T1500;
  wire[21:0] T1501;
  wire[20:0] T1502;
  wire[20:0] T1503;
  wire[19:0] T1504;
  wire[19:0] T1505;
  wire[18:0] T1506;
  wire[18:0] T1507;
  wire[17:0] T1508;
  wire[17:0] T1509;
  wire[16:0] T1510;
  wire[16:0] T1511;
  wire[15:0] T1512;
  wire[15:0] T1513;
  wire[14:0] T1514;
  wire[14:0] T1515;
  wire[13:0] T1516;
  wire[13:0] T1517;
  wire[12:0] T1518;
  wire[12:0] T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[10:0] T1522;
  wire[10:0] T1523;
  wire[9:0] T1524;
  wire[9:0] T1525;
  wire[8:0] T1526;
  wire[8:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[6:0] T1530;
  wire[6:0] T1531;
  wire[5:0] T1532;
  wire[5:0] T1533;
  wire[4:0] T1534;
  wire[4:0] T1535;
  wire[3:0] T1536;
  wire[3:0] T1537;
  wire[2:0] T1538;
  wire[2:0] T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[11:0] T1660;
  wire[11:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[11:0] T1668;
  wire[11:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[11:0] T1676;
  wire[11:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[11:0] T1684;
  wire[11:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[11:0] T1692;
  wire[11:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[11:0] T1700;
  wire[11:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[11:0] T1708;
  wire[11:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[11:0] T1716;
  wire[11:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[11:0] T1724;
  wire[11:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1490, T2};
  assign T2 = T3;
  assign T3 = {T1482, T4};
  assign T4 = T5;
  assign T5 = {T1474, T6};
  assign T6 = T7;
  assign T7 = {T1466, T8};
  assign T8 = T9;
  assign T9 = {T1458, T10};
  assign T10 = T11;
  assign T11 = {T1450, T12};
  assign T12 = T13;
  assign T13 = {T1442, T14};
  assign T14 = T15;
  assign T15 = {T1434, T16};
  assign T16 = T17;
  assign T17 = {T1426, T18};
  assign T18 = T19;
  assign T19 = {T1418, T20};
  assign T20 = T21;
  assign T21 = {T1410, T22};
  assign T22 = T23;
  assign T23 = {T1402, T24};
  assign T24 = T25;
  assign T25 = {T1394, T26};
  assign T26 = T27;
  assign T27 = {T1386, T28};
  assign T28 = T29;
  assign T29 = {T1378, T30};
  assign T30 = T31;
  assign T31 = {T1370, T32};
  assign T32 = T33;
  assign T33 = {T1362, T34};
  assign T34 = T35;
  assign T35 = {T1354, T36};
  assign T36 = T37;
  assign T37 = {T1346, T38};
  assign T38 = T39;
  assign T39 = {T1338, T40};
  assign T40 = T41;
  assign T41 = {T1330, T42};
  assign T42 = T43;
  assign T43 = {T1322, T44};
  assign T44 = T45;
  assign T45 = {T1314, T46};
  assign T46 = T47;
  assign T47 = {T1306, T48};
  assign T48 = T49;
  assign T49 = {T1298, T50};
  assign T50 = T51;
  assign T51 = {T1290, T52};
  assign T52 = T53;
  assign T53 = {T1282, T54};
  assign T54 = T55;
  assign T55 = {T1274, T56};
  assign T56 = T57;
  assign T57 = {T1266, T58};
  assign T58 = T59;
  assign T59 = {T1258, T60};
  assign T60 = T61;
  assign T61 = {T1250, T62};
  assign T62 = T63;
  assign T63 = {T1242, T64};
  assign T64 = T65;
  assign T65 = {T1234, T66};
  assign T66 = T67;
  assign T67 = {T1226, T68};
  assign T68 = T69;
  assign T69 = {T1218, T70};
  assign T70 = T71;
  assign T71 = {T1210, T72};
  assign T72 = T73;
  assign T73 = {T1202, T74};
  assign T74 = T75;
  assign T75 = {T1194, T76};
  assign T76 = T77;
  assign T77 = {T1186, T78};
  assign T78 = T79;
  assign T79 = {T1178, T80};
  assign T80 = T81;
  assign T81 = {T1170, T82};
  assign T82 = T83;
  assign T83 = {T1162, T84};
  assign T84 = T85;
  assign T85 = {T1154, T86};
  assign T86 = T87;
  assign T87 = {T1146, T88};
  assign T88 = T89;
  assign T89 = {T1138, T90};
  assign T90 = T91;
  assign T91 = {T1130, T92};
  assign T92 = T93;
  assign T93 = {T1122, T94};
  assign T94 = T95;
  assign T95 = {T1114, T96};
  assign T96 = T97;
  assign T97 = {T1106, T98};
  assign T98 = T99;
  assign T99 = {T1098, T100};
  assign T100 = T101;
  assign T101 = {T1090, T102};
  assign T102 = T103;
  assign T103 = {T1082, T104};
  assign T104 = T105;
  assign T105 = {T1074, T106};
  assign T106 = T107;
  assign T107 = {T1066, T108};
  assign T108 = T109;
  assign T109 = {T1058, T110};
  assign T110 = T111;
  assign T111 = {T1050, T112};
  assign T112 = T113;
  assign T113 = {T1042, T114};
  assign T114 = T115;
  assign T115 = {T1034, T116};
  assign T116 = T117;
  assign T117 = {T1026, T118};
  assign T118 = T119;
  assign T119 = {T1018, T120};
  assign T120 = T121;
  assign T121 = {T1010, T122};
  assign T122 = T123;
  assign T123 = {T1002, T124};
  assign T124 = T125;
  assign T125 = {T994, T126};
  assign T126 = T127;
  assign T127 = {T986, T128};
  assign T128 = T129;
  assign T129 = {T978, T130};
  assign T130 = T131;
  assign T131 = {T970, T132};
  assign T132 = T133;
  assign T133 = {T962, T134};
  assign T134 = T135;
  assign T135 = {T954, T136};
  assign T136 = T137;
  assign T137 = {T946, T138};
  assign T138 = T139;
  assign T139 = {T938, T140};
  assign T140 = T141;
  assign T141 = {T930, T142};
  assign T142 = T143;
  assign T143 = {T922, T144};
  assign T144 = T145;
  assign T145 = {T914, T146};
  assign T146 = T147;
  assign T147 = {T906, T148};
  assign T148 = T149;
  assign T149 = {T898, T150};
  assign T150 = T151;
  assign T151 = {T890, T152};
  assign T152 = T153;
  assign T153 = {T882, T154};
  assign T154 = T155;
  assign T155 = {T874, T156};
  assign T156 = T157;
  assign T157 = {T866, T158};
  assign T158 = T159;
  assign T159 = {T858, T160};
  assign T160 = T161;
  assign T161 = {T850, T162};
  assign T162 = T163;
  assign T163 = {T842, T164};
  assign T164 = T165;
  assign T165 = {T834, T166};
  assign T166 = T167;
  assign T167 = {T826, T168};
  assign T168 = T169;
  assign T169 = {T818, T170};
  assign T170 = T171;
  assign T171 = {T810, T172};
  assign T172 = T173;
  assign T173 = {T802, T174};
  assign T174 = T175;
  assign T175 = {T794, T176};
  assign T176 = T177;
  assign T177 = {T786, T178};
  assign T178 = T179;
  assign T179 = {T778, T180};
  assign T180 = T181;
  assign T181 = {T770, T182};
  assign T182 = T183;
  assign T183 = {T762, T184};
  assign T184 = T185;
  assign T185 = {T754, T186};
  assign T186 = T187;
  assign T187 = {T746, T188};
  assign T188 = T189;
  assign T189 = {T738, T190};
  assign T190 = T191;
  assign T191 = {T730, T192};
  assign T192 = T193;
  assign T193 = {T722, T194};
  assign T194 = T195;
  assign T195 = {T714, T196};
  assign T196 = T197;
  assign T197 = {T706, T198};
  assign T198 = T199;
  assign T199 = {T698, T200};
  assign T200 = T201;
  assign T201 = {T690, T202};
  assign T202 = T203;
  assign T203 = {T682, T204};
  assign T204 = T205;
  assign T205 = {T674, T206};
  assign T206 = T207;
  assign T207 = {T666, T208};
  assign T208 = T209;
  assign T209 = {T658, T210};
  assign T210 = T211;
  assign T211 = {T650, T212};
  assign T212 = T213;
  assign T213 = {T642, T214};
  assign T214 = T215;
  assign T215 = {T634, T216};
  assign T216 = T217;
  assign T217 = {T626, T218};
  assign T218 = T219;
  assign T219 = {T618, T220};
  assign T220 = T221;
  assign T221 = {T610, T222};
  assign T222 = T223;
  assign T223 = {T602, T224};
  assign T224 = T225;
  assign T225 = {T594, T226};
  assign T226 = T227;
  assign T227 = {T586, T228};
  assign T228 = T229;
  assign T229 = {T578, T230};
  assign T230 = T231;
  assign T231 = {T570, T232};
  assign T232 = T233;
  assign T233 = {T562, T234};
  assign T234 = T235;
  assign T235 = {T554, T236};
  assign T236 = T237;
  assign T237 = {T546, T238};
  assign T238 = T239;
  assign T239 = {T538, T240};
  assign T240 = T241;
  assign T241 = {T530, T242};
  assign T242 = T243;
  assign T243 = {T522, T244};
  assign T244 = T245;
  assign T245 = {T514, T246};
  assign T246 = T247;
  assign T247 = {T506, T248};
  assign T248 = T249;
  assign T249 = {T498, T250};
  assign T250 = T251;
  assign T251 = {T490, T252};
  assign T252 = T253;
  assign T253 = {T482, T254};
  assign T254 = T255;
  assign T255 = {T474, T256};
  assign T256 = T257;
  assign T257 = {T466, T258};
  assign T258 = T259;
  assign T259 = {T458, T260};
  assign T260 = T261;
  assign T261 = {T450, T262};
  assign T262 = T263;
  assign T263 = {T442, T264};
  assign T264 = T265;
  assign T265 = {T434, T266};
  assign T266 = T267;
  assign T267 = {T426, T268};
  assign T268 = T269;
  assign T269 = {T418, T270};
  assign T270 = T271;
  assign T271 = {T410, T272};
  assign T272 = T273;
  assign T273 = {T402, T274};
  assign T274 = T275;
  assign T275 = {T394, T276};
  assign T276 = T277;
  assign T277 = {T386, T278};
  assign T278 = T279;
  assign T279 = {T378, T280};
  assign T280 = T281;
  assign T281 = {T370, T282};
  assign T282 = T283;
  assign T283 = {T362, T284};
  assign T284 = T285;
  assign T285 = {T354, T286};
  assign T286 = T287;
  assign T287 = {T346, T288};
  assign T288 = T289;
  assign T289 = {T338, T290};
  assign T290 = T291;
  assign T291 = {T330, T292};
  assign T292 = T293;
  assign T293 = {T322, T294};
  assign T294 = T295;
  assign T295 = {T314, T296};
  assign T296 = T297;
  assign T297 = {T306, T298};
  assign T298 = T299;
  assign T299 = T300;
  assign T300 = T304[T301];
  assign T301 = T302;
  assign T302 = T303;
  assign T303 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T304 = T305;
  assign T305 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T306 = T307;
  assign T307 = T308;
  assign T308 = T312[T309];
  assign T309 = T310;
  assign T310 = T311;
  assign T311 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T312 = T313;
  assign T313 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T314 = T315;
  assign T315 = T316;
  assign T316 = T320[T317];
  assign T317 = T318;
  assign T318 = T319;
  assign T319 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T320 = T321;
  assign T321 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T322 = T323;
  assign T323 = T324;
  assign T324 = T328[T325];
  assign T325 = T326;
  assign T326 = T327;
  assign T327 = io_chanxy_config[4'h9/* 9*/:3'h6/* 6*/];
  assign T328 = T329;
  assign T329 = io_chanxy_in[5'h13/* 19*/:4'h9/* 9*/];
  assign T330 = T331;
  assign T331 = T332;
  assign T332 = T336[T333];
  assign T333 = T334;
  assign T334 = T335;
  assign T335 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T336 = T337;
  assign T337 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T338 = T339;
  assign T339 = T340;
  assign T340 = T344[T341];
  assign T341 = T342;
  assign T342 = T343;
  assign T343 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T344 = T345;
  assign T345 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T346 = T347;
  assign T347 = T348;
  assign T348 = T352[T349];
  assign T349 = T350;
  assign T350 = T351;
  assign T351 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T352 = T353;
  assign T353 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T354 = T355;
  assign T355 = T356;
  assign T356 = T360[T357];
  assign T357 = T358;
  assign T358 = T359;
  assign T359 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T360 = T361;
  assign T361 = io_chanxy_in[5'h1f/* 31*/:5'h1d/* 29*/];
  assign T362 = T363;
  assign T363 = T364;
  assign T364 = T368[T365];
  assign T365 = T366;
  assign T366 = T367;
  assign T367 = io_chanxy_config[5'h15/* 21*/:5'h12/* 18*/];
  assign T368 = T369;
  assign T369 = io_chanxy_in[6'h2a/* 42*/:6'h20/* 32*/];
  assign T370 = T371;
  assign T371 = T372;
  assign T372 = T376[T373];
  assign T373 = T374;
  assign T374 = T375;
  assign T375 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T376 = T377;
  assign T377 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T378 = T379;
  assign T379 = T380;
  assign T380 = T384[T381];
  assign T381 = T382;
  assign T382 = T383;
  assign T383 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T384 = T385;
  assign T385 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T386 = T387;
  assign T387 = T388;
  assign T388 = T392[T389];
  assign T389 = T390;
  assign T390 = T391;
  assign T391 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T392 = T393;
  assign T393 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T394 = T395;
  assign T395 = T396;
  assign T396 = T400[T397];
  assign T397 = T398;
  assign T398 = T399;
  assign T399 = io_chanxy_config[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T400 = T401;
  assign T401 = io_chanxy_in[6'h36/* 54*/:6'h34/* 52*/];
  assign T402 = T403;
  assign T403 = T404;
  assign T404 = T408[T405];
  assign T405 = T406;
  assign T406 = T407;
  assign T407 = io_chanxy_config[6'h21/* 33*/:5'h1e/* 30*/];
  assign T408 = T409;
  assign T409 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T410 = T411;
  assign T411 = T412;
  assign T412 = T416[T413];
  assign T413 = T414;
  assign T414 = T415;
  assign T415 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T416 = T417;
  assign T417 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T418 = T419;
  assign T419 = T420;
  assign T420 = T424[T421];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T424 = T425;
  assign T425 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T426 = T427;
  assign T427 = T428;
  assign T428 = T432[T429];
  assign T429 = T430;
  assign T430 = T431;
  assign T431 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T432 = T433;
  assign T433 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T434 = T435;
  assign T435 = T436;
  assign T436 = T440[T437];
  assign T437 = T438;
  assign T438 = T439;
  assign T439 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T440 = T441;
  assign T441 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = T448[T445];
  assign T445 = T446;
  assign T446 = T447;
  assign T447 = io_chanxy_config[6'h2d/* 45*/:6'h2a/* 42*/];
  assign T448 = T449;
  assign T449 = io_chanxy_in[7'h58/* 88*/:7'h4e/* 78*/];
  assign T450 = T451;
  assign T451 = T452;
  assign T452 = T456[T453];
  assign T453 = T454;
  assign T454 = T455;
  assign T455 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T456 = T457;
  assign T457 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T458 = T459;
  assign T459 = T460;
  assign T460 = T464[T461];
  assign T461 = T462;
  assign T462 = T463;
  assign T463 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T464 = T465;
  assign T465 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T472[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T472 = T473;
  assign T473 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T474 = T475;
  assign T475 = T476;
  assign T476 = T480[T477];
  assign T477 = T478;
  assign T478 = T479;
  assign T479 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T480 = T481;
  assign T481 = io_chanxy_in[7'h64/* 100*/:7'h62/* 98*/];
  assign T482 = T483;
  assign T483 = T484;
  assign T484 = T488[T485];
  assign T485 = T486;
  assign T486 = T487;
  assign T487 = io_chanxy_config[6'h39/* 57*/:6'h36/* 54*/];
  assign T488 = T489;
  assign T489 = io_chanxy_in[7'h6f/* 111*/:7'h65/* 101*/];
  assign T490 = T491;
  assign T491 = T492;
  assign T492 = T496[T493];
  assign T493 = T494;
  assign T494 = T495;
  assign T495 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T496 = T497;
  assign T497 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T498 = T499;
  assign T499 = T500;
  assign T500 = T504[T501];
  assign T501 = T502;
  assign T502 = T503;
  assign T503 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T504 = T505;
  assign T505 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T506 = T507;
  assign T507 = T508;
  assign T508 = T512[T509];
  assign T509 = T510;
  assign T510 = T511;
  assign T511 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T512 = T513;
  assign T513 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T514 = T515;
  assign T515 = T516;
  assign T516 = T520[T517];
  assign T517 = T518;
  assign T518 = T519;
  assign T519 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T520 = T521;
  assign T521 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T522 = T523;
  assign T523 = T524;
  assign T524 = T528[T525];
  assign T525 = T526;
  assign T526 = T527;
  assign T527 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T528 = T529;
  assign T529 = io_chanxy_in[8'h86/* 134*/:7'h7c/* 124*/];
  assign T530 = T531;
  assign T531 = T532;
  assign T532 = T536[T533];
  assign T533 = T534;
  assign T534 = T535;
  assign T535 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T536 = T537;
  assign T537 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T538 = T539;
  assign T539 = T540;
  assign T540 = T544[T541];
  assign T541 = T542;
  assign T542 = T543;
  assign T543 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T544 = T545;
  assign T545 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T546 = T547;
  assign T547 = T548;
  assign T548 = T552[T549];
  assign T549 = T550;
  assign T550 = T551;
  assign T551 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T552 = T553;
  assign T553 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T554 = T555;
  assign T555 = T556;
  assign T556 = T560[T557];
  assign T557 = T558;
  assign T558 = T559;
  assign T559 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T560 = T561;
  assign T561 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T562 = T563;
  assign T563 = T564;
  assign T564 = T568[T565];
  assign T565 = T566;
  assign T566 = T567;
  assign T567 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T568 = T569;
  assign T569 = io_chanxy_in[8'h9a/* 154*/:8'h90/* 144*/];
  assign T570 = T571;
  assign T571 = T572;
  assign T572 = T576[T573];
  assign T573 = T574;
  assign T574 = T575;
  assign T575 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T576 = T577;
  assign T577 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T578 = T579;
  assign T579 = T580;
  assign T580 = T584[T581];
  assign T581 = T582;
  assign T582 = T583;
  assign T583 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T584 = T585;
  assign T585 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T586 = T587;
  assign T587 = T588;
  assign T588 = T592[T589];
  assign T589 = T590;
  assign T590 = T591;
  assign T591 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T592 = T593;
  assign T593 = io_chanxy_in[8'ha0/* 160*/:8'h9f/* 159*/];
  assign T594 = T595;
  assign T595 = T596;
  assign T596 = T600[T597];
  assign T597 = T598;
  assign T598 = T599;
  assign T599 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T600 = T601;
  assign T601 = io_chanxy_in[8'ha2/* 162*/:8'ha1/* 161*/];
  assign T602 = T603;
  assign T603 = T604;
  assign T604 = T608[T605];
  assign T605 = T606;
  assign T606 = T607;
  assign T607 = io_chanxy_config[7'h56/* 86*/:7'h53/* 83*/];
  assign T608 = T609;
  assign T609 = io_chanxy_in[8'had/* 173*/:8'ha3/* 163*/];
  assign T610 = T611;
  assign T611 = T612;
  assign T612 = T616[T613];
  assign T613 = T614;
  assign T614 = T615;
  assign T615 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T616 = T617;
  assign T617 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T618 = T619;
  assign T619 = T620;
  assign T620 = T624[T621];
  assign T621 = T622;
  assign T622 = T623;
  assign T623 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T624 = T625;
  assign T625 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T626 = T627;
  assign T627 = T628;
  assign T628 = T632[T629];
  assign T629 = T630;
  assign T630 = T631;
  assign T631 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T632 = T633;
  assign T633 = io_chanxy_in[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T634 = T635;
  assign T635 = T636;
  assign T636 = T640[T637];
  assign T637 = T638;
  assign T638 = T639;
  assign T639 = io_chanxy_config[7'h5a/* 90*/:7'h5a/* 90*/];
  assign T640 = T641;
  assign T641 = io_chanxy_in[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T642 = T643;
  assign T643 = T644;
  assign T644 = T648[T645];
  assign T645 = T646;
  assign T646 = T647;
  assign T647 = io_chanxy_config[7'h5e/* 94*/:7'h5b/* 91*/];
  assign T648 = T649;
  assign T649 = io_chanxy_in[8'hc0/* 192*/:8'hb6/* 182*/];
  assign T650 = T651;
  assign T651 = T652;
  assign T652 = T656[T653];
  assign T653 = T654;
  assign T654 = T655;
  assign T655 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T656 = T657;
  assign T657 = io_chanxy_in[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T658 = T659;
  assign T659 = T660;
  assign T660 = T664[T661];
  assign T661 = T662;
  assign T662 = T663;
  assign T663 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T664 = T665;
  assign T665 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T666 = T667;
  assign T667 = T668;
  assign T668 = T672[T669];
  assign T669 = T670;
  assign T670 = T671;
  assign T671 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T672 = T673;
  assign T673 = io_chanxy_in[8'hc6/* 198*/:8'hc5/* 197*/];
  assign T674 = T675;
  assign T675 = T676;
  assign T676 = T680[T677];
  assign T677 = T678;
  assign T678 = T679;
  assign T679 = io_chanxy_config[7'h62/* 98*/:7'h62/* 98*/];
  assign T680 = T681;
  assign T681 = io_chanxy_in[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T682 = T683;
  assign T683 = T684;
  assign T684 = T688[T685];
  assign T685 = T686;
  assign T686 = T687;
  assign T687 = io_chanxy_config[7'h66/* 102*/:7'h63/* 99*/];
  assign T688 = T689;
  assign T689 = io_chanxy_in[8'hd2/* 210*/:8'hc9/* 201*/];
  assign T690 = T691;
  assign T691 = T692;
  assign T692 = T696[T693];
  assign T693 = T694;
  assign T694 = T695;
  assign T695 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T696 = T697;
  assign T697 = io_chanxy_in[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T698 = T699;
  assign T699 = T700;
  assign T700 = T704[T701];
  assign T701 = T702;
  assign T702 = T703;
  assign T703 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T704 = T705;
  assign T705 = io_chanxy_in[8'hd6/* 214*/:8'hd5/* 213*/];
  assign T706 = T707;
  assign T707 = T708;
  assign T708 = T712[T709];
  assign T709 = T710;
  assign T710 = T711;
  assign T711 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T712 = T713;
  assign T713 = io_chanxy_in[8'hd8/* 216*/:8'hd7/* 215*/];
  assign T714 = T715;
  assign T715 = T716;
  assign T716 = T720[T717];
  assign T717 = T718;
  assign T718 = T719;
  assign T719 = io_chanxy_config[7'h6a/* 106*/:7'h6a/* 106*/];
  assign T720 = T721;
  assign T721 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T722 = T723;
  assign T723 = T724;
  assign T724 = T728[T725];
  assign T725 = T726;
  assign T726 = T727;
  assign T727 = io_chanxy_config[7'h6e/* 110*/:7'h6b/* 107*/];
  assign T728 = T729;
  assign T729 = io_chanxy_in[8'he4/* 228*/:8'hdb/* 219*/];
  assign T730 = T731;
  assign T731 = T732;
  assign T732 = T736[T733];
  assign T733 = T734;
  assign T734 = T735;
  assign T735 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T736 = T737;
  assign T737 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T738 = T739;
  assign T739 = T740;
  assign T740 = T744[T741];
  assign T741 = T742;
  assign T742 = T743;
  assign T743 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T744 = T745;
  assign T745 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T746 = T747;
  assign T747 = T748;
  assign T748 = T752[T749];
  assign T749 = T750;
  assign T750 = T751;
  assign T751 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T752 = T753;
  assign T753 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T754 = T755;
  assign T755 = T756;
  assign T756 = T760[T757];
  assign T757 = T758;
  assign T758 = T759;
  assign T759 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T760 = T761;
  assign T761 = io_chanxy_in[8'hec/* 236*/:8'heb/* 235*/];
  assign T762 = T763;
  assign T763 = T764;
  assign T764 = T768[T765];
  assign T765 = T766;
  assign T766 = T767;
  assign T767 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T768 = T769;
  assign T769 = io_chanxy_in[8'hf6/* 246*/:8'hed/* 237*/];
  assign T770 = T771;
  assign T771 = T772;
  assign T772 = T776[T773];
  assign T773 = T774;
  assign T774 = T775;
  assign T775 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T776 = T777;
  assign T777 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T778 = T779;
  assign T779 = T780;
  assign T780 = T784[T781];
  assign T781 = T782;
  assign T782 = T783;
  assign T783 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T784 = T785;
  assign T785 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T786 = T787;
  assign T787 = T788;
  assign T788 = T792[T789];
  assign T789 = T790;
  assign T790 = T791;
  assign T791 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T792 = T793;
  assign T793 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T794 = T795;
  assign T795 = T796;
  assign T796 = T800[T797];
  assign T797 = T798;
  assign T798 = T799;
  assign T799 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T800 = T801;
  assign T801 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T802 = T803;
  assign T803 = T804;
  assign T804 = T808[T805];
  assign T805 = T806;
  assign T806 = T807;
  assign T807 = io_chanxy_config[7'h7e/* 126*/:7'h7b/* 123*/];
  assign T808 = T809;
  assign T809 = io_chanxy_in[9'h108/* 264*/:8'hff/* 255*/];
  assign T810 = T811;
  assign T811 = T812;
  assign T812 = T816[T813];
  assign T813 = T814;
  assign T814 = T815;
  assign T815 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T816 = T817;
  assign T817 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T818 = T819;
  assign T819 = T820;
  assign T820 = T824[T821];
  assign T821 = T822;
  assign T822 = T823;
  assign T823 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T824 = T825;
  assign T825 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T826 = T827;
  assign T827 = T828;
  assign T828 = T832[T829];
  assign T829 = T830;
  assign T830 = T831;
  assign T831 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T832 = T833;
  assign T833 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T834 = T835;
  assign T835 = T836;
  assign T836 = T840[T837];
  assign T837 = T838;
  assign T838 = T839;
  assign T839 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T840 = T841;
  assign T841 = io_chanxy_in[9'h110/* 272*/:9'h10f/* 271*/];
  assign T842 = T843;
  assign T843 = T844;
  assign T844 = T848[T845];
  assign T845 = T846;
  assign T846 = T847;
  assign T847 = io_chanxy_config[8'h86/* 134*/:8'h83/* 131*/];
  assign T848 = T849;
  assign T849 = io_chanxy_in[9'h11a/* 282*/:9'h111/* 273*/];
  assign T850 = T851;
  assign T851 = T852;
  assign T852 = T856[T853];
  assign T853 = T854;
  assign T854 = T855;
  assign T855 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T856 = T857;
  assign T857 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T858 = T859;
  assign T859 = T860;
  assign T860 = T864[T861];
  assign T861 = T862;
  assign T862 = T863;
  assign T863 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T864 = T865;
  assign T865 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T866 = T867;
  assign T867 = T868;
  assign T868 = T872[T869];
  assign T869 = T870;
  assign T870 = T871;
  assign T871 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T872 = T873;
  assign T873 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T874 = T875;
  assign T875 = T876;
  assign T876 = T880[T877];
  assign T877 = T878;
  assign T878 = T879;
  assign T879 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T880 = T881;
  assign T881 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T882 = T883;
  assign T883 = T884;
  assign T884 = T888[T885];
  assign T885 = T886;
  assign T886 = T887;
  assign T887 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T888 = T889;
  assign T889 = io_chanxy_in[9'h12c/* 300*/:9'h123/* 291*/];
  assign T890 = T891;
  assign T891 = T892;
  assign T892 = T896[T893];
  assign T893 = T894;
  assign T894 = T895;
  assign T895 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T896 = T897;
  assign T897 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T898 = T899;
  assign T899 = T900;
  assign T900 = T904[T901];
  assign T901 = T902;
  assign T902 = T903;
  assign T903 = io_chanxy_config[8'h91/* 145*/:8'h90/* 144*/];
  assign T904 = T905;
  assign T905 = io_chanxy_in[9'h131/* 305*/:9'h12f/* 303*/];
  assign T906 = T907;
  assign T907 = T908;
  assign T908 = T912[T909];
  assign T909 = T910;
  assign T910 = T911;
  assign T911 = io_chanxy_config[8'h93/* 147*/:8'h92/* 146*/];
  assign T912 = T913;
  assign T913 = io_chanxy_in[9'h134/* 308*/:9'h132/* 306*/];
  assign T914 = T915;
  assign T915 = T916;
  assign T916 = T920[T917];
  assign T917 = T918;
  assign T918 = T919;
  assign T919 = io_chanxy_config[8'h95/* 149*/:8'h94/* 148*/];
  assign T920 = T921;
  assign T921 = io_chanxy_in[9'h137/* 311*/:9'h135/* 309*/];
  assign T922 = T923;
  assign T923 = T924;
  assign T924 = T928[T925];
  assign T925 = T926;
  assign T926 = T927;
  assign T927 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T928 = T929;
  assign T929 = io_chanxy_in[9'h142/* 322*/:9'h138/* 312*/];
  assign T930 = T931;
  assign T931 = T932;
  assign T932 = T936[T933];
  assign T933 = T934;
  assign T934 = T935;
  assign T935 = io_chanxy_config[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T936 = T937;
  assign T937 = io_chanxy_in[9'h145/* 325*/:9'h143/* 323*/];
  assign T938 = T939;
  assign T939 = T940;
  assign T940 = T944[T941];
  assign T941 = T942;
  assign T942 = T943;
  assign T943 = io_chanxy_config[8'h9d/* 157*/:8'h9c/* 156*/];
  assign T944 = T945;
  assign T945 = io_chanxy_in[9'h148/* 328*/:9'h146/* 326*/];
  assign T946 = T947;
  assign T947 = T948;
  assign T948 = T952[T949];
  assign T949 = T950;
  assign T950 = T951;
  assign T951 = io_chanxy_config[8'h9f/* 159*/:8'h9e/* 158*/];
  assign T952 = T953;
  assign T953 = io_chanxy_in[9'h14b/* 331*/:9'h149/* 329*/];
  assign T954 = T955;
  assign T955 = T956;
  assign T956 = T960[T957];
  assign T957 = T958;
  assign T958 = T959;
  assign T959 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T960 = T961;
  assign T961 = io_chanxy_in[9'h14e/* 334*/:9'h14c/* 332*/];
  assign T962 = T963;
  assign T963 = T964;
  assign T964 = T968[T965];
  assign T965 = T966;
  assign T966 = T967;
  assign T967 = io_chanxy_config[8'ha5/* 165*/:8'ha2/* 162*/];
  assign T968 = T969;
  assign T969 = io_chanxy_in[9'h159/* 345*/:9'h14f/* 335*/];
  assign T970 = T971;
  assign T971 = T972;
  assign T972 = T976[T973];
  assign T973 = T974;
  assign T974 = T975;
  assign T975 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T976 = T977;
  assign T977 = io_chanxy_in[9'h15c/* 348*/:9'h15a/* 346*/];
  assign T978 = T979;
  assign T979 = T980;
  assign T980 = T984[T981];
  assign T981 = T982;
  assign T982 = T983;
  assign T983 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T984 = T985;
  assign T985 = io_chanxy_in[9'h15f/* 351*/:9'h15d/* 349*/];
  assign T986 = T987;
  assign T987 = T988;
  assign T988 = T992[T989];
  assign T989 = T990;
  assign T990 = T991;
  assign T991 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T992 = T993;
  assign T993 = io_chanxy_in[9'h162/* 354*/:9'h160/* 352*/];
  assign T994 = T995;
  assign T995 = T996;
  assign T996 = T1000[T997];
  assign T997 = T998;
  assign T998 = T999;
  assign T999 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T1000 = T1001;
  assign T1001 = io_chanxy_in[9'h165/* 357*/:9'h163/* 355*/];
  assign T1002 = T1003;
  assign T1003 = T1004;
  assign T1004 = T1008[T1005];
  assign T1005 = T1006;
  assign T1006 = T1007;
  assign T1007 = io_chanxy_config[8'hb1/* 177*/:8'hae/* 174*/];
  assign T1008 = T1009;
  assign T1009 = io_chanxy_in[9'h170/* 368*/:9'h166/* 358*/];
  assign T1010 = T1011;
  assign T1011 = T1012;
  assign T1012 = T1016[T1013];
  assign T1013 = T1014;
  assign T1014 = T1015;
  assign T1015 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T1016 = T1017;
  assign T1017 = io_chanxy_in[9'h173/* 371*/:9'h171/* 369*/];
  assign T1018 = T1019;
  assign T1019 = T1020;
  assign T1020 = T1024[T1021];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T1024 = T1025;
  assign T1025 = io_chanxy_in[9'h176/* 374*/:9'h174/* 372*/];
  assign T1026 = T1027;
  assign T1027 = T1028;
  assign T1028 = T1032[T1029];
  assign T1029 = T1030;
  assign T1030 = T1031;
  assign T1031 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T1032 = T1033;
  assign T1033 = io_chanxy_in[9'h179/* 377*/:9'h177/* 375*/];
  assign T1034 = T1035;
  assign T1035 = T1036;
  assign T1036 = T1040[T1037];
  assign T1037 = T1038;
  assign T1038 = T1039;
  assign T1039 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T1040 = T1041;
  assign T1041 = io_chanxy_in[9'h17c/* 380*/:9'h17a/* 378*/];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = T1048[T1045];
  assign T1045 = T1046;
  assign T1046 = T1047;
  assign T1047 = io_chanxy_config[8'hbd/* 189*/:8'hba/* 186*/];
  assign T1048 = T1049;
  assign T1049 = io_chanxy_in[9'h187/* 391*/:9'h17d/* 381*/];
  assign T1050 = T1051;
  assign T1051 = T1052;
  assign T1052 = T1056[T1053];
  assign T1053 = T1054;
  assign T1054 = T1055;
  assign T1055 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T1056 = T1057;
  assign T1057 = io_chanxy_in[9'h18a/* 394*/:9'h188/* 392*/];
  assign T1058 = T1059;
  assign T1059 = T1060;
  assign T1060 = T1064[T1061];
  assign T1061 = T1062;
  assign T1062 = T1063;
  assign T1063 = io_chanxy_config[8'hc1/* 193*/:8'hc0/* 192*/];
  assign T1064 = T1065;
  assign T1065 = io_chanxy_in[9'h18d/* 397*/:9'h18b/* 395*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1072[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = io_chanxy_config[8'hc3/* 195*/:8'hc2/* 194*/];
  assign T1072 = T1073;
  assign T1073 = io_chanxy_in[9'h190/* 400*/:9'h18e/* 398*/];
  assign T1074 = T1075;
  assign T1075 = T1076;
  assign T1076 = T1080[T1077];
  assign T1077 = T1078;
  assign T1078 = T1079;
  assign T1079 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T1080 = T1081;
  assign T1081 = io_chanxy_in[9'h193/* 403*/:9'h191/* 401*/];
  assign T1082 = T1083;
  assign T1083 = T1084;
  assign T1084 = T1088[T1085];
  assign T1085 = T1086;
  assign T1086 = T1087;
  assign T1087 = io_chanxy_config[8'hc9/* 201*/:8'hc6/* 198*/];
  assign T1088 = T1089;
  assign T1089 = io_chanxy_in[9'h19e/* 414*/:9'h194/* 404*/];
  assign T1090 = T1091;
  assign T1091 = T1092;
  assign T1092 = T1096[T1093];
  assign T1093 = T1094;
  assign T1094 = T1095;
  assign T1095 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T1096 = T1097;
  assign T1097 = io_chanxy_in[9'h1a1/* 417*/:9'h19f/* 415*/];
  assign T1098 = T1099;
  assign T1099 = T1100;
  assign T1100 = T1104[T1101];
  assign T1101 = T1102;
  assign T1102 = T1103;
  assign T1103 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T1104 = T1105;
  assign T1105 = io_chanxy_in[9'h1a4/* 420*/:9'h1a2/* 418*/];
  assign T1106 = T1107;
  assign T1107 = T1108;
  assign T1108 = T1112[T1109];
  assign T1109 = T1110;
  assign T1110 = T1111;
  assign T1111 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T1112 = T1113;
  assign T1113 = io_chanxy_in[9'h1a7/* 423*/:9'h1a5/* 421*/];
  assign T1114 = T1115;
  assign T1115 = T1116;
  assign T1116 = T1120[T1117];
  assign T1117 = T1118;
  assign T1118 = T1119;
  assign T1119 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T1120 = T1121;
  assign T1121 = io_chanxy_in[9'h1aa/* 426*/:9'h1a8/* 424*/];
  assign T1122 = T1123;
  assign T1123 = T1124;
  assign T1124 = T1128[T1125];
  assign T1125 = T1126;
  assign T1126 = T1127;
  assign T1127 = io_chanxy_config[8'hd5/* 213*/:8'hd2/* 210*/];
  assign T1128 = T1129;
  assign T1129 = io_chanxy_in[9'h1b5/* 437*/:9'h1ab/* 427*/];
  assign T1130 = T1131;
  assign T1131 = T1132;
  assign T1132 = T1136[T1133];
  assign T1133 = T1134;
  assign T1134 = T1135;
  assign T1135 = io_chanxy_config[8'hd7/* 215*/:8'hd6/* 214*/];
  assign T1136 = T1137;
  assign T1137 = io_chanxy_in[9'h1b8/* 440*/:9'h1b6/* 438*/];
  assign T1138 = T1139;
  assign T1139 = T1140;
  assign T1140 = T1144[T1141];
  assign T1141 = T1142;
  assign T1142 = T1143;
  assign T1143 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T1144 = T1145;
  assign T1145 = io_chanxy_in[9'h1ba/* 442*/:9'h1b9/* 441*/];
  assign T1146 = T1147;
  assign T1147 = T1148;
  assign T1148 = T1152[T1149];
  assign T1149 = T1150;
  assign T1150 = T1151;
  assign T1151 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T1152 = T1153;
  assign T1153 = io_chanxy_in[9'h1bc/* 444*/:9'h1bb/* 443*/];
  assign T1154 = T1155;
  assign T1155 = T1156;
  assign T1156 = T1160[T1157];
  assign T1157 = T1158;
  assign T1158 = T1159;
  assign T1159 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T1160 = T1161;
  assign T1161 = io_chanxy_in[9'h1be/* 446*/:9'h1bd/* 445*/];
  assign T1162 = T1163;
  assign T1163 = T1164;
  assign T1164 = T1168[T1165];
  assign T1165 = T1166;
  assign T1166 = T1167;
  assign T1167 = io_chanxy_config[8'hde/* 222*/:8'hdb/* 219*/];
  assign T1168 = T1169;
  assign T1169 = io_chanxy_in[9'h1c9/* 457*/:9'h1bf/* 447*/];
  assign T1170 = T1171;
  assign T1171 = T1172;
  assign T1172 = T1176[T1173];
  assign T1173 = T1174;
  assign T1174 = T1175;
  assign T1175 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T1176 = T1177;
  assign T1177 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T1178 = T1179;
  assign T1179 = T1180;
  assign T1180 = T1184[T1181];
  assign T1181 = T1182;
  assign T1182 = T1183;
  assign T1183 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T1184 = T1185;
  assign T1185 = io_chanxy_in[9'h1cd/* 461*/:9'h1cc/* 460*/];
  assign T1186 = T1187;
  assign T1187 = T1188;
  assign T1188 = T1192[T1189];
  assign T1189 = T1190;
  assign T1190 = T1191;
  assign T1191 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T1192 = T1193;
  assign T1193 = io_chanxy_in[9'h1cf/* 463*/:9'h1ce/* 462*/];
  assign T1194 = T1195;
  assign T1195 = T1196;
  assign T1196 = T1200[T1197];
  assign T1197 = T1198;
  assign T1198 = T1199;
  assign T1199 = io_chanxy_config[8'he2/* 226*/:8'he2/* 226*/];
  assign T1200 = T1201;
  assign T1201 = io_chanxy_in[9'h1d1/* 465*/:9'h1d0/* 464*/];
  assign T1202 = T1203;
  assign T1203 = T1204;
  assign T1204 = T1208[T1205];
  assign T1205 = T1206;
  assign T1206 = T1207;
  assign T1207 = io_chanxy_config[8'he6/* 230*/:8'he3/* 227*/];
  assign T1208 = T1209;
  assign T1209 = io_chanxy_in[9'h1dc/* 476*/:9'h1d2/* 466*/];
  assign T1210 = T1211;
  assign T1211 = T1212;
  assign T1212 = T1216[T1213];
  assign T1213 = T1214;
  assign T1214 = T1215;
  assign T1215 = io_chanxy_config[8'he7/* 231*/:8'he7/* 231*/];
  assign T1216 = T1217;
  assign T1217 = io_chanxy_in[9'h1de/* 478*/:9'h1dd/* 477*/];
  assign T1218 = T1219;
  assign T1219 = T1220;
  assign T1220 = T1224[T1221];
  assign T1221 = T1222;
  assign T1222 = T1223;
  assign T1223 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T1224 = T1225;
  assign T1225 = io_chanxy_in[9'h1e0/* 480*/:9'h1df/* 479*/];
  assign T1226 = T1227;
  assign T1227 = T1228;
  assign T1228 = T1232[T1229];
  assign T1229 = T1230;
  assign T1230 = T1231;
  assign T1231 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T1232 = T1233;
  assign T1233 = io_chanxy_in[9'h1e2/* 482*/:9'h1e1/* 481*/];
  assign T1234 = T1235;
  assign T1235 = T1236;
  assign T1236 = T1240[T1237];
  assign T1237 = T1238;
  assign T1238 = T1239;
  assign T1239 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T1240 = T1241;
  assign T1241 = io_chanxy_in[9'h1e4/* 484*/:9'h1e3/* 483*/];
  assign T1242 = T1243;
  assign T1243 = T1244;
  assign T1244 = T1248[T1245];
  assign T1245 = T1246;
  assign T1246 = T1247;
  assign T1247 = io_chanxy_config[8'hee/* 238*/:8'heb/* 235*/];
  assign T1248 = T1249;
  assign T1249 = io_chanxy_in[9'h1ef/* 495*/:9'h1e5/* 485*/];
  assign T1250 = T1251;
  assign T1251 = T1252;
  assign T1252 = T1256[T1253];
  assign T1253 = T1254;
  assign T1254 = T1255;
  assign T1255 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T1256 = T1257;
  assign T1257 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T1258 = T1259;
  assign T1259 = T1260;
  assign T1260 = T1264[T1261];
  assign T1261 = T1262;
  assign T1262 = T1263;
  assign T1263 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T1264 = T1265;
  assign T1265 = io_chanxy_in[9'h1f3/* 499*/:9'h1f2/* 498*/];
  assign T1266 = T1267;
  assign T1267 = T1268;
  assign T1268 = T1272[T1269];
  assign T1269 = T1270;
  assign T1270 = T1271;
  assign T1271 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T1272 = T1273;
  assign T1273 = io_chanxy_in[9'h1f5/* 501*/:9'h1f4/* 500*/];
  assign T1274 = T1275;
  assign T1275 = T1276;
  assign T1276 = T1280[T1277];
  assign T1277 = T1278;
  assign T1278 = T1279;
  assign T1279 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1280 = T1281;
  assign T1281 = io_chanxy_in[9'h1f7/* 503*/:9'h1f6/* 502*/];
  assign T1282 = T1283;
  assign T1283 = T1284;
  assign T1284 = T1288[T1285];
  assign T1285 = T1286;
  assign T1286 = T1287;
  assign T1287 = io_chanxy_config[8'hf6/* 246*/:8'hf3/* 243*/];
  assign T1288 = T1289;
  assign T1289 = io_chanxy_in[10'h201/* 513*/:9'h1f8/* 504*/];
  assign T1290 = T1291;
  assign T1291 = T1292;
  assign T1292 = T1296[T1293];
  assign T1293 = T1294;
  assign T1294 = T1295;
  assign T1295 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T1296 = T1297;
  assign T1297 = io_chanxy_in[10'h203/* 515*/:10'h202/* 514*/];
  assign T1298 = T1299;
  assign T1299 = T1300;
  assign T1300 = T1304[T1301];
  assign T1301 = T1302;
  assign T1302 = T1303;
  assign T1303 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1304 = T1305;
  assign T1305 = io_chanxy_in[10'h205/* 517*/:10'h204/* 516*/];
  assign T1306 = T1307;
  assign T1307 = T1308;
  assign T1308 = T1312[T1309];
  assign T1309 = T1310;
  assign T1310 = T1311;
  assign T1311 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T1312 = T1313;
  assign T1313 = io_chanxy_in[10'h207/* 519*/:10'h206/* 518*/];
  assign T1314 = T1315;
  assign T1315 = T1316;
  assign T1316 = T1320[T1317];
  assign T1317 = T1318;
  assign T1318 = T1319;
  assign T1319 = io_chanxy_config[8'hfa/* 250*/:8'hfa/* 250*/];
  assign T1320 = T1321;
  assign T1321 = io_chanxy_in[10'h209/* 521*/:10'h208/* 520*/];
  assign T1322 = T1323;
  assign T1323 = T1324;
  assign T1324 = T1328[T1325];
  assign T1325 = T1326;
  assign T1326 = T1327;
  assign T1327 = io_chanxy_config[8'hfe/* 254*/:8'hfb/* 251*/];
  assign T1328 = T1329;
  assign T1329 = io_chanxy_in[10'h213/* 531*/:10'h20a/* 522*/];
  assign T1330 = T1331;
  assign T1331 = T1332;
  assign T1332 = T1336[T1333];
  assign T1333 = T1334;
  assign T1334 = T1335;
  assign T1335 = io_chanxy_config[8'hff/* 255*/:8'hff/* 255*/];
  assign T1336 = T1337;
  assign T1337 = io_chanxy_in[10'h215/* 533*/:10'h214/* 532*/];
  assign T1338 = T1339;
  assign T1339 = T1340;
  assign T1340 = T1344[T1341];
  assign T1341 = T1342;
  assign T1342 = T1343;
  assign T1343 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1344 = T1345;
  assign T1345 = io_chanxy_in[10'h217/* 535*/:10'h216/* 534*/];
  assign T1346 = T1347;
  assign T1347 = T1348;
  assign T1348 = T1352[T1349];
  assign T1349 = T1350;
  assign T1350 = T1351;
  assign T1351 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1352 = T1353;
  assign T1353 = io_chanxy_in[10'h219/* 537*/:10'h218/* 536*/];
  assign T1354 = T1355;
  assign T1355 = T1356;
  assign T1356 = T1360[T1357];
  assign T1357 = T1358;
  assign T1358 = T1359;
  assign T1359 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1360 = T1361;
  assign T1361 = io_chanxy_in[10'h21b/* 539*/:10'h21a/* 538*/];
  assign T1362 = T1363;
  assign T1363 = T1364;
  assign T1364 = T1368[T1365];
  assign T1365 = T1366;
  assign T1366 = T1367;
  assign T1367 = io_chanxy_config[9'h106/* 262*/:9'h103/* 259*/];
  assign T1368 = T1369;
  assign T1369 = io_chanxy_in[10'h225/* 549*/:10'h21c/* 540*/];
  assign T1370 = T1371;
  assign T1371 = T1372;
  assign T1372 = T1376[T1373];
  assign T1373 = T1374;
  assign T1374 = T1375;
  assign T1375 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1376 = T1377;
  assign T1377 = io_chanxy_in[10'h227/* 551*/:10'h226/* 550*/];
  assign T1378 = T1379;
  assign T1379 = T1380;
  assign T1380 = T1384[T1381];
  assign T1381 = T1382;
  assign T1382 = T1383;
  assign T1383 = io_chanxy_config[9'h108/* 264*/:9'h108/* 264*/];
  assign T1384 = T1385;
  assign T1385 = io_chanxy_in[10'h229/* 553*/:10'h228/* 552*/];
  assign T1386 = T1387;
  assign T1387 = T1388;
  assign T1388 = T1392[T1389];
  assign T1389 = T1390;
  assign T1390 = T1391;
  assign T1391 = io_chanxy_config[9'h109/* 265*/:9'h109/* 265*/];
  assign T1392 = T1393;
  assign T1393 = io_chanxy_in[10'h22b/* 555*/:10'h22a/* 554*/];
  assign T1394 = T1395;
  assign T1395 = T1396;
  assign T1396 = T1400[T1397];
  assign T1397 = T1398;
  assign T1398 = T1399;
  assign T1399 = io_chanxy_config[9'h10a/* 266*/:9'h10a/* 266*/];
  assign T1400 = T1401;
  assign T1401 = io_chanxy_in[10'h22d/* 557*/:10'h22c/* 556*/];
  assign T1402 = T1403;
  assign T1403 = T1404;
  assign T1404 = T1408[T1405];
  assign T1405 = T1406;
  assign T1406 = T1407;
  assign T1407 = io_chanxy_config[9'h10e/* 270*/:9'h10b/* 267*/];
  assign T1408 = T1409;
  assign T1409 = io_chanxy_in[10'h237/* 567*/:10'h22e/* 558*/];
  assign T1410 = T1411;
  assign T1411 = T1412;
  assign T1412 = T1416[T1413];
  assign T1413 = T1414;
  assign T1414 = T1415;
  assign T1415 = io_chanxy_config[9'h10f/* 271*/:9'h10f/* 271*/];
  assign T1416 = T1417;
  assign T1417 = io_chanxy_in[10'h239/* 569*/:10'h238/* 568*/];
  assign T1418 = T1419;
  assign T1419 = T1420;
  assign T1420 = T1424[T1421];
  assign T1421 = T1422;
  assign T1422 = T1423;
  assign T1423 = io_chanxy_config[9'h110/* 272*/:9'h110/* 272*/];
  assign T1424 = T1425;
  assign T1425 = io_chanxy_in[10'h23b/* 571*/:10'h23a/* 570*/];
  assign T1426 = T1427;
  assign T1427 = T1428;
  assign T1428 = T1432[T1429];
  assign T1429 = T1430;
  assign T1430 = T1431;
  assign T1431 = io_chanxy_config[9'h111/* 273*/:9'h111/* 273*/];
  assign T1432 = T1433;
  assign T1433 = io_chanxy_in[10'h23d/* 573*/:10'h23c/* 572*/];
  assign T1434 = T1435;
  assign T1435 = T1436;
  assign T1436 = T1440[T1437];
  assign T1437 = T1438;
  assign T1438 = T1439;
  assign T1439 = io_chanxy_config[9'h112/* 274*/:9'h112/* 274*/];
  assign T1440 = T1441;
  assign T1441 = io_chanxy_in[10'h23f/* 575*/:10'h23e/* 574*/];
  assign T1442 = T1443;
  assign T1443 = T1444;
  assign T1444 = T1448[T1445];
  assign T1445 = T1446;
  assign T1446 = T1447;
  assign T1447 = io_chanxy_config[9'h116/* 278*/:9'h113/* 275*/];
  assign T1448 = T1449;
  assign T1449 = io_chanxy_in[10'h249/* 585*/:10'h240/* 576*/];
  assign T1450 = T1451;
  assign T1451 = T1452;
  assign T1452 = T1456[T1453];
  assign T1453 = T1454;
  assign T1454 = T1455;
  assign T1455 = io_chanxy_config[9'h117/* 279*/:9'h117/* 279*/];
  assign T1456 = T1457;
  assign T1457 = io_chanxy_in[10'h24b/* 587*/:10'h24a/* 586*/];
  assign T1458 = T1459;
  assign T1459 = T1460;
  assign T1460 = T1464[T1461];
  assign T1461 = T1462;
  assign T1462 = T1463;
  assign T1463 = io_chanxy_config[9'h118/* 280*/:9'h118/* 280*/];
  assign T1464 = T1465;
  assign T1465 = io_chanxy_in[10'h24d/* 589*/:10'h24c/* 588*/];
  assign T1466 = T1467;
  assign T1467 = T1468;
  assign T1468 = T1472[T1469];
  assign T1469 = T1470;
  assign T1470 = T1471;
  assign T1471 = io_chanxy_config[9'h119/* 281*/:9'h119/* 281*/];
  assign T1472 = T1473;
  assign T1473 = io_chanxy_in[10'h24f/* 591*/:10'h24e/* 590*/];
  assign T1474 = T1475;
  assign T1475 = T1476;
  assign T1476 = T1480[T1477];
  assign T1477 = T1478;
  assign T1478 = T1479;
  assign T1479 = io_chanxy_config[9'h11a/* 282*/:9'h11a/* 282*/];
  assign T1480 = T1481;
  assign T1481 = io_chanxy_in[10'h251/* 593*/:10'h250/* 592*/];
  assign T1482 = T1483;
  assign T1483 = T1484;
  assign T1484 = T1488[T1485];
  assign T1485 = T1486;
  assign T1486 = T1487;
  assign T1487 = io_chanxy_config[9'h11e/* 286*/:9'h11b/* 283*/];
  assign T1488 = T1489;
  assign T1489 = io_chanxy_in[10'h25b/* 603*/:10'h252/* 594*/];
  assign T1490 = T1491;
  assign T1491 = T1492;
  assign T1492 = T1496[T1493];
  assign T1493 = T1494;
  assign T1494 = T1495;
  assign T1495 = io_chanxy_config[9'h11f/* 287*/:9'h11f/* 287*/];
  assign T1496 = T1497;
  assign T1497 = io_chanxy_in[10'h25d/* 605*/:10'h25c/* 604*/];
  assign io_ipin_out = T1498;
  assign T1498 = T1499;
  assign T1499 = {T1718, T1500};
  assign T1500 = T1501;
  assign T1501 = {T1710, T1502};
  assign T1502 = T1503;
  assign T1503 = {T1702, T1504};
  assign T1504 = T1505;
  assign T1505 = {T1694, T1506};
  assign T1506 = T1507;
  assign T1507 = {T1686, T1508};
  assign T1508 = T1509;
  assign T1509 = {T1678, T1510};
  assign T1510 = T1511;
  assign T1511 = {T1670, T1512};
  assign T1512 = T1513;
  assign T1513 = {T1662, T1514};
  assign T1514 = T1515;
  assign T1515 = {T1654, T1516};
  assign T1516 = T1517;
  assign T1517 = {T1646, T1518};
  assign T1518 = T1519;
  assign T1519 = {T1638, T1520};
  assign T1520 = T1521;
  assign T1521 = {T1630, T1522};
  assign T1522 = T1523;
  assign T1523 = {T1622, T1524};
  assign T1524 = T1525;
  assign T1525 = {T1614, T1526};
  assign T1526 = T1527;
  assign T1527 = {T1606, T1528};
  assign T1528 = T1529;
  assign T1529 = {T1598, T1530};
  assign T1530 = T1531;
  assign T1531 = {T1590, T1532};
  assign T1532 = T1533;
  assign T1533 = {T1582, T1534};
  assign T1534 = T1535;
  assign T1535 = {T1574, T1536};
  assign T1536 = T1537;
  assign T1537 = {T1566, T1538};
  assign T1538 = T1539;
  assign T1539 = {T1558, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1550, T1542};
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_0(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [26:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [605:0] io_chanxy_in,
    output[149:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[287:0] T0;
  wire[863:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[149:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h34b/* 843*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_27 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


module sbcb_sp_1(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[1:0] T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[1:0] T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[1:0] T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire[2:0] T230;
  wire[2:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire[2:0] T238;
  wire[2:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[10:0] T246;
  wire[10:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  wire[1:0] T260;
  wire[1:0] T261;
  wire[2:0] T262;
  wire[2:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire[2:0] T270;
  wire[2:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[1:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire[2:0] T278;
  wire[2:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[10:0] T286;
  wire[10:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[1:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[2:0] T302;
  wire[2:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[1:0] T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire[2:0] T310;
  wire[2:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[1:0] T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire[2:0] T318;
  wire[2:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[10:0] T326;
  wire[10:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[1:0] T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[1:0] T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[1:0] T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire[2:0] T350;
  wire[2:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[10:0] T366;
  wire[10:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire[2:0] T398;
  wire[2:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[10:0] T406;
  wire[10:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[1:0] T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire[2:0] T414;
  wire[2:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[1:0] T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire[2:0] T422;
  wire[2:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[2:0] T430;
  wire[2:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[2:0] T438;
  wire[2:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[10:0] T446;
  wire[10:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire[1:0] T462;
  wire[1:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire[1:0] T470;
  wire[1:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire[1:0] T478;
  wire[1:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[3:0] T483;
  wire[3:0] T484;
  wire[3:0] T485;
  wire[10:0] T486;
  wire[10:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire[1:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire[3:0] T523;
  wire[3:0] T524;
  wire[3:0] T525;
  wire[10:0] T526;
  wire[10:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[3:0] T563;
  wire[3:0] T564;
  wire[3:0] T565;
  wire[10:0] T566;
  wire[10:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire[1:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire[1:0] T582;
  wire[1:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire[1:0] T598;
  wire[1:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[3:0] T603;
  wire[3:0] T604;
  wire[3:0] T605;
  wire[9:0] T606;
  wire[9:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[1:0] T614;
  wire[1:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[1:0] T622;
  wire[1:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire[1:0] T638;
  wire[1:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[3:0] T643;
  wire[3:0] T644;
  wire[3:0] T645;
  wire[9:0] T646;
  wire[9:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire[1:0] T654;
  wire[1:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire[1:0] T662;
  wire[1:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[1:0] T678;
  wire[1:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[3:0] T683;
  wire[3:0] T684;
  wire[3:0] T685;
  wire[9:0] T686;
  wire[9:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire[3:0] T723;
  wire[3:0] T724;
  wire[3:0] T725;
  wire[9:0] T726;
  wire[9:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire[3:0] T763;
  wire[3:0] T764;
  wire[3:0] T765;
  wire[9:0] T766;
  wire[9:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire[3:0] T803;
  wire[3:0] T804;
  wire[3:0] T805;
  wire[9:0] T806;
  wire[9:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[10:0] T814;
  wire[10:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[10:0] T822;
  wire[10:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[10:0] T830;
  wire[10:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[10:0] T838;
  wire[10:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[10:0] T846;
  wire[10:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[3:0] T851;
  wire[3:0] T852;
  wire[3:0] T853;
  wire[10:0] T854;
  wire[10:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[10:0] T862;
  wire[10:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[10:0] T870;
  wire[10:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[10:0] T878;
  wire[10:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[9:0] T886;
  wire[9:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[9:0] T894;
  wire[9:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[9:0] T902;
  wire[9:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[9:0] T910;
  wire[9:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[9:0] T918;
  wire[9:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[3:0] T932;
  wire[3:0] T933;
  wire[10:0] T934;
  wire[10:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[10:0] T942;
  wire[10:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[10:0] T950;
  wire[10:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[10:0] T958;
  wire[10:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[10:0] T966;
  wire[10:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[10:0] T974;
  wire[10:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[10:0] T982;
  wire[10:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[10:0] T990;
  wire[10:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[10:0] T998;
  wire[10:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire[3:0] T1011;
  wire[3:0] T1012;
  wire[3:0] T1013;
  wire[9:0] T1014;
  wire[9:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[9:0] T1030;
  wire[9:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[9:0] T1046;
  wire[9:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[5'h16/* 22*/:4'hc/* 12*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[5'h1f/* 31*/:5'h1d/* 29*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[6'h22/* 34*/:6'h20/* 32*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[6'h2d/* 45*/:6'h23/* 35*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[6'h36/* 54*/:6'h34/* 52*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[6'h39/* 57*/:6'h37/* 55*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[7'h44/* 68*/:6'h3a/* 58*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[7'h50/* 80*/:7'h4e/* 78*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[7'h5b/* 91*/:7'h51/* 81*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[7'h64/* 100*/:7'h62/* 98*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[6'h37/* 55*/:6'h36/* 54*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[7'h67/* 103*/:7'h65/* 101*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[7'h72/* 114*/:7'h68/* 104*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[7'h7e/* 126*/:7'h7c/* 124*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[8'h89/* 137*/:7'h7f/* 127*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h4b/* 75*/:7'h4b/* 75*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[8'h91/* 145*/:8'h90/* 144*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[8'h9c/* 156*/:8'h92/* 146*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[8'ha0/* 160*/:8'h9f/* 159*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[8'ha2/* 162*/:8'ha1/* 161*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[7'h53/* 83*/:7'h53/* 83*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[8'ha4/* 164*/:8'ha3/* 163*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[8'haf/* 175*/:8'ha5/* 165*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[7'h5a/* 90*/:7'h5a/* 90*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[7'h5b/* 91*/:7'h5b/* 91*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[8'hc2/* 194*/:8'hb8/* 184*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[8'hc6/* 198*/:8'hc5/* 197*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[7'h62/* 98*/:7'h62/* 98*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[7'h63/* 99*/:7'h63/* 99*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[8'hca/* 202*/:8'hc9/* 201*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[8'hd4/* 212*/:8'hcb/* 203*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[8'hd6/* 214*/:8'hd5/* 213*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[8'hd8/* 216*/:8'hd7/* 215*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[7'h6a/* 106*/:7'h6a/* 106*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[7'h6b/* 107*/:7'h6b/* 107*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[8'hdc/* 220*/:8'hdb/* 219*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[8'he6/* 230*/:8'hdd/* 221*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[8'hec/* 236*/:8'heb/* 235*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[7'h73/* 115*/:7'h73/* 115*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[8'hee/* 238*/:8'hed/* 237*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[8'hf8/* 248*/:8'hef/* 239*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[7'h7b/* 123*/:7'h7b/* 123*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h10a/* 266*/:9'h101/* 257*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h110/* 272*/:9'h10f/* 271*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'h83/* 131*/:8'h83/* 131*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h112/* 274*/:9'h111/* 273*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h11c/* 284*/:9'h113/* 275*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h12e/* 302*/:9'h125/* 293*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h144/* 324*/:9'h13a/* 314*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h14f/* 335*/:9'h145/* 325*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h15a/* 346*/:9'h150/* 336*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h165/* 357*/:9'h15b/* 347*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h170/* 368*/:9'h166/* 358*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h17b/* 379*/:9'h171/* 369*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h186/* 390*/:9'h17c/* 380*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h191/* 401*/:9'h187/* 391*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h19b/* 411*/:9'h192/* 402*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h1a5/* 421*/:9'h19c/* 412*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h1af/* 431*/:9'h1a6/* 422*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1b9/* 441*/:9'h1b0/* 432*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1c3/* 451*/:9'h1ba/* 442*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1cd/* 461*/:9'h1c4/* 452*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1e3/* 483*/:9'h1d9/* 473*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1ee/* 494*/:9'h1e4/* 484*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1f9/* 505*/:9'h1ef/* 495*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h204/* 516*/:9'h1fa/* 506*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h20f/* 527*/:10'h205/* 517*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h21a/* 538*/:10'h210/* 528*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h225/* 549*/:10'h21b/* 539*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h230/* 560*/:10'h226/* 550*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h23a/* 570*/:10'h231/* 561*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h244/* 580*/:10'h23b/* 571*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h24e/* 590*/:10'h245/* 581*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h258/* 600*/:10'h24f/* 591*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h262/* 610*/:10'h259/* 601*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h263/* 611*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_1(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_2(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[1:0] T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[10:0] T222;
  wire[10:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[1:0] T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire[2:0] T230;
  wire[2:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire[2:0] T238;
  wire[2:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire[2:0] T246;
  wire[2:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[10:0] T262;
  wire[10:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire[2:0] T270;
  wire[2:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[1:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire[2:0] T278;
  wire[2:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[1:0] T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire[2:0] T286;
  wire[2:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[10:0] T302;
  wire[10:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[1:0] T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire[2:0] T310;
  wire[2:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[1:0] T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire[2:0] T318;
  wire[2:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[2:0] T326;
  wire[2:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[1:0] T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[10:0] T342;
  wire[10:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[1:0] T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire[2:0] T350;
  wire[2:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[10:0] T382;
  wire[10:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire[2:0] T398;
  wire[2:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[1:0] T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire[2:0] T406;
  wire[2:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[1:0] T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire[2:0] T414;
  wire[2:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[10:0] T422;
  wire[10:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[2:0] T430;
  wire[2:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[2:0] T438;
  wire[2:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire[2:0] T446;
  wire[2:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[3:0] T459;
  wire[3:0] T460;
  wire[3:0] T461;
  wire[10:0] T462;
  wire[10:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire[1:0] T470;
  wire[1:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire[1:0] T478;
  wire[1:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire[1:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire[1:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire[3:0] T499;
  wire[3:0] T500;
  wire[3:0] T501;
  wire[10:0] T502;
  wire[10:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire[3:0] T539;
  wire[3:0] T540;
  wire[3:0] T541;
  wire[10:0] T542;
  wire[10:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire[1:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[3:0] T579;
  wire[3:0] T580;
  wire[3:0] T581;
  wire[9:0] T582;
  wire[9:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire[1:0] T598;
  wire[1:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire[1:0] T606;
  wire[1:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[1:0] T614;
  wire[1:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[3:0] T619;
  wire[3:0] T620;
  wire[3:0] T621;
  wire[9:0] T622;
  wire[9:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire[1:0] T638;
  wire[1:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire[1:0] T646;
  wire[1:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire[1:0] T654;
  wire[1:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[3:0] T659;
  wire[3:0] T660;
  wire[3:0] T661;
  wire[9:0] T662;
  wire[9:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[1:0] T678;
  wire[1:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire[1:0] T686;
  wire[1:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire[3:0] T699;
  wire[3:0] T700;
  wire[3:0] T701;
  wire[9:0] T702;
  wire[9:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire[3:0] T739;
  wire[3:0] T740;
  wire[3:0] T741;
  wire[9:0] T742;
  wire[9:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire[3:0] T779;
  wire[3:0] T780;
  wire[3:0] T781;
  wire[9:0] T782;
  wire[9:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[10:0] T814;
  wire[10:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[10:0] T822;
  wire[10:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[10:0] T830;
  wire[10:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[10:0] T838;
  wire[10:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[10:0] T846;
  wire[10:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[3:0] T851;
  wire[3:0] T852;
  wire[3:0] T853;
  wire[10:0] T854;
  wire[10:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[10:0] T862;
  wire[10:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[10:0] T870;
  wire[10:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[10:0] T878;
  wire[10:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[9:0] T886;
  wire[9:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[9:0] T894;
  wire[9:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[9:0] T902;
  wire[9:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[9:0] T910;
  wire[9:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[9:0] T918;
  wire[9:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[3:0] T932;
  wire[3:0] T933;
  wire[10:0] T934;
  wire[10:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[10:0] T942;
  wire[10:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[10:0] T950;
  wire[10:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[10:0] T958;
  wire[10:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[10:0] T966;
  wire[10:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[10:0] T974;
  wire[10:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[10:0] T982;
  wire[10:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[10:0] T990;
  wire[10:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[10:0] T998;
  wire[10:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire[3:0] T1011;
  wire[3:0] T1012;
  wire[3:0] T1013;
  wire[9:0] T1014;
  wire[9:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[9:0] T1030;
  wire[9:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[9:0] T1046;
  wire[9:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h5/* 5*/:2'h2/* 2*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[4'hd/* 13*/:2'h3/* 3*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[5'h10/* 16*/:4'he/* 14*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[5'h13/* 19*/:5'h11/* 17*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h11/* 17*/:4'he/* 14*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[6'h24/* 36*/:5'h1a/* 26*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[6'h27/* 39*/:6'h25/* 37*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[5'h15/* 21*/:5'h14/* 20*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[6'h2a/* 42*/:6'h28/* 40*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[5'h1d/* 29*/:5'h1a/* 26*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[6'h3b/* 59*/:6'h31/* 49*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[6'h3e/* 62*/:6'h3c/* 60*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[7'h41/* 65*/:6'h3f/* 63*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[6'h29/* 41*/:6'h26/* 38*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[7'h52/* 82*/:7'h48/* 72*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[7'h55/* 85*/:7'h53/* 83*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[7'h58/* 88*/:7'h56/* 86*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[6'h35/* 53*/:6'h32/* 50*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[7'h69/* 105*/:7'h5f/* 95*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[6'h37/* 55*/:6'h36/* 54*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[7'h6c/* 108*/:7'h6a/* 106*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[6'h39/* 57*/:6'h38/* 56*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h41/* 65*/:6'h3e/* 62*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[8'h80/* 128*/:7'h76/* 118*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[8'h83/* 131*/:8'h81/* 129*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[8'h86/* 134*/:8'h84/* 132*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h4c/* 76*/:7'h49/* 73*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[8'h96/* 150*/:8'h8c/* 140*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h4d/* 77*/:7'h4d/* 77*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[8'h98/* 152*/:8'h97/* 151*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h4e/* 78*/:7'h4e/* 78*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[8'h9a/* 154*/:8'h99/* 153*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[7'h54/* 84*/:7'h51/* 81*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[8'ha9/* 169*/:8'h9f/* 159*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[7'h55/* 85*/:7'h55/* 85*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[8'hab/* 171*/:8'haa/* 170*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[8'had/* 173*/:8'hac/* 172*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[7'h5c/* 92*/:7'h59/* 89*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[8'hbc/* 188*/:8'hb2/* 178*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[7'h5d/* 93*/:7'h5d/* 93*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[8'hbe/* 190*/:8'hbd/* 189*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[8'hc0/* 192*/:8'hbf/* 191*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[7'h64/* 100*/:7'h61/* 97*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[8'hce/* 206*/:8'hc5/* 197*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[7'h65/* 101*/:7'h65/* 101*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[8'hd0/* 208*/:8'hcf/* 207*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[7'h66/* 102*/:7'h66/* 102*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[8'hd2/* 210*/:8'hd1/* 209*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[8'hd6/* 214*/:8'hd5/* 213*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[7'h6c/* 108*/:7'h69/* 105*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[8'he0/* 224*/:8'hd7/* 215*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[7'h6d/* 109*/:7'h6d/* 109*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[8'he2/* 226*/:8'he1/* 225*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[7'h6e/* 110*/:7'h6e/* 110*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[8'he4/* 228*/:8'he3/* 227*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[7'h74/* 116*/:7'h71/* 113*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[8'hf2/* 242*/:8'he9/* 233*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[7'h75/* 117*/:7'h75/* 117*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[8'hf4/* 244*/:8'hf3/* 243*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[8'hf6/* 246*/:8'hf5/* 245*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[7'h7c/* 124*/:7'h79/* 121*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h104/* 260*/:8'hfb/* 251*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[7'h7d/* 125*/:7'h7d/* 125*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h106/* 262*/:9'h105/* 261*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h108/* 264*/:9'h107/* 263*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'h84/* 132*/:8'h81/* 129*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h116/* 278*/:9'h10d/* 269*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h118/* 280*/:9'h117/* 279*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h11a/* 282*/:9'h119/* 281*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'h8c/* 140*/:8'h89/* 137*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h128/* 296*/:9'h11f/* 287*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'h8d/* 141*/:8'h8d/* 141*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h12a/* 298*/:9'h129/* 297*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h12c/* 300*/:9'h12b/* 299*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h144/* 324*/:9'h13a/* 314*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h14f/* 335*/:9'h145/* 325*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h15a/* 346*/:9'h150/* 336*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h165/* 357*/:9'h15b/* 347*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h170/* 368*/:9'h166/* 358*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h17b/* 379*/:9'h171/* 369*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h186/* 390*/:9'h17c/* 380*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h191/* 401*/:9'h187/* 391*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h19b/* 411*/:9'h192/* 402*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h1a5/* 421*/:9'h19c/* 412*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h1af/* 431*/:9'h1a6/* 422*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1b9/* 441*/:9'h1b0/* 432*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1c3/* 451*/:9'h1ba/* 442*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1cd/* 461*/:9'h1c4/* 452*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1e3/* 483*/:9'h1d9/* 473*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1ee/* 494*/:9'h1e4/* 484*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1f9/* 505*/:9'h1ef/* 495*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h204/* 516*/:9'h1fa/* 506*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h20f/* 527*/:10'h205/* 517*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h21a/* 538*/:10'h210/* 528*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h225/* 549*/:10'h21b/* 539*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h230/* 560*/:10'h226/* 550*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h23a/* 570*/:10'h231/* 561*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h244/* 580*/:10'h23b/* 571*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h24e/* 590*/:10'h245/* 581*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h258/* 600*/:10'h24f/* 591*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h262/* 610*/:10'h259/* 601*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h263/* 611*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_2(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_2 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_3(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[1:0] T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[1:0] T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[10:0] T230;
  wire[10:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire[2:0] T238;
  wire[2:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire[2:0] T246;
  wire[2:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  wire[1:0] T260;
  wire[1:0] T261;
  wire[2:0] T262;
  wire[2:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[1:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire[2:0] T278;
  wire[2:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[1:0] T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire[2:0] T286;
  wire[2:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[1:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[2:0] T302;
  wire[2:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[10:0] T310;
  wire[10:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[1:0] T315;
  wire[1:0] T316;
  wire[1:0] T317;
  wire[2:0] T318;
  wire[2:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[2:0] T326;
  wire[2:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[1:0] T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[1:0] T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[10:0] T350;
  wire[10:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[10:0] T390;
  wire[10:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[1:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire[2:0] T398;
  wire[2:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[1:0] T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire[2:0] T406;
  wire[2:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[1:0] T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire[2:0] T414;
  wire[2:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[1:0] T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire[2:0] T422;
  wire[2:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[10:0] T430;
  wire[10:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire[2:0] T438;
  wire[2:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire[2:0] T446;
  wire[2:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire[1:0] T462;
  wire[1:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[3:0] T467;
  wire[3:0] T468;
  wire[3:0] T469;
  wire[10:0] T470;
  wire[10:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire[1:0] T478;
  wire[1:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire[1:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire[1:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[10:0] T510;
  wire[10:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire[3:0] T547;
  wire[3:0] T548;
  wire[3:0] T549;
  wire[10:0] T550;
  wire[10:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire[1:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire[1:0] T582;
  wire[1:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[3:0] T587;
  wire[3:0] T588;
  wire[3:0] T589;
  wire[9:0] T590;
  wire[9:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire[1:0] T598;
  wire[1:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire[1:0] T606;
  wire[1:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[1:0] T614;
  wire[1:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[1:0] T622;
  wire[1:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[3:0] T627;
  wire[3:0] T628;
  wire[3:0] T629;
  wire[9:0] T630;
  wire[9:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire[1:0] T638;
  wire[1:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire[1:0] T646;
  wire[1:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire[1:0] T654;
  wire[1:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire[1:0] T662;
  wire[1:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[3:0] T667;
  wire[3:0] T668;
  wire[3:0] T669;
  wire[9:0] T670;
  wire[9:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[1:0] T678;
  wire[1:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire[1:0] T686;
  wire[1:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire[3:0] T707;
  wire[3:0] T708;
  wire[3:0] T709;
  wire[9:0] T710;
  wire[9:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire[3:0] T747;
  wire[3:0] T748;
  wire[3:0] T749;
  wire[9:0] T750;
  wire[9:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire[3:0] T787;
  wire[3:0] T788;
  wire[3:0] T789;
  wire[9:0] T790;
  wire[9:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[10:0] T814;
  wire[10:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[10:0] T822;
  wire[10:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[10:0] T830;
  wire[10:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[10:0] T838;
  wire[10:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[10:0] T846;
  wire[10:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[3:0] T851;
  wire[3:0] T852;
  wire[3:0] T853;
  wire[10:0] T854;
  wire[10:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[10:0] T862;
  wire[10:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[10:0] T870;
  wire[10:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[10:0] T878;
  wire[10:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[9:0] T886;
  wire[9:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[9:0] T894;
  wire[9:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[9:0] T902;
  wire[9:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[9:0] T910;
  wire[9:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[9:0] T918;
  wire[9:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[3:0] T932;
  wire[3:0] T933;
  wire[10:0] T934;
  wire[10:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[10:0] T942;
  wire[10:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[10:0] T950;
  wire[10:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[10:0] T958;
  wire[10:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[10:0] T966;
  wire[10:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[10:0] T974;
  wire[10:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[10:0] T982;
  wire[10:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[10:0] T990;
  wire[10:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[10:0] T998;
  wire[10:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire[3:0] T1011;
  wire[3:0] T1012;
  wire[3:0] T1013;
  wire[9:0] T1014;
  wire[9:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[9:0] T1030;
  wire[9:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[9:0] T1046;
  wire[9:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[5'h10/* 16*/:3'h6/* 6*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[5'h13/* 19*/:5'h11/* 17*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[6'h27/* 39*/:5'h1d/* 29*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[5'h15/* 21*/:5'h14/* 20*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[6'h2a/* 42*/:6'h28/* 40*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[6'h3e/* 62*/:6'h34/* 52*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[7'h41/* 65*/:6'h3f/* 63*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[7'h55/* 85*/:7'h4b/* 75*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[7'h58/* 88*/:7'h56/* 86*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[7'h6c/* 108*/:7'h62/* 98*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[6'h39/* 57*/:6'h38/* 56*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[8'h83/* 131*/:7'h79/* 121*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[8'h86/* 134*/:8'h84/* 132*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h4d/* 77*/:7'h4a/* 74*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[8'h98/* 152*/:8'h8e/* 142*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h4e/* 78*/:7'h4e/* 78*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[8'h9a/* 154*/:8'h99/* 153*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[8'ha0/* 160*/:8'h9f/* 159*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[7'h55/* 85*/:7'h52/* 82*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[8'hab/* 171*/:8'ha1/* 161*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[8'had/* 173*/:8'hac/* 172*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[8'hbe/* 190*/:8'hb4/* 180*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[8'hc0/* 192*/:8'hbf/* 191*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[8'hc6/* 198*/:8'hc5/* 197*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[7'h65/* 101*/:7'h62/* 98*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[8'hd0/* 208*/:8'hc7/* 199*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[7'h66/* 102*/:7'h66/* 102*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[8'hd2/* 210*/:8'hd1/* 209*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[8'hd6/* 214*/:8'hd5/* 213*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[8'hd8/* 216*/:8'hd7/* 215*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[7'h6d/* 109*/:7'h6a/* 106*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[8'he2/* 226*/:8'hd9/* 217*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[7'h6e/* 110*/:7'h6e/* 110*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[8'he4/* 228*/:8'he3/* 227*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[8'hf4/* 244*/:8'heb/* 235*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[8'hf6/* 246*/:8'hf5/* 245*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[7'h7d/* 125*/:7'h7a/* 122*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h106/* 262*/:8'hfd/* 253*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h108/* 264*/:9'h107/* 263*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h118/* 280*/:9'h10f/* 271*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h11a/* 282*/:9'h119/* 281*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h12a/* 298*/:9'h121/* 289*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h12c/* 300*/:9'h12b/* 299*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h144/* 324*/:9'h13a/* 314*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h14f/* 335*/:9'h145/* 325*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h15a/* 346*/:9'h150/* 336*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h165/* 357*/:9'h15b/* 347*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h170/* 368*/:9'h166/* 358*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h17b/* 379*/:9'h171/* 369*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h186/* 390*/:9'h17c/* 380*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h191/* 401*/:9'h187/* 391*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h19b/* 411*/:9'h192/* 402*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h1a5/* 421*/:9'h19c/* 412*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h1af/* 431*/:9'h1a6/* 422*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1b9/* 441*/:9'h1b0/* 432*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1c3/* 451*/:9'h1ba/* 442*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1cd/* 461*/:9'h1c4/* 452*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1e3/* 483*/:9'h1d9/* 473*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1ee/* 494*/:9'h1e4/* 484*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1f9/* 505*/:9'h1ef/* 495*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h204/* 516*/:9'h1fa/* 506*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h20f/* 527*/:10'h205/* 517*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h21a/* 538*/:10'h210/* 528*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h225/* 549*/:10'h21b/* 539*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h230/* 560*/:10'h226/* 550*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h23a/* 570*/:10'h231/* 561*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h244/* 580*/:10'h23b/* 571*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h24e/* 590*/:10'h245/* 581*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h258/* 600*/:10'h24f/* 591*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h262/* 610*/:10'h259/* 601*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h263/* 611*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_3(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_3 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_4(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[1:0] T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[1:0] T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[1:0] T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire[2:0] T230;
  wire[2:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[10:0] T238;
  wire[10:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire[2:0] T246;
  wire[2:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[1:0] T259;
  wire[1:0] T260;
  wire[1:0] T261;
  wire[2:0] T262;
  wire[2:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[1:0] T267;
  wire[1:0] T268;
  wire[1:0] T269;
  wire[2:0] T270;
  wire[2:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[1:0] T283;
  wire[1:0] T284;
  wire[1:0] T285;
  wire[2:0] T286;
  wire[2:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire[1:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[1:0] T299;
  wire[1:0] T300;
  wire[1:0] T301;
  wire[2:0] T302;
  wire[2:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[1:0] T307;
  wire[1:0] T308;
  wire[1:0] T309;
  wire[2:0] T310;
  wire[2:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[10:0] T318;
  wire[10:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[1:0] T323;
  wire[1:0] T324;
  wire[1:0] T325;
  wire[2:0] T326;
  wire[2:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[1:0] T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[1:0] T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[1:0] T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire[2:0] T350;
  wire[2:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[10:0] T358;
  wire[10:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[1:0] T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire[2:0] T382;
  wire[2:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[1:0] T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire[2:0] T390;
  wire[2:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[10:0] T398;
  wire[10:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[1:0] T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire[2:0] T406;
  wire[2:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[1:0] T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire[2:0] T414;
  wire[2:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[1:0] T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire[2:0] T422;
  wire[2:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[1:0] T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire[2:0] T430;
  wire[2:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[10:0] T438;
  wire[10:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[1:0] T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire[2:0] T446;
  wire[2:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire[1:0] T462;
  wire[1:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire[1:0] T470;
  wire[1:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[3:0] T475;
  wire[3:0] T476;
  wire[3:0] T477;
  wire[10:0] T478;
  wire[10:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire[1:0] T486;
  wire[1:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire[1:0] T494;
  wire[1:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire[3:0] T515;
  wire[3:0] T516;
  wire[3:0] T517;
  wire[10:0] T518;
  wire[10:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire[3:0] T555;
  wire[3:0] T556;
  wire[3:0] T557;
  wire[10:0] T558;
  wire[10:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire[1:0] T574;
  wire[1:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire[1:0] T582;
  wire[1:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire[1:0] T590;
  wire[1:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[3:0] T595;
  wire[3:0] T596;
  wire[3:0] T597;
  wire[9:0] T598;
  wire[9:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire[1:0] T606;
  wire[1:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire[1:0] T614;
  wire[1:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[1:0] T622;
  wire[1:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[3:0] T635;
  wire[3:0] T636;
  wire[3:0] T637;
  wire[9:0] T638;
  wire[9:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire[1:0] T646;
  wire[1:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire[1:0] T654;
  wire[1:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire[1:0] T662;
  wire[1:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire[3:0] T675;
  wire[3:0] T676;
  wire[3:0] T677;
  wire[9:0] T678;
  wire[9:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire[1:0] T686;
  wire[1:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire[3:0] T715;
  wire[3:0] T716;
  wire[3:0] T717;
  wire[9:0] T718;
  wire[9:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire[3:0] T755;
  wire[3:0] T756;
  wire[3:0] T757;
  wire[9:0] T758;
  wire[9:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire[3:0] T795;
  wire[3:0] T796;
  wire[3:0] T797;
  wire[9:0] T798;
  wire[9:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[10:0] T814;
  wire[10:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[10:0] T822;
  wire[10:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[10:0] T830;
  wire[10:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[10:0] T838;
  wire[10:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[10:0] T846;
  wire[10:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[3:0] T851;
  wire[3:0] T852;
  wire[3:0] T853;
  wire[10:0] T854;
  wire[10:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[10:0] T862;
  wire[10:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[10:0] T870;
  wire[10:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[10:0] T878;
  wire[10:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[9:0] T886;
  wire[9:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[9:0] T894;
  wire[9:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[9:0] T902;
  wire[9:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[9:0] T910;
  wire[9:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[9:0] T918;
  wire[9:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[3:0] T932;
  wire[3:0] T933;
  wire[10:0] T934;
  wire[10:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[10:0] T942;
  wire[10:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[10:0] T950;
  wire[10:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[10:0] T958;
  wire[10:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[10:0] T966;
  wire[10:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[10:0] T974;
  wire[10:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[10:0] T982;
  wire[10:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[10:0] T990;
  wire[10:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[10:0] T998;
  wire[10:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire[3:0] T1011;
  wire[3:0] T1012;
  wire[3:0] T1013;
  wire[9:0] T1014;
  wire[9:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[9:0] T1030;
  wire[9:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[9:0] T1046;
  wire[9:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'h9/* 9*/:3'h6/* 6*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[5'h13/* 19*/:4'h9/* 9*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[5'h1f/* 31*/:5'h1d/* 29*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[5'h15/* 21*/:5'h12/* 18*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[6'h2a/* 42*/:6'h20/* 32*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[6'h36/* 54*/:6'h34/* 52*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h21/* 33*/:5'h1e/* 30*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[6'h2d/* 45*/:6'h2a/* 42*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[7'h58/* 88*/:7'h4e/* 78*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[7'h64/* 100*/:7'h62/* 98*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[6'h39/* 57*/:6'h36/* 54*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[7'h6f/* 111*/:7'h65/* 101*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[8'h86/* 134*/:7'h7c/* 124*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[8'h9a/* 154*/:8'h90/* 144*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[8'ha0/* 160*/:8'h9f/* 159*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[8'ha2/* 162*/:8'ha1/* 161*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[7'h56/* 86*/:7'h53/* 83*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[8'had/* 173*/:8'ha3/* 163*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[7'h5a/* 90*/:7'h5a/* 90*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[7'h5e/* 94*/:7'h5b/* 91*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[8'hc0/* 192*/:8'hb6/* 182*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[8'hc6/* 198*/:8'hc5/* 197*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[7'h62/* 98*/:7'h62/* 98*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[7'h66/* 102*/:7'h63/* 99*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[8'hd2/* 210*/:8'hc9/* 201*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[8'hd6/* 214*/:8'hd5/* 213*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[8'hd8/* 216*/:8'hd7/* 215*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[7'h6a/* 106*/:7'h6a/* 106*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[7'h6e/* 110*/:7'h6b/* 107*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[8'he4/* 228*/:8'hdb/* 219*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[8'hea/* 234*/:8'he9/* 233*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[8'hec/* 236*/:8'heb/* 235*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[8'hf6/* 246*/:8'hed/* 237*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[7'h7e/* 126*/:7'h7b/* 123*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h108/* 264*/:8'hff/* 255*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h110/* 272*/:9'h10f/* 271*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'h86/* 134*/:8'h83/* 131*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h11a/* 282*/:9'h111/* 273*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h12c/* 300*/:9'h123/* 291*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h144/* 324*/:9'h13a/* 314*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h14f/* 335*/:9'h145/* 325*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h15a/* 346*/:9'h150/* 336*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h165/* 357*/:9'h15b/* 347*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h170/* 368*/:9'h166/* 358*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h17b/* 379*/:9'h171/* 369*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h186/* 390*/:9'h17c/* 380*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h191/* 401*/:9'h187/* 391*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h19b/* 411*/:9'h192/* 402*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h1a5/* 421*/:9'h19c/* 412*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h1af/* 431*/:9'h1a6/* 422*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1b9/* 441*/:9'h1b0/* 432*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1c3/* 451*/:9'h1ba/* 442*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1cd/* 461*/:9'h1c4/* 452*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1e3/* 483*/:9'h1d9/* 473*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1ee/* 494*/:9'h1e4/* 484*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1f9/* 505*/:9'h1ef/* 495*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h204/* 516*/:9'h1fa/* 506*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h20f/* 527*/:10'h205/* 517*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h21a/* 538*/:10'h210/* 528*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h225/* 549*/:10'h21b/* 539*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h230/* 560*/:10'h226/* 550*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h23a/* 570*/:10'h231/* 561*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h244/* 580*/:10'h23b/* 571*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h24e/* 590*/:10'h245/* 581*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h258/* 600*/:10'h24f/* 591*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h262/* 610*/:10'h259/* 601*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h263/* 611*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_4(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_5(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_6(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_2 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_7(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_3 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_8(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_5(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [557:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[149:0] io_chanxy_out);

  wire[149:0] T0;
  wire[149:0] T1;
  wire[148:0] T2;
  wire[148:0] T3;
  wire[147:0] T4;
  wire[147:0] T5;
  wire[146:0] T6;
  wire[146:0] T7;
  wire[145:0] T8;
  wire[145:0] T9;
  wire[144:0] T10;
  wire[144:0] T11;
  wire[143:0] T12;
  wire[143:0] T13;
  wire[142:0] T14;
  wire[142:0] T15;
  wire[141:0] T16;
  wire[141:0] T17;
  wire[140:0] T18;
  wire[140:0] T19;
  wire[139:0] T20;
  wire[139:0] T21;
  wire[138:0] T22;
  wire[138:0] T23;
  wire[137:0] T24;
  wire[137:0] T25;
  wire[136:0] T26;
  wire[136:0] T27;
  wire[135:0] T28;
  wire[135:0] T29;
  wire[134:0] T30;
  wire[134:0] T31;
  wire[133:0] T32;
  wire[133:0] T33;
  wire[132:0] T34;
  wire[132:0] T35;
  wire[131:0] T36;
  wire[131:0] T37;
  wire[130:0] T38;
  wire[130:0] T39;
  wire[129:0] T40;
  wire[129:0] T41;
  wire[128:0] T42;
  wire[128:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[126:0] T46;
  wire[126:0] T47;
  wire[125:0] T48;
  wire[125:0] T49;
  wire[124:0] T50;
  wire[124:0] T51;
  wire[123:0] T52;
  wire[123:0] T53;
  wire[122:0] T54;
  wire[122:0] T55;
  wire[121:0] T56;
  wire[121:0] T57;
  wire[120:0] T58;
  wire[120:0] T59;
  wire[119:0] T60;
  wire[119:0] T61;
  wire[118:0] T62;
  wire[118:0] T63;
  wire[117:0] T64;
  wire[117:0] T65;
  wire[116:0] T66;
  wire[116:0] T67;
  wire[115:0] T68;
  wire[115:0] T69;
  wire[114:0] T70;
  wire[114:0] T71;
  wire[113:0] T72;
  wire[113:0] T73;
  wire[112:0] T74;
  wire[112:0] T75;
  wire[111:0] T76;
  wire[111:0] T77;
  wire[110:0] T78;
  wire[110:0] T79;
  wire[109:0] T80;
  wire[109:0] T81;
  wire[108:0] T82;
  wire[108:0] T83;
  wire[107:0] T84;
  wire[107:0] T85;
  wire[106:0] T86;
  wire[106:0] T87;
  wire[105:0] T88;
  wire[105:0] T89;
  wire[104:0] T90;
  wire[104:0] T91;
  wire[103:0] T92;
  wire[103:0] T93;
  wire[102:0] T94;
  wire[102:0] T95;
  wire[101:0] T96;
  wire[101:0] T97;
  wire[100:0] T98;
  wire[100:0] T99;
  wire[99:0] T100;
  wire[99:0] T101;
  wire[98:0] T102;
  wire[98:0] T103;
  wire[97:0] T104;
  wire[97:0] T105;
  wire[96:0] T106;
  wire[96:0] T107;
  wire[95:0] T108;
  wire[95:0] T109;
  wire[94:0] T110;
  wire[94:0] T111;
  wire[93:0] T112;
  wire[93:0] T113;
  wire[92:0] T114;
  wire[92:0] T115;
  wire[91:0] T116;
  wire[91:0] T117;
  wire[90:0] T118;
  wire[90:0] T119;
  wire[89:0] T120;
  wire[89:0] T121;
  wire[88:0] T122;
  wire[88:0] T123;
  wire[87:0] T124;
  wire[87:0] T125;
  wire[86:0] T126;
  wire[86:0] T127;
  wire[85:0] T128;
  wire[85:0] T129;
  wire[84:0] T130;
  wire[84:0] T131;
  wire[83:0] T132;
  wire[83:0] T133;
  wire[82:0] T134;
  wire[82:0] T135;
  wire[81:0] T136;
  wire[81:0] T137;
  wire[80:0] T138;
  wire[80:0] T139;
  wire[79:0] T140;
  wire[79:0] T141;
  wire[78:0] T142;
  wire[78:0] T143;
  wire[77:0] T144;
  wire[77:0] T145;
  wire[76:0] T146;
  wire[76:0] T147;
  wire[75:0] T148;
  wire[75:0] T149;
  wire[74:0] T150;
  wire[74:0] T151;
  wire[73:0] T152;
  wire[73:0] T153;
  wire[72:0] T154;
  wire[72:0] T155;
  wire[71:0] T156;
  wire[71:0] T157;
  wire[70:0] T158;
  wire[70:0] T159;
  wire[69:0] T160;
  wire[69:0] T161;
  wire[68:0] T162;
  wire[68:0] T163;
  wire[67:0] T164;
  wire[67:0] T165;
  wire[66:0] T166;
  wire[66:0] T167;
  wire[65:0] T168;
  wire[65:0] T169;
  wire[64:0] T170;
  wire[64:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[62:0] T174;
  wire[62:0] T175;
  wire[61:0] T176;
  wire[61:0] T177;
  wire[60:0] T178;
  wire[60:0] T179;
  wire[59:0] T180;
  wire[59:0] T181;
  wire[58:0] T182;
  wire[58:0] T183;
  wire[57:0] T184;
  wire[57:0] T185;
  wire[56:0] T186;
  wire[56:0] T187;
  wire[55:0] T188;
  wire[55:0] T189;
  wire[54:0] T190;
  wire[54:0] T191;
  wire[53:0] T192;
  wire[53:0] T193;
  wire[52:0] T194;
  wire[52:0] T195;
  wire[51:0] T196;
  wire[51:0] T197;
  wire[50:0] T198;
  wire[50:0] T199;
  wire[49:0] T200;
  wire[49:0] T201;
  wire[48:0] T202;
  wire[48:0] T203;
  wire[47:0] T204;
  wire[47:0] T205;
  wire[46:0] T206;
  wire[46:0] T207;
  wire[45:0] T208;
  wire[45:0] T209;
  wire[44:0] T210;
  wire[44:0] T211;
  wire[43:0] T212;
  wire[43:0] T213;
  wire[42:0] T214;
  wire[42:0] T215;
  wire[41:0] T216;
  wire[41:0] T217;
  wire[40:0] T218;
  wire[40:0] T219;
  wire[39:0] T220;
  wire[39:0] T221;
  wire[38:0] T222;
  wire[38:0] T223;
  wire[37:0] T224;
  wire[37:0] T225;
  wire[36:0] T226;
  wire[36:0] T227;
  wire[35:0] T228;
  wire[35:0] T229;
  wire[34:0] T230;
  wire[34:0] T231;
  wire[33:0] T232;
  wire[33:0] T233;
  wire[32:0] T234;
  wire[32:0] T235;
  wire[31:0] T236;
  wire[31:0] T237;
  wire[30:0] T238;
  wire[30:0] T239;
  wire[29:0] T240;
  wire[29:0] T241;
  wire[28:0] T242;
  wire[28:0] T243;
  wire[27:0] T244;
  wire[27:0] T245;
  wire[26:0] T246;
  wire[26:0] T247;
  wire[25:0] T248;
  wire[25:0] T249;
  wire[24:0] T250;
  wire[24:0] T251;
  wire[23:0] T252;
  wire[23:0] T253;
  wire[22:0] T254;
  wire[22:0] T255;
  wire[21:0] T256;
  wire[21:0] T257;
  wire[20:0] T258;
  wire[20:0] T259;
  wire[19:0] T260;
  wire[19:0] T261;
  wire[18:0] T262;
  wire[18:0] T263;
  wire[17:0] T264;
  wire[17:0] T265;
  wire[16:0] T266;
  wire[16:0] T267;
  wire[15:0] T268;
  wire[15:0] T269;
  wire[14:0] T270;
  wire[14:0] T271;
  wire[13:0] T272;
  wire[13:0] T273;
  wire[12:0] T274;
  wire[12:0] T275;
  wire[11:0] T276;
  wire[11:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire[9:0] T280;
  wire[9:0] T281;
  wire[8:0] T282;
  wire[8:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[6:0] T286;
  wire[6:0] T287;
  wire[5:0] T288;
  wire[5:0] T289;
  wire[4:0] T290;
  wire[4:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire[1:0] T296;
  wire[1:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[1:0] T304;
  wire[1:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire[1:0] T312;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire[1:0] T328;
  wire[1:0] T329;
  wire T330;
  wire T331;
  wire T332;
  wire[3:0] T333;
  wire[3:0] T334;
  wire[3:0] T335;
  wire[8:0] T336;
  wire[8:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[1:0] T344;
  wire[1:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire[1:0] T352;
  wire[1:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire[1:0] T360;
  wire[1:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[1:0] T368;
  wire[1:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire[3:0] T373;
  wire[3:0] T374;
  wire[3:0] T375;
  wire[8:0] T376;
  wire[8:0] T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire[1:0] T384;
  wire[1:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire[1:0] T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire[1:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[1:0] T408;
  wire[1:0] T409;
  wire T410;
  wire T411;
  wire T412;
  wire[3:0] T413;
  wire[3:0] T414;
  wire[3:0] T415;
  wire[8:0] T416;
  wire[8:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[1:0] T424;
  wire[1:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire[1:0] T432;
  wire[1:0] T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire[1:0] T448;
  wire[1:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire[3:0] T453;
  wire[3:0] T454;
  wire[3:0] T455;
  wire[8:0] T456;
  wire[8:0] T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire[1:0] T464;
  wire[1:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire[1:0] T480;
  wire[1:0] T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[1:0] T488;
  wire[1:0] T489;
  wire T490;
  wire T491;
  wire T492;
  wire[3:0] T493;
  wire[3:0] T494;
  wire[3:0] T495;
  wire[8:0] T496;
  wire[8:0] T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire[1:0] T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire[1:0] T512;
  wire[1:0] T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire[1:0] T520;
  wire[1:0] T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire[1:0] T528;
  wire[1:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire[3:0] T533;
  wire[3:0] T534;
  wire[3:0] T535;
  wire[8:0] T536;
  wire[8:0] T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire[1:0] T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[1:0] T552;
  wire[1:0] T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire[1:0] T560;
  wire[1:0] T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire[1:0] T568;
  wire[1:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire[3:0] T573;
  wire[3:0] T574;
  wire[3:0] T575;
  wire[8:0] T576;
  wire[8:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire[1:0] T584;
  wire[1:0] T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[1:0] T592;
  wire[1:0] T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire[1:0] T600;
  wire[1:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire[1:0] T608;
  wire[1:0] T609;
  wire T610;
  wire T611;
  wire T612;
  wire[3:0] T613;
  wire[3:0] T614;
  wire[3:0] T615;
  wire[8:0] T616;
  wire[8:0] T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[1:0] T624;
  wire[1:0] T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[1:0] T632;
  wire[1:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire[1:0] T640;
  wire[1:0] T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire[1:0] T648;
  wire[1:0] T649;
  wire T650;
  wire T651;
  wire T652;
  wire[3:0] T653;
  wire[3:0] T654;
  wire[3:0] T655;
  wire[8:0] T656;
  wire[8:0] T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire[1:0] T664;
  wire[1:0] T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire[1:0] T672;
  wire[1:0] T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire[1:0] T680;
  wire[1:0] T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire[1:0] T688;
  wire[1:0] T689;
  wire T690;
  wire T691;
  wire T692;
  wire[3:0] T693;
  wire[3:0] T694;
  wire[3:0] T695;
  wire[8:0] T696;
  wire[8:0] T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire[1:0] T704;
  wire[1:0] T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire[1:0] T712;
  wire[1:0] T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[1:0] T720;
  wire[1:0] T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire T726;
  wire T727;
  wire[1:0] T728;
  wire[1:0] T729;
  wire T730;
  wire T731;
  wire T732;
  wire[3:0] T733;
  wire[3:0] T734;
  wire[3:0] T735;
  wire[8:0] T736;
  wire[8:0] T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire[1:0] T744;
  wire[1:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire[1:0] T752;
  wire[1:0] T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire[1:0] T760;
  wire[1:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire[1:0] T768;
  wire[1:0] T769;
  wire T770;
  wire T771;
  wire T772;
  wire[3:0] T773;
  wire[3:0] T774;
  wire[3:0] T775;
  wire[8:0] T776;
  wire[8:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[1:0] T784;
  wire[1:0] T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire[1:0] T792;
  wire[1:0] T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire[1:0] T800;
  wire[1:0] T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire[1:0] T808;
  wire[1:0] T809;
  wire T810;
  wire T811;
  wire T812;
  wire[3:0] T813;
  wire[3:0] T814;
  wire[3:0] T815;
  wire[8:0] T816;
  wire[8:0] T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire T822;
  wire T823;
  wire[1:0] T824;
  wire[1:0] T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire[1:0] T832;
  wire[1:0] T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire T838;
  wire T839;
  wire[1:0] T840;
  wire[1:0] T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire T847;
  wire[1:0] T848;
  wire[1:0] T849;
  wire T850;
  wire T851;
  wire T852;
  wire[3:0] T853;
  wire[3:0] T854;
  wire[3:0] T855;
  wire[8:0] T856;
  wire[8:0] T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire[1:0] T864;
  wire[1:0] T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire[1:0] T872;
  wire[1:0] T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire[1:0] T880;
  wire[1:0] T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire[1:0] T888;
  wire[1:0] T889;
  wire T890;
  wire T891;
  wire T892;
  wire[3:0] T893;
  wire[3:0] T894;
  wire[3:0] T895;
  wire[8:0] T896;
  wire[8:0] T897;
  wire T898;
  wire T899;
  wire T900;
  wire[1:0] T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire[2:0] T904;
  wire[2:0] T905;
  wire T906;
  wire T907;
  wire T908;
  wire[1:0] T909;
  wire[1:0] T910;
  wire[1:0] T911;
  wire[2:0] T912;
  wire[2:0] T913;
  wire T914;
  wire T915;
  wire T916;
  wire[1:0] T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire[2:0] T920;
  wire[2:0] T921;
  wire T922;
  wire T923;
  wire T924;
  wire[1:0] T925;
  wire[1:0] T926;
  wire[1:0] T927;
  wire[2:0] T928;
  wire[2:0] T929;
  wire T930;
  wire T931;
  wire T932;
  wire[1:0] T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire[2:0] T936;
  wire[2:0] T937;
  wire T938;
  wire T939;
  wire T940;
  wire[1:0] T941;
  wire[1:0] T942;
  wire[1:0] T943;
  wire[2:0] T944;
  wire[2:0] T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire[1:0] T952;
  wire[1:0] T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire[1:0] T960;
  wire[1:0] T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire T966;
  wire T967;
  wire[1:0] T968;
  wire[1:0] T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire[1:0] T976;
  wire[1:0] T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire[1:0] T984;
  wire[1:0] T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire[1:0] T992;
  wire[1:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[1:0] T1000;
  wire[1:0] T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire T1006;
  wire T1007;
  wire[1:0] T1008;
  wire[1:0] T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire T1015;
  wire[1:0] T1016;
  wire[1:0] T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire[1:0] T1021;
  wire[1:0] T1022;
  wire[1:0] T1023;
  wire[2:0] T1024;
  wire[2:0] T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire[1:0] T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire[2:0] T1032;
  wire[2:0] T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire[1:0] T1037;
  wire[1:0] T1038;
  wire[1:0] T1039;
  wire[2:0] T1040;
  wire[2:0] T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire[1:0] T1045;
  wire[1:0] T1046;
  wire[1:0] T1047;
  wire[2:0] T1048;
  wire[2:0] T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire[1:0] T1053;
  wire[1:0] T1054;
  wire[1:0] T1055;
  wire[2:0] T1056;
  wire[2:0] T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire[1:0] T1061;
  wire[1:0] T1062;
  wire[1:0] T1063;
  wire[2:0] T1064;
  wire[2:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire[1:0] T1072;
  wire[1:0] T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire T1078;
  wire T1079;
  wire[1:0] T1080;
  wire[1:0] T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire[1:0] T1088;
  wire[1:0] T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire[1:0] T1096;
  wire[1:0] T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire[1:0] T1104;
  wire[1:0] T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire[1:0] T1112;
  wire[1:0] T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire[1:0] T1120;
  wire[1:0] T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire T1127;
  wire[1:0] T1128;
  wire[1:0] T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire[1:0] T1136;
  wire[1:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire[1:0] T1141;
  wire[1:0] T1142;
  wire[1:0] T1143;
  wire[2:0] T1144;
  wire[2:0] T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire[1:0] T1149;
  wire[1:0] T1150;
  wire[1:0] T1151;
  wire[2:0] T1152;
  wire[2:0] T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire[1:0] T1157;
  wire[1:0] T1158;
  wire[1:0] T1159;
  wire[2:0] T1160;
  wire[2:0] T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire[1:0] T1165;
  wire[1:0] T1166;
  wire[1:0] T1167;
  wire[2:0] T1168;
  wire[2:0] T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire[1:0] T1173;
  wire[1:0] T1174;
  wire[1:0] T1175;
  wire[2:0] T1176;
  wire[2:0] T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire[1:0] T1181;
  wire[1:0] T1182;
  wire[1:0] T1183;
  wire[2:0] T1184;
  wire[2:0] T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire[1:0] T1192;
  wire[1:0] T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire[1:0] T1200;
  wire[1:0] T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[1:0] T1208;
  wire[1:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire[1:0] T1216;
  wire[1:0] T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire[1:0] T1224;
  wire[1:0] T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire[1:0] T1232;
  wire[1:0] T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire[1:0] T1240;
  wire[1:0] T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire[1:0] T1248;
  wire[1:0] T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire[1:0] T1256;
  wire[1:0] T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire[3:0] T1261;
  wire[3:0] T1262;
  wire[3:0] T1263;
  wire[10:0] T1264;
  wire[10:0] T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire[1:0] T1269;
  wire[1:0] T1270;
  wire[1:0] T1271;
  wire[2:0] T1272;
  wire[2:0] T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire[3:0] T1277;
  wire[3:0] T1278;
  wire[3:0] T1279;
  wire[10:0] T1280;
  wire[10:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire[1:0] T1285;
  wire[1:0] T1286;
  wire[1:0] T1287;
  wire[2:0] T1288;
  wire[2:0] T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire[3:0] T1293;
  wire[3:0] T1294;
  wire[3:0] T1295;
  wire[10:0] T1296;
  wire[10:0] T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire[1:0] T1301;
  wire[1:0] T1302;
  wire[1:0] T1303;
  wire[2:0] T1304;
  wire[2:0] T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire[3:0] T1309;
  wire[3:0] T1310;
  wire[3:0] T1311;
  wire[10:0] T1312;
  wire[10:0] T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire[1:0] T1317;
  wire[1:0] T1318;
  wire[1:0] T1319;
  wire[2:0] T1320;
  wire[2:0] T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire[3:0] T1325;
  wire[3:0] T1326;
  wire[3:0] T1327;
  wire[10:0] T1328;
  wire[10:0] T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire[1:0] T1333;
  wire[1:0] T1334;
  wire[1:0] T1335;
  wire[2:0] T1336;
  wire[2:0] T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire[3:0] T1341;
  wire[3:0] T1342;
  wire[3:0] T1343;
  wire[10:0] T1344;
  wire[10:0] T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire[1:0] T1349;
  wire[1:0] T1350;
  wire[1:0] T1351;
  wire[2:0] T1352;
  wire[2:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire[3:0] T1357;
  wire[3:0] T1358;
  wire[3:0] T1359;
  wire[10:0] T1360;
  wire[10:0] T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  wire T1366;
  wire T1367;
  wire[1:0] T1368;
  wire[1:0] T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire[3:0] T1373;
  wire[3:0] T1374;
  wire[3:0] T1375;
  wire[10:0] T1376;
  wire[10:0] T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire[1:0] T1384;
  wire[1:0] T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire[3:0] T1389;
  wire[3:0] T1390;
  wire[3:0] T1391;
  wire[10:0] T1392;
  wire[10:0] T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[1:0] T1400;
  wire[1:0] T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire[3:0] T1405;
  wire[3:0] T1406;
  wire[3:0] T1407;
  wire[9:0] T1408;
  wire[9:0] T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire T1414;
  wire T1415;
  wire[1:0] T1416;
  wire[1:0] T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire[3:0] T1421;
  wire[3:0] T1422;
  wire[3:0] T1423;
  wire[9:0] T1424;
  wire[9:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[1:0] T1432;
  wire[1:0] T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire[3:0] T1437;
  wire[3:0] T1438;
  wire[3:0] T1439;
  wire[9:0] T1440;
  wire[9:0] T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire[1:0] T1448;
  wire[1:0] T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire[3:0] T1453;
  wire[3:0] T1454;
  wire[3:0] T1455;
  wire[9:0] T1456;
  wire[9:0] T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire[1:0] T1464;
  wire[1:0] T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire[3:0] T1469;
  wire[3:0] T1470;
  wire[3:0] T1471;
  wire[9:0] T1472;
  wire[9:0] T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire T1478;
  wire T1479;
  wire[1:0] T1480;
  wire[1:0] T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire[3:0] T1485;
  wire[3:0] T1486;
  wire[3:0] T1487;
  wire[9:0] T1488;
  wire[9:0] T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[1:0] T1496;
  wire[1:0] T1497;
  wire[22:0] T1498;
  wire[22:0] T1499;
  wire[21:0] T1500;
  wire[21:0] T1501;
  wire[20:0] T1502;
  wire[20:0] T1503;
  wire[19:0] T1504;
  wire[19:0] T1505;
  wire[18:0] T1506;
  wire[18:0] T1507;
  wire[17:0] T1508;
  wire[17:0] T1509;
  wire[16:0] T1510;
  wire[16:0] T1511;
  wire[15:0] T1512;
  wire[15:0] T1513;
  wire[14:0] T1514;
  wire[14:0] T1515;
  wire[13:0] T1516;
  wire[13:0] T1517;
  wire[12:0] T1518;
  wire[12:0] T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[10:0] T1522;
  wire[10:0] T1523;
  wire[9:0] T1524;
  wire[9:0] T1525;
  wire[8:0] T1526;
  wire[8:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[6:0] T1530;
  wire[6:0] T1531;
  wire[5:0] T1532;
  wire[5:0] T1533;
  wire[4:0] T1534;
  wire[4:0] T1535;
  wire[3:0] T1536;
  wire[3:0] T1537;
  wire[2:0] T1538;
  wire[2:0] T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[11:0] T1660;
  wire[11:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[11:0] T1668;
  wire[11:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[11:0] T1676;
  wire[11:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[11:0] T1684;
  wire[11:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[11:0] T1692;
  wire[11:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[11:0] T1700;
  wire[11:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[11:0] T1708;
  wire[11:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[11:0] T1716;
  wire[11:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[11:0] T1724;
  wire[11:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1490, T2};
  assign T2 = T3;
  assign T3 = {T1482, T4};
  assign T4 = T5;
  assign T5 = {T1474, T6};
  assign T6 = T7;
  assign T7 = {T1466, T8};
  assign T8 = T9;
  assign T9 = {T1458, T10};
  assign T10 = T11;
  assign T11 = {T1450, T12};
  assign T12 = T13;
  assign T13 = {T1442, T14};
  assign T14 = T15;
  assign T15 = {T1434, T16};
  assign T16 = T17;
  assign T17 = {T1426, T18};
  assign T18 = T19;
  assign T19 = {T1418, T20};
  assign T20 = T21;
  assign T21 = {T1410, T22};
  assign T22 = T23;
  assign T23 = {T1402, T24};
  assign T24 = T25;
  assign T25 = {T1394, T26};
  assign T26 = T27;
  assign T27 = {T1386, T28};
  assign T28 = T29;
  assign T29 = {T1378, T30};
  assign T30 = T31;
  assign T31 = {T1370, T32};
  assign T32 = T33;
  assign T33 = {T1362, T34};
  assign T34 = T35;
  assign T35 = {T1354, T36};
  assign T36 = T37;
  assign T37 = {T1346, T38};
  assign T38 = T39;
  assign T39 = {T1338, T40};
  assign T40 = T41;
  assign T41 = {T1330, T42};
  assign T42 = T43;
  assign T43 = {T1322, T44};
  assign T44 = T45;
  assign T45 = {T1314, T46};
  assign T46 = T47;
  assign T47 = {T1306, T48};
  assign T48 = T49;
  assign T49 = {T1298, T50};
  assign T50 = T51;
  assign T51 = {T1290, T52};
  assign T52 = T53;
  assign T53 = {T1282, T54};
  assign T54 = T55;
  assign T55 = {T1274, T56};
  assign T56 = T57;
  assign T57 = {T1266, T58};
  assign T58 = T59;
  assign T59 = {T1258, T60};
  assign T60 = T61;
  assign T61 = {T1250, T62};
  assign T62 = T63;
  assign T63 = {T1242, T64};
  assign T64 = T65;
  assign T65 = {T1234, T66};
  assign T66 = T67;
  assign T67 = {T1226, T68};
  assign T68 = T69;
  assign T69 = {T1218, T70};
  assign T70 = T71;
  assign T71 = {T1210, T72};
  assign T72 = T73;
  assign T73 = {T1202, T74};
  assign T74 = T75;
  assign T75 = {T1194, T76};
  assign T76 = T77;
  assign T77 = {T1186, T78};
  assign T78 = T79;
  assign T79 = {T1178, T80};
  assign T80 = T81;
  assign T81 = {T1170, T82};
  assign T82 = T83;
  assign T83 = {T1162, T84};
  assign T84 = T85;
  assign T85 = {T1154, T86};
  assign T86 = T87;
  assign T87 = {T1146, T88};
  assign T88 = T89;
  assign T89 = {T1138, T90};
  assign T90 = T91;
  assign T91 = {T1130, T92};
  assign T92 = T93;
  assign T93 = {T1122, T94};
  assign T94 = T95;
  assign T95 = {T1114, T96};
  assign T96 = T97;
  assign T97 = {T1106, T98};
  assign T98 = T99;
  assign T99 = {T1098, T100};
  assign T100 = T101;
  assign T101 = {T1090, T102};
  assign T102 = T103;
  assign T103 = {T1082, T104};
  assign T104 = T105;
  assign T105 = {T1074, T106};
  assign T106 = T107;
  assign T107 = {T1066, T108};
  assign T108 = T109;
  assign T109 = {T1058, T110};
  assign T110 = T111;
  assign T111 = {T1050, T112};
  assign T112 = T113;
  assign T113 = {T1042, T114};
  assign T114 = T115;
  assign T115 = {T1034, T116};
  assign T116 = T117;
  assign T117 = {T1026, T118};
  assign T118 = T119;
  assign T119 = {T1018, T120};
  assign T120 = T121;
  assign T121 = {T1010, T122};
  assign T122 = T123;
  assign T123 = {T1002, T124};
  assign T124 = T125;
  assign T125 = {T994, T126};
  assign T126 = T127;
  assign T127 = {T986, T128};
  assign T128 = T129;
  assign T129 = {T978, T130};
  assign T130 = T131;
  assign T131 = {T970, T132};
  assign T132 = T133;
  assign T133 = {T962, T134};
  assign T134 = T135;
  assign T135 = {T954, T136};
  assign T136 = T137;
  assign T137 = {T946, T138};
  assign T138 = T139;
  assign T139 = {T938, T140};
  assign T140 = T141;
  assign T141 = {T930, T142};
  assign T142 = T143;
  assign T143 = {T922, T144};
  assign T144 = T145;
  assign T145 = {T914, T146};
  assign T146 = T147;
  assign T147 = {T906, T148};
  assign T148 = T149;
  assign T149 = {T898, T150};
  assign T150 = T151;
  assign T151 = {T890, T152};
  assign T152 = T153;
  assign T153 = {T882, T154};
  assign T154 = T155;
  assign T155 = {T874, T156};
  assign T156 = T157;
  assign T157 = {T866, T158};
  assign T158 = T159;
  assign T159 = {T858, T160};
  assign T160 = T161;
  assign T161 = {T850, T162};
  assign T162 = T163;
  assign T163 = {T842, T164};
  assign T164 = T165;
  assign T165 = {T834, T166};
  assign T166 = T167;
  assign T167 = {T826, T168};
  assign T168 = T169;
  assign T169 = {T818, T170};
  assign T170 = T171;
  assign T171 = {T810, T172};
  assign T172 = T173;
  assign T173 = {T802, T174};
  assign T174 = T175;
  assign T175 = {T794, T176};
  assign T176 = T177;
  assign T177 = {T786, T178};
  assign T178 = T179;
  assign T179 = {T778, T180};
  assign T180 = T181;
  assign T181 = {T770, T182};
  assign T182 = T183;
  assign T183 = {T762, T184};
  assign T184 = T185;
  assign T185 = {T754, T186};
  assign T186 = T187;
  assign T187 = {T746, T188};
  assign T188 = T189;
  assign T189 = {T738, T190};
  assign T190 = T191;
  assign T191 = {T730, T192};
  assign T192 = T193;
  assign T193 = {T722, T194};
  assign T194 = T195;
  assign T195 = {T714, T196};
  assign T196 = T197;
  assign T197 = {T706, T198};
  assign T198 = T199;
  assign T199 = {T698, T200};
  assign T200 = T201;
  assign T201 = {T690, T202};
  assign T202 = T203;
  assign T203 = {T682, T204};
  assign T204 = T205;
  assign T205 = {T674, T206};
  assign T206 = T207;
  assign T207 = {T666, T208};
  assign T208 = T209;
  assign T209 = {T658, T210};
  assign T210 = T211;
  assign T211 = {T650, T212};
  assign T212 = T213;
  assign T213 = {T642, T214};
  assign T214 = T215;
  assign T215 = {T634, T216};
  assign T216 = T217;
  assign T217 = {T626, T218};
  assign T218 = T219;
  assign T219 = {T618, T220};
  assign T220 = T221;
  assign T221 = {T610, T222};
  assign T222 = T223;
  assign T223 = {T602, T224};
  assign T224 = T225;
  assign T225 = {T594, T226};
  assign T226 = T227;
  assign T227 = {T586, T228};
  assign T228 = T229;
  assign T229 = {T578, T230};
  assign T230 = T231;
  assign T231 = {T570, T232};
  assign T232 = T233;
  assign T233 = {T562, T234};
  assign T234 = T235;
  assign T235 = {T554, T236};
  assign T236 = T237;
  assign T237 = {T546, T238};
  assign T238 = T239;
  assign T239 = {T538, T240};
  assign T240 = T241;
  assign T241 = {T530, T242};
  assign T242 = T243;
  assign T243 = {T522, T244};
  assign T244 = T245;
  assign T245 = {T514, T246};
  assign T246 = T247;
  assign T247 = {T506, T248};
  assign T248 = T249;
  assign T249 = {T498, T250};
  assign T250 = T251;
  assign T251 = {T490, T252};
  assign T252 = T253;
  assign T253 = {T482, T254};
  assign T254 = T255;
  assign T255 = {T474, T256};
  assign T256 = T257;
  assign T257 = {T466, T258};
  assign T258 = T259;
  assign T259 = {T458, T260};
  assign T260 = T261;
  assign T261 = {T450, T262};
  assign T262 = T263;
  assign T263 = {T442, T264};
  assign T264 = T265;
  assign T265 = {T434, T266};
  assign T266 = T267;
  assign T267 = {T426, T268};
  assign T268 = T269;
  assign T269 = {T418, T270};
  assign T270 = T271;
  assign T271 = {T410, T272};
  assign T272 = T273;
  assign T273 = {T402, T274};
  assign T274 = T275;
  assign T275 = {T394, T276};
  assign T276 = T277;
  assign T277 = {T386, T278};
  assign T278 = T279;
  assign T279 = {T378, T280};
  assign T280 = T281;
  assign T281 = {T370, T282};
  assign T282 = T283;
  assign T283 = {T362, T284};
  assign T284 = T285;
  assign T285 = {T354, T286};
  assign T286 = T287;
  assign T287 = {T346, T288};
  assign T288 = T289;
  assign T289 = {T338, T290};
  assign T290 = T291;
  assign T291 = {T330, T292};
  assign T292 = T293;
  assign T293 = {T322, T294};
  assign T294 = T295;
  assign T295 = {T314, T296};
  assign T296 = T297;
  assign T297 = {T306, T298};
  assign T298 = T299;
  assign T299 = T300;
  assign T300 = T304[T301];
  assign T301 = T302;
  assign T302 = T303;
  assign T303 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T304 = T305;
  assign T305 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T306 = T307;
  assign T307 = T308;
  assign T308 = T312[T309];
  assign T309 = T310;
  assign T310 = T311;
  assign T311 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T312 = T313;
  assign T313 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T314 = T315;
  assign T315 = T316;
  assign T316 = T320[T317];
  assign T317 = T318;
  assign T318 = T319;
  assign T319 = io_chanxy_config[2'h2/* 2*/:2'h2/* 2*/];
  assign T320 = T321;
  assign T321 = io_chanxy_in[3'h5/* 5*/:3'h4/* 4*/];
  assign T322 = T323;
  assign T323 = T324;
  assign T324 = T328[T325];
  assign T325 = T326;
  assign T326 = T327;
  assign T327 = io_chanxy_config[2'h3/* 3*/:2'h3/* 3*/];
  assign T328 = T329;
  assign T329 = io_chanxy_in[3'h7/* 7*/:3'h6/* 6*/];
  assign T330 = T331;
  assign T331 = T332;
  assign T332 = T336[T333];
  assign T333 = T334;
  assign T334 = T335;
  assign T335 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T336 = T337;
  assign T337 = io_chanxy_in[5'h10/* 16*/:4'h8/* 8*/];
  assign T338 = T339;
  assign T339 = T340;
  assign T340 = T344[T341];
  assign T341 = T342;
  assign T342 = T343;
  assign T343 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T344 = T345;
  assign T345 = io_chanxy_in[5'h12/* 18*/:5'h11/* 17*/];
  assign T346 = T347;
  assign T347 = T348;
  assign T348 = T352[T349];
  assign T349 = T350;
  assign T350 = T351;
  assign T351 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T352 = T353;
  assign T353 = io_chanxy_in[5'h14/* 20*/:5'h13/* 19*/];
  assign T354 = T355;
  assign T355 = T356;
  assign T356 = T360[T357];
  assign T357 = T358;
  assign T358 = T359;
  assign T359 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T360 = T361;
  assign T361 = io_chanxy_in[5'h16/* 22*/:5'h15/* 21*/];
  assign T362 = T363;
  assign T363 = T364;
  assign T364 = T368[T365];
  assign T365 = T366;
  assign T366 = T367;
  assign T367 = io_chanxy_config[4'hb/* 11*/:4'hb/* 11*/];
  assign T368 = T369;
  assign T369 = io_chanxy_in[5'h18/* 24*/:5'h17/* 23*/];
  assign T370 = T371;
  assign T371 = T372;
  assign T372 = T376[T373];
  assign T373 = T374;
  assign T374 = T375;
  assign T375 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T376 = T377;
  assign T377 = io_chanxy_in[6'h21/* 33*/:5'h19/* 25*/];
  assign T378 = T379;
  assign T379 = T380;
  assign T380 = T384[T381];
  assign T381 = T382;
  assign T382 = T383;
  assign T383 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T384 = T385;
  assign T385 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T386 = T387;
  assign T387 = T388;
  assign T388 = T392[T389];
  assign T389 = T390;
  assign T390 = T391;
  assign T391 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T392 = T393;
  assign T393 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T394 = T395;
  assign T395 = T396;
  assign T396 = T400[T397];
  assign T397 = T398;
  assign T398 = T399;
  assign T399 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T400 = T401;
  assign T401 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T402 = T403;
  assign T403 = T404;
  assign T404 = T408[T405];
  assign T405 = T406;
  assign T406 = T407;
  assign T407 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T408 = T409;
  assign T409 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T410 = T411;
  assign T411 = T412;
  assign T412 = T416[T413];
  assign T413 = T414;
  assign T414 = T415;
  assign T415 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T416 = T417;
  assign T417 = io_chanxy_in[6'h32/* 50*/:6'h2a/* 42*/];
  assign T418 = T419;
  assign T419 = T420;
  assign T420 = T424[T421];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T424 = T425;
  assign T425 = io_chanxy_in[6'h34/* 52*/:6'h33/* 51*/];
  assign T426 = T427;
  assign T427 = T428;
  assign T428 = T432[T429];
  assign T429 = T430;
  assign T430 = T431;
  assign T431 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T432 = T433;
  assign T433 = io_chanxy_in[6'h36/* 54*/:6'h35/* 53*/];
  assign T434 = T435;
  assign T435 = T436;
  assign T436 = T440[T437];
  assign T437 = T438;
  assign T438 = T439;
  assign T439 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T440 = T441;
  assign T441 = io_chanxy_in[6'h38/* 56*/:6'h37/* 55*/];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = T448[T445];
  assign T445 = T446;
  assign T446 = T447;
  assign T447 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T448 = T449;
  assign T449 = io_chanxy_in[6'h3a/* 58*/:6'h39/* 57*/];
  assign T450 = T451;
  assign T451 = T452;
  assign T452 = T456[T453];
  assign T453 = T454;
  assign T454 = T455;
  assign T455 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T456 = T457;
  assign T457 = io_chanxy_in[7'h43/* 67*/:6'h3b/* 59*/];
  assign T458 = T459;
  assign T459 = T460;
  assign T460 = T464[T461];
  assign T461 = T462;
  assign T462 = T463;
  assign T463 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T464 = T465;
  assign T465 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T472[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T472 = T473;
  assign T473 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T474 = T475;
  assign T475 = T476;
  assign T476 = T480[T477];
  assign T477 = T478;
  assign T478 = T479;
  assign T479 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T480 = T481;
  assign T481 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T482 = T483;
  assign T483 = T484;
  assign T484 = T488[T485];
  assign T485 = T486;
  assign T486 = T487;
  assign T487 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T488 = T489;
  assign T489 = io_chanxy_in[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T490 = T491;
  assign T491 = T492;
  assign T492 = T496[T493];
  assign T493 = T494;
  assign T494 = T495;
  assign T495 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T496 = T497;
  assign T497 = io_chanxy_in[7'h54/* 84*/:7'h4c/* 76*/];
  assign T498 = T499;
  assign T499 = T500;
  assign T500 = T504[T501];
  assign T501 = T502;
  assign T502 = T503;
  assign T503 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T504 = T505;
  assign T505 = io_chanxy_in[7'h56/* 86*/:7'h55/* 85*/];
  assign T506 = T507;
  assign T507 = T508;
  assign T508 = T512[T509];
  assign T509 = T510;
  assign T510 = T511;
  assign T511 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T512 = T513;
  assign T513 = io_chanxy_in[7'h58/* 88*/:7'h57/* 87*/];
  assign T514 = T515;
  assign T515 = T516;
  assign T516 = T520[T517];
  assign T517 = T518;
  assign T518 = T519;
  assign T519 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T520 = T521;
  assign T521 = io_chanxy_in[7'h5a/* 90*/:7'h59/* 89*/];
  assign T522 = T523;
  assign T523 = T524;
  assign T524 = T528[T525];
  assign T525 = T526;
  assign T526 = T527;
  assign T527 = io_chanxy_config[6'h2b/* 43*/:6'h2b/* 43*/];
  assign T528 = T529;
  assign T529 = io_chanxy_in[7'h5c/* 92*/:7'h5b/* 91*/];
  assign T530 = T531;
  assign T531 = T532;
  assign T532 = T536[T533];
  assign T533 = T534;
  assign T534 = T535;
  assign T535 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T536 = T537;
  assign T537 = io_chanxy_in[7'h65/* 101*/:7'h5d/* 93*/];
  assign T538 = T539;
  assign T539 = T540;
  assign T540 = T544[T541];
  assign T541 = T542;
  assign T542 = T543;
  assign T543 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T544 = T545;
  assign T545 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T546 = T547;
  assign T547 = T548;
  assign T548 = T552[T549];
  assign T549 = T550;
  assign T550 = T551;
  assign T551 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T552 = T553;
  assign T553 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T554 = T555;
  assign T555 = T556;
  assign T556 = T560[T557];
  assign T557 = T558;
  assign T558 = T559;
  assign T559 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T560 = T561;
  assign T561 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T562 = T563;
  assign T563 = T564;
  assign T564 = T568[T565];
  assign T565 = T566;
  assign T566 = T567;
  assign T567 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T568 = T569;
  assign T569 = io_chanxy_in[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T570 = T571;
  assign T571 = T572;
  assign T572 = T576[T573];
  assign T573 = T574;
  assign T574 = T575;
  assign T575 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T576 = T577;
  assign T577 = io_chanxy_in[7'h76/* 118*/:7'h6e/* 110*/];
  assign T578 = T579;
  assign T579 = T580;
  assign T580 = T584[T581];
  assign T581 = T582;
  assign T582 = T583;
  assign T583 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T584 = T585;
  assign T585 = io_chanxy_in[7'h78/* 120*/:7'h77/* 119*/];
  assign T586 = T587;
  assign T587 = T588;
  assign T588 = T592[T589];
  assign T589 = T590;
  assign T590 = T591;
  assign T591 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T592 = T593;
  assign T593 = io_chanxy_in[7'h7a/* 122*/:7'h79/* 121*/];
  assign T594 = T595;
  assign T595 = T596;
  assign T596 = T600[T597];
  assign T597 = T598;
  assign T598 = T599;
  assign T599 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T600 = T601;
  assign T601 = io_chanxy_in[7'h7c/* 124*/:7'h7b/* 123*/];
  assign T602 = T603;
  assign T603 = T604;
  assign T604 = T608[T605];
  assign T605 = T606;
  assign T606 = T607;
  assign T607 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T608 = T609;
  assign T609 = io_chanxy_in[7'h7e/* 126*/:7'h7d/* 125*/];
  assign T610 = T611;
  assign T611 = T612;
  assign T612 = T616[T613];
  assign T613 = T614;
  assign T614 = T615;
  assign T615 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T616 = T617;
  assign T617 = io_chanxy_in[8'h87/* 135*/:7'h7f/* 127*/];
  assign T618 = T619;
  assign T619 = T620;
  assign T620 = T624[T621];
  assign T621 = T622;
  assign T622 = T623;
  assign T623 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T624 = T625;
  assign T625 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T626 = T627;
  assign T627 = T628;
  assign T628 = T632[T629];
  assign T629 = T630;
  assign T630 = T631;
  assign T631 = io_chanxy_config[7'h41/* 65*/:7'h41/* 65*/];
  assign T632 = T633;
  assign T633 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T634 = T635;
  assign T635 = T636;
  assign T636 = T640[T637];
  assign T637 = T638;
  assign T638 = T639;
  assign T639 = io_chanxy_config[7'h42/* 66*/:7'h42/* 66*/];
  assign T640 = T641;
  assign T641 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T642 = T643;
  assign T643 = T644;
  assign T644 = T648[T645];
  assign T645 = T646;
  assign T646 = T647;
  assign T647 = io_chanxy_config[7'h43/* 67*/:7'h43/* 67*/];
  assign T648 = T649;
  assign T649 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T650 = T651;
  assign T651 = T652;
  assign T652 = T656[T653];
  assign T653 = T654;
  assign T654 = T655;
  assign T655 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T656 = T657;
  assign T657 = io_chanxy_in[8'h98/* 152*/:8'h90/* 144*/];
  assign T658 = T659;
  assign T659 = T660;
  assign T660 = T664[T661];
  assign T661 = T662;
  assign T662 = T663;
  assign T663 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T664 = T665;
  assign T665 = io_chanxy_in[8'h9a/* 154*/:8'h99/* 153*/];
  assign T666 = T667;
  assign T667 = T668;
  assign T668 = T672[T669];
  assign T669 = T670;
  assign T670 = T671;
  assign T671 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T672 = T673;
  assign T673 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T674 = T675;
  assign T675 = T676;
  assign T676 = T680[T677];
  assign T677 = T678;
  assign T678 = T679;
  assign T679 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T680 = T681;
  assign T681 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T682 = T683;
  assign T683 = T684;
  assign T684 = T688[T685];
  assign T685 = T686;
  assign T686 = T687;
  assign T687 = io_chanxy_config[7'h4b/* 75*/:7'h4b/* 75*/];
  assign T688 = T689;
  assign T689 = io_chanxy_in[8'ha0/* 160*/:8'h9f/* 159*/];
  assign T690 = T691;
  assign T691 = T692;
  assign T692 = T696[T693];
  assign T693 = T694;
  assign T694 = T695;
  assign T695 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T696 = T697;
  assign T697 = io_chanxy_in[8'ha9/* 169*/:8'ha1/* 161*/];
  assign T698 = T699;
  assign T699 = T700;
  assign T700 = T704[T701];
  assign T701 = T702;
  assign T702 = T703;
  assign T703 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T704 = T705;
  assign T705 = io_chanxy_in[8'hab/* 171*/:8'haa/* 170*/];
  assign T706 = T707;
  assign T707 = T708;
  assign T708 = T712[T709];
  assign T709 = T710;
  assign T710 = T711;
  assign T711 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T712 = T713;
  assign T713 = io_chanxy_in[8'had/* 173*/:8'hac/* 172*/];
  assign T714 = T715;
  assign T715 = T716;
  assign T716 = T720[T717];
  assign T717 = T718;
  assign T718 = T719;
  assign T719 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T720 = T721;
  assign T721 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T722 = T723;
  assign T723 = T724;
  assign T724 = T728[T725];
  assign T725 = T726;
  assign T726 = T727;
  assign T727 = io_chanxy_config[7'h53/* 83*/:7'h53/* 83*/];
  assign T728 = T729;
  assign T729 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T730 = T731;
  assign T731 = T732;
  assign T732 = T736[T733];
  assign T733 = T734;
  assign T734 = T735;
  assign T735 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T736 = T737;
  assign T737 = io_chanxy_in[8'hba/* 186*/:8'hb2/* 178*/];
  assign T738 = T739;
  assign T739 = T740;
  assign T740 = T744[T741];
  assign T741 = T742;
  assign T742 = T743;
  assign T743 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T744 = T745;
  assign T745 = io_chanxy_in[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T746 = T747;
  assign T747 = T748;
  assign T748 = T752[T749];
  assign T749 = T750;
  assign T750 = T751;
  assign T751 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T752 = T753;
  assign T753 = io_chanxy_in[8'hbe/* 190*/:8'hbd/* 189*/];
  assign T754 = T755;
  assign T755 = T756;
  assign T756 = T760[T757];
  assign T757 = T758;
  assign T758 = T759;
  assign T759 = io_chanxy_config[7'h5a/* 90*/:7'h5a/* 90*/];
  assign T760 = T761;
  assign T761 = io_chanxy_in[8'hc0/* 192*/:8'hbf/* 191*/];
  assign T762 = T763;
  assign T763 = T764;
  assign T764 = T768[T765];
  assign T765 = T766;
  assign T766 = T767;
  assign T767 = io_chanxy_config[7'h5b/* 91*/:7'h5b/* 91*/];
  assign T768 = T769;
  assign T769 = io_chanxy_in[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T770 = T771;
  assign T771 = T772;
  assign T772 = T776[T773];
  assign T773 = T774;
  assign T774 = T775;
  assign T775 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T776 = T777;
  assign T777 = io_chanxy_in[8'hcb/* 203*/:8'hc3/* 195*/];
  assign T778 = T779;
  assign T779 = T780;
  assign T780 = T784[T781];
  assign T781 = T782;
  assign T782 = T783;
  assign T783 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T784 = T785;
  assign T785 = io_chanxy_in[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T786 = T787;
  assign T787 = T788;
  assign T788 = T792[T789];
  assign T789 = T790;
  assign T790 = T791;
  assign T791 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T792 = T793;
  assign T793 = io_chanxy_in[8'hcf/* 207*/:8'hce/* 206*/];
  assign T794 = T795;
  assign T795 = T796;
  assign T796 = T800[T797];
  assign T797 = T798;
  assign T798 = T799;
  assign T799 = io_chanxy_config[7'h62/* 98*/:7'h62/* 98*/];
  assign T800 = T801;
  assign T801 = io_chanxy_in[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T802 = T803;
  assign T803 = T804;
  assign T804 = T808[T805];
  assign T805 = T806;
  assign T806 = T807;
  assign T807 = io_chanxy_config[7'h63/* 99*/:7'h63/* 99*/];
  assign T808 = T809;
  assign T809 = io_chanxy_in[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T810 = T811;
  assign T811 = T812;
  assign T812 = T816[T813];
  assign T813 = T814;
  assign T814 = T815;
  assign T815 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T816 = T817;
  assign T817 = io_chanxy_in[8'hdc/* 220*/:8'hd4/* 212*/];
  assign T818 = T819;
  assign T819 = T820;
  assign T820 = T824[T821];
  assign T821 = T822;
  assign T822 = T823;
  assign T823 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T824 = T825;
  assign T825 = io_chanxy_in[8'hde/* 222*/:8'hdd/* 221*/];
  assign T826 = T827;
  assign T827 = T828;
  assign T828 = T832[T829];
  assign T829 = T830;
  assign T830 = T831;
  assign T831 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T832 = T833;
  assign T833 = io_chanxy_in[8'he0/* 224*/:8'hdf/* 223*/];
  assign T834 = T835;
  assign T835 = T836;
  assign T836 = T840[T837];
  assign T837 = T838;
  assign T838 = T839;
  assign T839 = io_chanxy_config[7'h6a/* 106*/:7'h6a/* 106*/];
  assign T840 = T841;
  assign T841 = io_chanxy_in[8'he2/* 226*/:8'he1/* 225*/];
  assign T842 = T843;
  assign T843 = T844;
  assign T844 = T848[T845];
  assign T845 = T846;
  assign T846 = T847;
  assign T847 = io_chanxy_config[7'h6b/* 107*/:7'h6b/* 107*/];
  assign T848 = T849;
  assign T849 = io_chanxy_in[8'he4/* 228*/:8'he3/* 227*/];
  assign T850 = T851;
  assign T851 = T852;
  assign T852 = T856[T853];
  assign T853 = T854;
  assign T854 = T855;
  assign T855 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T856 = T857;
  assign T857 = io_chanxy_in[8'hed/* 237*/:8'he5/* 229*/];
  assign T858 = T859;
  assign T859 = T860;
  assign T860 = T864[T861];
  assign T861 = T862;
  assign T862 = T863;
  assign T863 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T864 = T865;
  assign T865 = io_chanxy_in[8'hef/* 239*/:8'hee/* 238*/];
  assign T866 = T867;
  assign T867 = T868;
  assign T868 = T872[T869];
  assign T869 = T870;
  assign T870 = T871;
  assign T871 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T872 = T873;
  assign T873 = io_chanxy_in[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T874 = T875;
  assign T875 = T876;
  assign T876 = T880[T877];
  assign T877 = T878;
  assign T878 = T879;
  assign T879 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T880 = T881;
  assign T881 = io_chanxy_in[8'hf3/* 243*/:8'hf2/* 242*/];
  assign T882 = T883;
  assign T883 = T884;
  assign T884 = T888[T885];
  assign T885 = T886;
  assign T886 = T887;
  assign T887 = io_chanxy_config[7'h73/* 115*/:7'h73/* 115*/];
  assign T888 = T889;
  assign T889 = io_chanxy_in[8'hf5/* 245*/:8'hf4/* 244*/];
  assign T890 = T891;
  assign T891 = T892;
  assign T892 = T896[T893];
  assign T893 = T894;
  assign T894 = T895;
  assign T895 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T896 = T897;
  assign T897 = io_chanxy_in[8'hfe/* 254*/:8'hf6/* 246*/];
  assign T898 = T899;
  assign T899 = T900;
  assign T900 = T904[T901];
  assign T901 = T902;
  assign T902 = T903;
  assign T903 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T904 = T905;
  assign T905 = io_chanxy_in[9'h101/* 257*/:8'hff/* 255*/];
  assign T906 = T907;
  assign T907 = T908;
  assign T908 = T912[T909];
  assign T909 = T910;
  assign T910 = T911;
  assign T911 = io_chanxy_config[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T912 = T913;
  assign T913 = io_chanxy_in[9'h104/* 260*/:9'h102/* 258*/];
  assign T914 = T915;
  assign T915 = T916;
  assign T916 = T920[T917];
  assign T917 = T918;
  assign T918 = T919;
  assign T919 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T920 = T921;
  assign T921 = io_chanxy_in[9'h107/* 263*/:9'h105/* 261*/];
  assign T922 = T923;
  assign T923 = T924;
  assign T924 = T928[T925];
  assign T925 = T926;
  assign T926 = T927;
  assign T927 = io_chanxy_config[7'h7f/* 127*/:7'h7e/* 126*/];
  assign T928 = T929;
  assign T929 = io_chanxy_in[9'h10a/* 266*/:9'h108/* 264*/];
  assign T930 = T931;
  assign T931 = T932;
  assign T932 = T936[T933];
  assign T933 = T934;
  assign T934 = T935;
  assign T935 = io_chanxy_config[8'h81/* 129*/:8'h80/* 128*/];
  assign T936 = T937;
  assign T937 = io_chanxy_in[9'h10d/* 269*/:9'h10b/* 267*/];
  assign T938 = T939;
  assign T939 = T940;
  assign T940 = T944[T941];
  assign T941 = T942;
  assign T942 = T943;
  assign T943 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T944 = T945;
  assign T945 = io_chanxy_in[9'h110/* 272*/:9'h10e/* 270*/];
  assign T946 = T947;
  assign T947 = T948;
  assign T948 = T952[T949];
  assign T949 = T950;
  assign T950 = T951;
  assign T951 = io_chanxy_config[8'h84/* 132*/:8'h84/* 132*/];
  assign T952 = T953;
  assign T953 = io_chanxy_in[9'h112/* 274*/:9'h111/* 273*/];
  assign T954 = T955;
  assign T955 = T956;
  assign T956 = T960[T957];
  assign T957 = T958;
  assign T958 = T959;
  assign T959 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T960 = T961;
  assign T961 = io_chanxy_in[9'h114/* 276*/:9'h113/* 275*/];
  assign T962 = T963;
  assign T963 = T964;
  assign T964 = T968[T965];
  assign T965 = T966;
  assign T966 = T967;
  assign T967 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T968 = T969;
  assign T969 = io_chanxy_in[9'h116/* 278*/:9'h115/* 277*/];
  assign T970 = T971;
  assign T971 = T972;
  assign T972 = T976[T973];
  assign T973 = T974;
  assign T974 = T975;
  assign T975 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T976 = T977;
  assign T977 = io_chanxy_in[9'h118/* 280*/:9'h117/* 279*/];
  assign T978 = T979;
  assign T979 = T980;
  assign T980 = T984[T981];
  assign T981 = T982;
  assign T982 = T983;
  assign T983 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T984 = T985;
  assign T985 = io_chanxy_in[9'h11a/* 282*/:9'h119/* 281*/];
  assign T986 = T987;
  assign T987 = T988;
  assign T988 = T992[T989];
  assign T989 = T990;
  assign T990 = T991;
  assign T991 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T992 = T993;
  assign T993 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T994 = T995;
  assign T995 = T996;
  assign T996 = T1000[T997];
  assign T997 = T998;
  assign T998 = T999;
  assign T999 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T1000 = T1001;
  assign T1001 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T1002 = T1003;
  assign T1003 = T1004;
  assign T1004 = T1008[T1005];
  assign T1005 = T1006;
  assign T1006 = T1007;
  assign T1007 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T1008 = T1009;
  assign T1009 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T1010 = T1011;
  assign T1011 = T1012;
  assign T1012 = T1016[T1013];
  assign T1013 = T1014;
  assign T1014 = T1015;
  assign T1015 = io_chanxy_config[8'h8c/* 140*/:8'h8c/* 140*/];
  assign T1016 = T1017;
  assign T1017 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T1018 = T1019;
  assign T1019 = T1020;
  assign T1020 = T1024[T1021];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = io_chanxy_config[8'h8e/* 142*/:8'h8d/* 141*/];
  assign T1024 = T1025;
  assign T1025 = io_chanxy_in[9'h125/* 293*/:9'h123/* 291*/];
  assign T1026 = T1027;
  assign T1027 = T1028;
  assign T1028 = T1032[T1029];
  assign T1029 = T1030;
  assign T1030 = T1031;
  assign T1031 = io_chanxy_config[8'h90/* 144*/:8'h8f/* 143*/];
  assign T1032 = T1033;
  assign T1033 = io_chanxy_in[9'h128/* 296*/:9'h126/* 294*/];
  assign T1034 = T1035;
  assign T1035 = T1036;
  assign T1036 = T1040[T1037];
  assign T1037 = T1038;
  assign T1038 = T1039;
  assign T1039 = io_chanxy_config[8'h92/* 146*/:8'h91/* 145*/];
  assign T1040 = T1041;
  assign T1041 = io_chanxy_in[9'h12b/* 299*/:9'h129/* 297*/];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = T1048[T1045];
  assign T1045 = T1046;
  assign T1046 = T1047;
  assign T1047 = io_chanxy_config[8'h94/* 148*/:8'h93/* 147*/];
  assign T1048 = T1049;
  assign T1049 = io_chanxy_in[9'h12e/* 302*/:9'h12c/* 300*/];
  assign T1050 = T1051;
  assign T1051 = T1052;
  assign T1052 = T1056[T1053];
  assign T1053 = T1054;
  assign T1054 = T1055;
  assign T1055 = io_chanxy_config[8'h96/* 150*/:8'h95/* 149*/];
  assign T1056 = T1057;
  assign T1057 = io_chanxy_in[9'h131/* 305*/:9'h12f/* 303*/];
  assign T1058 = T1059;
  assign T1059 = T1060;
  assign T1060 = T1064[T1061];
  assign T1061 = T1062;
  assign T1062 = T1063;
  assign T1063 = io_chanxy_config[8'h98/* 152*/:8'h97/* 151*/];
  assign T1064 = T1065;
  assign T1065 = io_chanxy_in[9'h134/* 308*/:9'h132/* 306*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1072[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T1072 = T1073;
  assign T1073 = io_chanxy_in[9'h136/* 310*/:9'h135/* 309*/];
  assign T1074 = T1075;
  assign T1075 = T1076;
  assign T1076 = T1080[T1077];
  assign T1077 = T1078;
  assign T1078 = T1079;
  assign T1079 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T1080 = T1081;
  assign T1081 = io_chanxy_in[9'h138/* 312*/:9'h137/* 311*/];
  assign T1082 = T1083;
  assign T1083 = T1084;
  assign T1084 = T1088[T1085];
  assign T1085 = T1086;
  assign T1086 = T1087;
  assign T1087 = io_chanxy_config[8'h9b/* 155*/:8'h9b/* 155*/];
  assign T1088 = T1089;
  assign T1089 = io_chanxy_in[9'h13a/* 314*/:9'h139/* 313*/];
  assign T1090 = T1091;
  assign T1091 = T1092;
  assign T1092 = T1096[T1093];
  assign T1093 = T1094;
  assign T1094 = T1095;
  assign T1095 = io_chanxy_config[8'h9c/* 156*/:8'h9c/* 156*/];
  assign T1096 = T1097;
  assign T1097 = io_chanxy_in[9'h13c/* 316*/:9'h13b/* 315*/];
  assign T1098 = T1099;
  assign T1099 = T1100;
  assign T1100 = T1104[T1101];
  assign T1101 = T1102;
  assign T1102 = T1103;
  assign T1103 = io_chanxy_config[8'h9d/* 157*/:8'h9d/* 157*/];
  assign T1104 = T1105;
  assign T1105 = io_chanxy_in[9'h13e/* 318*/:9'h13d/* 317*/];
  assign T1106 = T1107;
  assign T1107 = T1108;
  assign T1108 = T1112[T1109];
  assign T1109 = T1110;
  assign T1110 = T1111;
  assign T1111 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T1112 = T1113;
  assign T1113 = io_chanxy_in[9'h140/* 320*/:9'h13f/* 319*/];
  assign T1114 = T1115;
  assign T1115 = T1116;
  assign T1116 = T1120[T1117];
  assign T1117 = T1118;
  assign T1118 = T1119;
  assign T1119 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T1120 = T1121;
  assign T1121 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T1122 = T1123;
  assign T1123 = T1124;
  assign T1124 = T1128[T1125];
  assign T1125 = T1126;
  assign T1126 = T1127;
  assign T1127 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T1128 = T1129;
  assign T1129 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T1130 = T1131;
  assign T1131 = T1132;
  assign T1132 = T1136[T1133];
  assign T1133 = T1134;
  assign T1134 = T1135;
  assign T1135 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T1136 = T1137;
  assign T1137 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T1138 = T1139;
  assign T1139 = T1140;
  assign T1140 = T1144[T1141];
  assign T1141 = T1142;
  assign T1142 = T1143;
  assign T1143 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T1144 = T1145;
  assign T1145 = io_chanxy_in[9'h149/* 329*/:9'h147/* 327*/];
  assign T1146 = T1147;
  assign T1147 = T1148;
  assign T1148 = T1152[T1149];
  assign T1149 = T1150;
  assign T1150 = T1151;
  assign T1151 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T1152 = T1153;
  assign T1153 = io_chanxy_in[9'h14c/* 332*/:9'h14a/* 330*/];
  assign T1154 = T1155;
  assign T1155 = T1156;
  assign T1156 = T1160[T1157];
  assign T1157 = T1158;
  assign T1158 = T1159;
  assign T1159 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T1160 = T1161;
  assign T1161 = io_chanxy_in[9'h14f/* 335*/:9'h14d/* 333*/];
  assign T1162 = T1163;
  assign T1163 = T1164;
  assign T1164 = T1168[T1165];
  assign T1165 = T1166;
  assign T1166 = T1167;
  assign T1167 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T1168 = T1169;
  assign T1169 = io_chanxy_in[9'h152/* 338*/:9'h150/* 336*/];
  assign T1170 = T1171;
  assign T1171 = T1172;
  assign T1172 = T1176[T1173];
  assign T1173 = T1174;
  assign T1174 = T1175;
  assign T1175 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T1176 = T1177;
  assign T1177 = io_chanxy_in[9'h155/* 341*/:9'h153/* 339*/];
  assign T1178 = T1179;
  assign T1179 = T1180;
  assign T1180 = T1184[T1181];
  assign T1181 = T1182;
  assign T1182 = T1183;
  assign T1183 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T1184 = T1185;
  assign T1185 = io_chanxy_in[9'h158/* 344*/:9'h156/* 342*/];
  assign T1186 = T1187;
  assign T1187 = T1188;
  assign T1188 = T1192[T1189];
  assign T1189 = T1190;
  assign T1190 = T1191;
  assign T1191 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T1192 = T1193;
  assign T1193 = io_chanxy_in[9'h15a/* 346*/:9'h159/* 345*/];
  assign T1194 = T1195;
  assign T1195 = T1196;
  assign T1196 = T1200[T1197];
  assign T1197 = T1198;
  assign T1198 = T1199;
  assign T1199 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T1200 = T1201;
  assign T1201 = io_chanxy_in[9'h15c/* 348*/:9'h15b/* 347*/];
  assign T1202 = T1203;
  assign T1203 = T1204;
  assign T1204 = T1208[T1205];
  assign T1205 = T1206;
  assign T1206 = T1207;
  assign T1207 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T1208 = T1209;
  assign T1209 = io_chanxy_in[9'h15e/* 350*/:9'h15d/* 349*/];
  assign T1210 = T1211;
  assign T1211 = T1212;
  assign T1212 = T1216[T1213];
  assign T1213 = T1214;
  assign T1214 = T1215;
  assign T1215 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T1216 = T1217;
  assign T1217 = io_chanxy_in[9'h160/* 352*/:9'h15f/* 351*/];
  assign T1218 = T1219;
  assign T1219 = T1220;
  assign T1220 = T1224[T1221];
  assign T1221 = T1222;
  assign T1222 = T1223;
  assign T1223 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T1224 = T1225;
  assign T1225 = io_chanxy_in[9'h162/* 354*/:9'h161/* 353*/];
  assign T1226 = T1227;
  assign T1227 = T1228;
  assign T1228 = T1232[T1229];
  assign T1229 = T1230;
  assign T1230 = T1231;
  assign T1231 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1232 = T1233;
  assign T1233 = io_chanxy_in[9'h164/* 356*/:9'h163/* 355*/];
  assign T1234 = T1235;
  assign T1235 = T1236;
  assign T1236 = T1240[T1237];
  assign T1237 = T1238;
  assign T1238 = T1239;
  assign T1239 = io_chanxy_config[8'hb4/* 180*/:8'hb4/* 180*/];
  assign T1240 = T1241;
  assign T1241 = io_chanxy_in[9'h166/* 358*/:9'h165/* 357*/];
  assign T1242 = T1243;
  assign T1243 = T1244;
  assign T1244 = T1248[T1245];
  assign T1245 = T1246;
  assign T1246 = T1247;
  assign T1247 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T1248 = T1249;
  assign T1249 = io_chanxy_in[9'h168/* 360*/:9'h167/* 359*/];
  assign T1250 = T1251;
  assign T1251 = T1252;
  assign T1252 = T1256[T1253];
  assign T1253 = T1254;
  assign T1254 = T1255;
  assign T1255 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T1256 = T1257;
  assign T1257 = io_chanxy_in[9'h16a/* 362*/:9'h169/* 361*/];
  assign T1258 = T1259;
  assign T1259 = T1260;
  assign T1260 = T1264[T1261];
  assign T1261 = T1262;
  assign T1262 = T1263;
  assign T1263 = io_chanxy_config[8'hba/* 186*/:8'hb7/* 183*/];
  assign T1264 = T1265;
  assign T1265 = io_chanxy_in[9'h175/* 373*/:9'h16b/* 363*/];
  assign T1266 = T1267;
  assign T1267 = T1268;
  assign T1268 = T1272[T1269];
  assign T1269 = T1270;
  assign T1270 = T1271;
  assign T1271 = io_chanxy_config[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T1272 = T1273;
  assign T1273 = io_chanxy_in[9'h178/* 376*/:9'h176/* 374*/];
  assign T1274 = T1275;
  assign T1275 = T1276;
  assign T1276 = T1280[T1277];
  assign T1277 = T1278;
  assign T1278 = T1279;
  assign T1279 = io_chanxy_config[8'hc0/* 192*/:8'hbd/* 189*/];
  assign T1280 = T1281;
  assign T1281 = io_chanxy_in[9'h183/* 387*/:9'h179/* 377*/];
  assign T1282 = T1283;
  assign T1283 = T1284;
  assign T1284 = T1288[T1285];
  assign T1285 = T1286;
  assign T1286 = T1287;
  assign T1287 = io_chanxy_config[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T1288 = T1289;
  assign T1289 = io_chanxy_in[9'h186/* 390*/:9'h184/* 388*/];
  assign T1290 = T1291;
  assign T1291 = T1292;
  assign T1292 = T1296[T1293];
  assign T1293 = T1294;
  assign T1294 = T1295;
  assign T1295 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T1296 = T1297;
  assign T1297 = io_chanxy_in[9'h191/* 401*/:9'h187/* 391*/];
  assign T1298 = T1299;
  assign T1299 = T1300;
  assign T1300 = T1304[T1301];
  assign T1301 = T1302;
  assign T1302 = T1303;
  assign T1303 = io_chanxy_config[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T1304 = T1305;
  assign T1305 = io_chanxy_in[9'h194/* 404*/:9'h192/* 402*/];
  assign T1306 = T1307;
  assign T1307 = T1308;
  assign T1308 = T1312[T1309];
  assign T1309 = T1310;
  assign T1310 = T1311;
  assign T1311 = io_chanxy_config[8'hcc/* 204*/:8'hc9/* 201*/];
  assign T1312 = T1313;
  assign T1313 = io_chanxy_in[9'h19f/* 415*/:9'h195/* 405*/];
  assign T1314 = T1315;
  assign T1315 = T1316;
  assign T1316 = T1320[T1317];
  assign T1317 = T1318;
  assign T1318 = T1319;
  assign T1319 = io_chanxy_config[8'hce/* 206*/:8'hcd/* 205*/];
  assign T1320 = T1321;
  assign T1321 = io_chanxy_in[9'h1a2/* 418*/:9'h1a0/* 416*/];
  assign T1322 = T1323;
  assign T1323 = T1324;
  assign T1324 = T1328[T1325];
  assign T1325 = T1326;
  assign T1326 = T1327;
  assign T1327 = io_chanxy_config[8'hd2/* 210*/:8'hcf/* 207*/];
  assign T1328 = T1329;
  assign T1329 = io_chanxy_in[9'h1ad/* 429*/:9'h1a3/* 419*/];
  assign T1330 = T1331;
  assign T1331 = T1332;
  assign T1332 = T1336[T1333];
  assign T1333 = T1334;
  assign T1334 = T1335;
  assign T1335 = io_chanxy_config[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T1336 = T1337;
  assign T1337 = io_chanxy_in[9'h1b0/* 432*/:9'h1ae/* 430*/];
  assign T1338 = T1339;
  assign T1339 = T1340;
  assign T1340 = T1344[T1341];
  assign T1341 = T1342;
  assign T1342 = T1343;
  assign T1343 = io_chanxy_config[8'hd8/* 216*/:8'hd5/* 213*/];
  assign T1344 = T1345;
  assign T1345 = io_chanxy_in[9'h1bb/* 443*/:9'h1b1/* 433*/];
  assign T1346 = T1347;
  assign T1347 = T1348;
  assign T1348 = T1352[T1349];
  assign T1349 = T1350;
  assign T1350 = T1351;
  assign T1351 = io_chanxy_config[8'hda/* 218*/:8'hd9/* 217*/];
  assign T1352 = T1353;
  assign T1353 = io_chanxy_in[9'h1be/* 446*/:9'h1bc/* 444*/];
  assign T1354 = T1355;
  assign T1355 = T1356;
  assign T1356 = T1360[T1357];
  assign T1357 = T1358;
  assign T1358 = T1359;
  assign T1359 = io_chanxy_config[8'hde/* 222*/:8'hdb/* 219*/];
  assign T1360 = T1361;
  assign T1361 = io_chanxy_in[9'h1c9/* 457*/:9'h1bf/* 447*/];
  assign T1362 = T1363;
  assign T1363 = T1364;
  assign T1364 = T1368[T1365];
  assign T1365 = T1366;
  assign T1366 = T1367;
  assign T1367 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T1368 = T1369;
  assign T1369 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T1370 = T1371;
  assign T1371 = T1372;
  assign T1372 = T1376[T1373];
  assign T1373 = T1374;
  assign T1374 = T1375;
  assign T1375 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T1376 = T1377;
  assign T1377 = io_chanxy_in[9'h1d6/* 470*/:9'h1cc/* 460*/];
  assign T1378 = T1379;
  assign T1379 = T1380;
  assign T1380 = T1384[T1381];
  assign T1381 = T1382;
  assign T1382 = T1383;
  assign T1383 = io_chanxy_config[8'he4/* 228*/:8'he4/* 228*/];
  assign T1384 = T1385;
  assign T1385 = io_chanxy_in[9'h1d8/* 472*/:9'h1d7/* 471*/];
  assign T1386 = T1387;
  assign T1387 = T1388;
  assign T1388 = T1392[T1389];
  assign T1389 = T1390;
  assign T1390 = T1391;
  assign T1391 = io_chanxy_config[8'he8/* 232*/:8'he5/* 229*/];
  assign T1392 = T1393;
  assign T1393 = io_chanxy_in[9'h1e3/* 483*/:9'h1d9/* 473*/];
  assign T1394 = T1395;
  assign T1395 = T1396;
  assign T1396 = T1400[T1397];
  assign T1397 = T1398;
  assign T1398 = T1399;
  assign T1399 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T1400 = T1401;
  assign T1401 = io_chanxy_in[9'h1e5/* 485*/:9'h1e4/* 484*/];
  assign T1402 = T1403;
  assign T1403 = T1404;
  assign T1404 = T1408[T1405];
  assign T1405 = T1406;
  assign T1406 = T1407;
  assign T1407 = io_chanxy_config[8'hed/* 237*/:8'hea/* 234*/];
  assign T1408 = T1409;
  assign T1409 = io_chanxy_in[9'h1ef/* 495*/:9'h1e6/* 486*/];
  assign T1410 = T1411;
  assign T1411 = T1412;
  assign T1412 = T1416[T1413];
  assign T1413 = T1414;
  assign T1414 = T1415;
  assign T1415 = io_chanxy_config[8'hee/* 238*/:8'hee/* 238*/];
  assign T1416 = T1417;
  assign T1417 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T1418 = T1419;
  assign T1419 = T1420;
  assign T1420 = T1424[T1421];
  assign T1421 = T1422;
  assign T1422 = T1423;
  assign T1423 = io_chanxy_config[8'hf2/* 242*/:8'hef/* 239*/];
  assign T1424 = T1425;
  assign T1425 = io_chanxy_in[9'h1fb/* 507*/:9'h1f2/* 498*/];
  assign T1426 = T1427;
  assign T1427 = T1428;
  assign T1428 = T1432[T1429];
  assign T1429 = T1430;
  assign T1430 = T1431;
  assign T1431 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T1432 = T1433;
  assign T1433 = io_chanxy_in[9'h1fd/* 509*/:9'h1fc/* 508*/];
  assign T1434 = T1435;
  assign T1435 = T1436;
  assign T1436 = T1440[T1437];
  assign T1437 = T1438;
  assign T1438 = T1439;
  assign T1439 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1440 = T1441;
  assign T1441 = io_chanxy_in[10'h207/* 519*/:9'h1fe/* 510*/];
  assign T1442 = T1443;
  assign T1443 = T1444;
  assign T1444 = T1448[T1445];
  assign T1445 = T1446;
  assign T1446 = T1447;
  assign T1447 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1448 = T1449;
  assign T1449 = io_chanxy_in[10'h209/* 521*/:10'h208/* 520*/];
  assign T1450 = T1451;
  assign T1451 = T1452;
  assign T1452 = T1456[T1453];
  assign T1453 = T1454;
  assign T1454 = T1455;
  assign T1455 = io_chanxy_config[8'hfc/* 252*/:8'hf9/* 249*/];
  assign T1456 = T1457;
  assign T1457 = io_chanxy_in[10'h213/* 531*/:10'h20a/* 522*/];
  assign T1458 = T1459;
  assign T1459 = T1460;
  assign T1460 = T1464[T1461];
  assign T1461 = T1462;
  assign T1462 = T1463;
  assign T1463 = io_chanxy_config[8'hfd/* 253*/:8'hfd/* 253*/];
  assign T1464 = T1465;
  assign T1465 = io_chanxy_in[10'h215/* 533*/:10'h214/* 532*/];
  assign T1466 = T1467;
  assign T1467 = T1468;
  assign T1468 = T1472[T1469];
  assign T1469 = T1470;
  assign T1470 = T1471;
  assign T1471 = io_chanxy_config[9'h101/* 257*/:8'hfe/* 254*/];
  assign T1472 = T1473;
  assign T1473 = io_chanxy_in[10'h21f/* 543*/:10'h216/* 534*/];
  assign T1474 = T1475;
  assign T1475 = T1476;
  assign T1476 = T1480[T1477];
  assign T1477 = T1478;
  assign T1478 = T1479;
  assign T1479 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1480 = T1481;
  assign T1481 = io_chanxy_in[10'h221/* 545*/:10'h220/* 544*/];
  assign T1482 = T1483;
  assign T1483 = T1484;
  assign T1484 = T1488[T1485];
  assign T1485 = T1486;
  assign T1486 = T1487;
  assign T1487 = io_chanxy_config[9'h106/* 262*/:9'h103/* 259*/];
  assign T1488 = T1489;
  assign T1489 = io_chanxy_in[10'h22b/* 555*/:10'h222/* 546*/];
  assign T1490 = T1491;
  assign T1491 = T1492;
  assign T1492 = T1496[T1493];
  assign T1493 = T1494;
  assign T1494 = T1495;
  assign T1495 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1496 = T1497;
  assign T1497 = io_chanxy_in[10'h22d/* 557*/:10'h22c/* 556*/];
  assign io_ipin_out = T1498;
  assign T1498 = T1499;
  assign T1499 = {T1718, T1500};
  assign T1500 = T1501;
  assign T1501 = {T1710, T1502};
  assign T1502 = T1503;
  assign T1503 = {T1702, T1504};
  assign T1504 = T1505;
  assign T1505 = {T1694, T1506};
  assign T1506 = T1507;
  assign T1507 = {T1686, T1508};
  assign T1508 = T1509;
  assign T1509 = {T1678, T1510};
  assign T1510 = T1511;
  assign T1511 = {T1670, T1512};
  assign T1512 = T1513;
  assign T1513 = {T1662, T1514};
  assign T1514 = T1515;
  assign T1515 = {T1654, T1516};
  assign T1516 = T1517;
  assign T1517 = {T1646, T1518};
  assign T1518 = T1519;
  assign T1519 = {T1638, T1520};
  assign T1520 = T1521;
  assign T1521 = {T1630, T1522};
  assign T1522 = T1523;
  assign T1523 = {T1622, T1524};
  assign T1524 = T1525;
  assign T1525 = {T1614, T1526};
  assign T1526 = T1527;
  assign T1527 = {T1606, T1528};
  assign T1528 = T1529;
  assign T1529 = {T1598, T1530};
  assign T1530 = T1531;
  assign T1531 = {T1590, T1532};
  assign T1532 = T1533;
  assign T1533 = {T1582, T1534};
  assign T1534 = T1535;
  assign T1535 = {T1574, T1536};
  assign T1536 = T1537;
  assign T1537 = {T1566, T1538};
  assign T1538 = T1539;
  assign T1539 = {T1558, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1550, T1542};
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_9(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [557:0] io_chanxy_in,
    output[149:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[149:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_5 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_6(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [557:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[149:0] io_chanxy_out);

  wire[149:0] T0;
  wire[149:0] T1;
  wire[148:0] T2;
  wire[148:0] T3;
  wire[147:0] T4;
  wire[147:0] T5;
  wire[146:0] T6;
  wire[146:0] T7;
  wire[145:0] T8;
  wire[145:0] T9;
  wire[144:0] T10;
  wire[144:0] T11;
  wire[143:0] T12;
  wire[143:0] T13;
  wire[142:0] T14;
  wire[142:0] T15;
  wire[141:0] T16;
  wire[141:0] T17;
  wire[140:0] T18;
  wire[140:0] T19;
  wire[139:0] T20;
  wire[139:0] T21;
  wire[138:0] T22;
  wire[138:0] T23;
  wire[137:0] T24;
  wire[137:0] T25;
  wire[136:0] T26;
  wire[136:0] T27;
  wire[135:0] T28;
  wire[135:0] T29;
  wire[134:0] T30;
  wire[134:0] T31;
  wire[133:0] T32;
  wire[133:0] T33;
  wire[132:0] T34;
  wire[132:0] T35;
  wire[131:0] T36;
  wire[131:0] T37;
  wire[130:0] T38;
  wire[130:0] T39;
  wire[129:0] T40;
  wire[129:0] T41;
  wire[128:0] T42;
  wire[128:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[126:0] T46;
  wire[126:0] T47;
  wire[125:0] T48;
  wire[125:0] T49;
  wire[124:0] T50;
  wire[124:0] T51;
  wire[123:0] T52;
  wire[123:0] T53;
  wire[122:0] T54;
  wire[122:0] T55;
  wire[121:0] T56;
  wire[121:0] T57;
  wire[120:0] T58;
  wire[120:0] T59;
  wire[119:0] T60;
  wire[119:0] T61;
  wire[118:0] T62;
  wire[118:0] T63;
  wire[117:0] T64;
  wire[117:0] T65;
  wire[116:0] T66;
  wire[116:0] T67;
  wire[115:0] T68;
  wire[115:0] T69;
  wire[114:0] T70;
  wire[114:0] T71;
  wire[113:0] T72;
  wire[113:0] T73;
  wire[112:0] T74;
  wire[112:0] T75;
  wire[111:0] T76;
  wire[111:0] T77;
  wire[110:0] T78;
  wire[110:0] T79;
  wire[109:0] T80;
  wire[109:0] T81;
  wire[108:0] T82;
  wire[108:0] T83;
  wire[107:0] T84;
  wire[107:0] T85;
  wire[106:0] T86;
  wire[106:0] T87;
  wire[105:0] T88;
  wire[105:0] T89;
  wire[104:0] T90;
  wire[104:0] T91;
  wire[103:0] T92;
  wire[103:0] T93;
  wire[102:0] T94;
  wire[102:0] T95;
  wire[101:0] T96;
  wire[101:0] T97;
  wire[100:0] T98;
  wire[100:0] T99;
  wire[99:0] T100;
  wire[99:0] T101;
  wire[98:0] T102;
  wire[98:0] T103;
  wire[97:0] T104;
  wire[97:0] T105;
  wire[96:0] T106;
  wire[96:0] T107;
  wire[95:0] T108;
  wire[95:0] T109;
  wire[94:0] T110;
  wire[94:0] T111;
  wire[93:0] T112;
  wire[93:0] T113;
  wire[92:0] T114;
  wire[92:0] T115;
  wire[91:0] T116;
  wire[91:0] T117;
  wire[90:0] T118;
  wire[90:0] T119;
  wire[89:0] T120;
  wire[89:0] T121;
  wire[88:0] T122;
  wire[88:0] T123;
  wire[87:0] T124;
  wire[87:0] T125;
  wire[86:0] T126;
  wire[86:0] T127;
  wire[85:0] T128;
  wire[85:0] T129;
  wire[84:0] T130;
  wire[84:0] T131;
  wire[83:0] T132;
  wire[83:0] T133;
  wire[82:0] T134;
  wire[82:0] T135;
  wire[81:0] T136;
  wire[81:0] T137;
  wire[80:0] T138;
  wire[80:0] T139;
  wire[79:0] T140;
  wire[79:0] T141;
  wire[78:0] T142;
  wire[78:0] T143;
  wire[77:0] T144;
  wire[77:0] T145;
  wire[76:0] T146;
  wire[76:0] T147;
  wire[75:0] T148;
  wire[75:0] T149;
  wire[74:0] T150;
  wire[74:0] T151;
  wire[73:0] T152;
  wire[73:0] T153;
  wire[72:0] T154;
  wire[72:0] T155;
  wire[71:0] T156;
  wire[71:0] T157;
  wire[70:0] T158;
  wire[70:0] T159;
  wire[69:0] T160;
  wire[69:0] T161;
  wire[68:0] T162;
  wire[68:0] T163;
  wire[67:0] T164;
  wire[67:0] T165;
  wire[66:0] T166;
  wire[66:0] T167;
  wire[65:0] T168;
  wire[65:0] T169;
  wire[64:0] T170;
  wire[64:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[62:0] T174;
  wire[62:0] T175;
  wire[61:0] T176;
  wire[61:0] T177;
  wire[60:0] T178;
  wire[60:0] T179;
  wire[59:0] T180;
  wire[59:0] T181;
  wire[58:0] T182;
  wire[58:0] T183;
  wire[57:0] T184;
  wire[57:0] T185;
  wire[56:0] T186;
  wire[56:0] T187;
  wire[55:0] T188;
  wire[55:0] T189;
  wire[54:0] T190;
  wire[54:0] T191;
  wire[53:0] T192;
  wire[53:0] T193;
  wire[52:0] T194;
  wire[52:0] T195;
  wire[51:0] T196;
  wire[51:0] T197;
  wire[50:0] T198;
  wire[50:0] T199;
  wire[49:0] T200;
  wire[49:0] T201;
  wire[48:0] T202;
  wire[48:0] T203;
  wire[47:0] T204;
  wire[47:0] T205;
  wire[46:0] T206;
  wire[46:0] T207;
  wire[45:0] T208;
  wire[45:0] T209;
  wire[44:0] T210;
  wire[44:0] T211;
  wire[43:0] T212;
  wire[43:0] T213;
  wire[42:0] T214;
  wire[42:0] T215;
  wire[41:0] T216;
  wire[41:0] T217;
  wire[40:0] T218;
  wire[40:0] T219;
  wire[39:0] T220;
  wire[39:0] T221;
  wire[38:0] T222;
  wire[38:0] T223;
  wire[37:0] T224;
  wire[37:0] T225;
  wire[36:0] T226;
  wire[36:0] T227;
  wire[35:0] T228;
  wire[35:0] T229;
  wire[34:0] T230;
  wire[34:0] T231;
  wire[33:0] T232;
  wire[33:0] T233;
  wire[32:0] T234;
  wire[32:0] T235;
  wire[31:0] T236;
  wire[31:0] T237;
  wire[30:0] T238;
  wire[30:0] T239;
  wire[29:0] T240;
  wire[29:0] T241;
  wire[28:0] T242;
  wire[28:0] T243;
  wire[27:0] T244;
  wire[27:0] T245;
  wire[26:0] T246;
  wire[26:0] T247;
  wire[25:0] T248;
  wire[25:0] T249;
  wire[24:0] T250;
  wire[24:0] T251;
  wire[23:0] T252;
  wire[23:0] T253;
  wire[22:0] T254;
  wire[22:0] T255;
  wire[21:0] T256;
  wire[21:0] T257;
  wire[20:0] T258;
  wire[20:0] T259;
  wire[19:0] T260;
  wire[19:0] T261;
  wire[18:0] T262;
  wire[18:0] T263;
  wire[17:0] T264;
  wire[17:0] T265;
  wire[16:0] T266;
  wire[16:0] T267;
  wire[15:0] T268;
  wire[15:0] T269;
  wire[14:0] T270;
  wire[14:0] T271;
  wire[13:0] T272;
  wire[13:0] T273;
  wire[12:0] T274;
  wire[12:0] T275;
  wire[11:0] T276;
  wire[11:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire[9:0] T280;
  wire[9:0] T281;
  wire[8:0] T282;
  wire[8:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[6:0] T286;
  wire[6:0] T287;
  wire[5:0] T288;
  wire[5:0] T289;
  wire[4:0] T290;
  wire[4:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire[1:0] T296;
  wire[1:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire[1:0] T301;
  wire[1:0] T302;
  wire[1:0] T303;
  wire[2:0] T304;
  wire[2:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire[1:0] T309;
  wire[1:0] T310;
  wire[1:0] T311;
  wire[2:0] T312;
  wire[2:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire[1:0] T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire[2:0] T320;
  wire[2:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire[1:0] T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire[2:0] T328;
  wire[2:0] T329;
  wire T330;
  wire T331;
  wire T332;
  wire[1:0] T333;
  wire[1:0] T334;
  wire[1:0] T335;
  wire[2:0] T336;
  wire[2:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire[1:0] T341;
  wire[1:0] T342;
  wire[1:0] T343;
  wire[2:0] T344;
  wire[2:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire[1:0] T352;
  wire[1:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire[1:0] T360;
  wire[1:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[1:0] T368;
  wire[1:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire[1:0] T384;
  wire[1:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire[1:0] T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire[1:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[1:0] T408;
  wire[1:0] T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire[1:0] T416;
  wire[1:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire[1:0] T421;
  wire[1:0] T422;
  wire[1:0] T423;
  wire[2:0] T424;
  wire[2:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire[1:0] T429;
  wire[1:0] T430;
  wire[1:0] T431;
  wire[2:0] T432;
  wire[2:0] T433;
  wire T434;
  wire T435;
  wire T436;
  wire[1:0] T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire[2:0] T440;
  wire[2:0] T441;
  wire T442;
  wire T443;
  wire T444;
  wire[1:0] T445;
  wire[1:0] T446;
  wire[1:0] T447;
  wire[2:0] T448;
  wire[2:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire[1:0] T453;
  wire[1:0] T454;
  wire[1:0] T455;
  wire[2:0] T456;
  wire[2:0] T457;
  wire T458;
  wire T459;
  wire T460;
  wire[1:0] T461;
  wire[1:0] T462;
  wire[1:0] T463;
  wire[2:0] T464;
  wire[2:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire[1:0] T480;
  wire[1:0] T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[1:0] T488;
  wire[1:0] T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire[1:0] T496;
  wire[1:0] T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire[1:0] T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire[1:0] T512;
  wire[1:0] T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire[1:0] T520;
  wire[1:0] T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire[1:0] T528;
  wire[1:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[1:0] T536;
  wire[1:0] T537;
  wire T538;
  wire T539;
  wire T540;
  wire[1:0] T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire[2:0] T544;
  wire[2:0] T545;
  wire T546;
  wire T547;
  wire T548;
  wire[1:0] T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire[2:0] T552;
  wire[2:0] T553;
  wire T554;
  wire T555;
  wire T556;
  wire[1:0] T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire[2:0] T560;
  wire[2:0] T561;
  wire T562;
  wire T563;
  wire T564;
  wire[1:0] T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire[2:0] T568;
  wire[2:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire[1:0] T573;
  wire[1:0] T574;
  wire[1:0] T575;
  wire[2:0] T576;
  wire[2:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire[1:0] T581;
  wire[1:0] T582;
  wire[1:0] T583;
  wire[2:0] T584;
  wire[2:0] T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[1:0] T592;
  wire[1:0] T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire[1:0] T600;
  wire[1:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire[1:0] T608;
  wire[1:0] T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire[1:0] T616;
  wire[1:0] T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[1:0] T624;
  wire[1:0] T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[1:0] T632;
  wire[1:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire[1:0] T640;
  wire[1:0] T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire[1:0] T648;
  wire[1:0] T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire[1:0] T656;
  wire[1:0] T657;
  wire T658;
  wire T659;
  wire T660;
  wire[3:0] T661;
  wire[3:0] T662;
  wire[3:0] T663;
  wire[10:0] T664;
  wire[10:0] T665;
  wire T666;
  wire T667;
  wire T668;
  wire[1:0] T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire[2:0] T672;
  wire[2:0] T673;
  wire T674;
  wire T675;
  wire T676;
  wire[3:0] T677;
  wire[3:0] T678;
  wire[3:0] T679;
  wire[10:0] T680;
  wire[10:0] T681;
  wire T682;
  wire T683;
  wire T684;
  wire[1:0] T685;
  wire[1:0] T686;
  wire[1:0] T687;
  wire[2:0] T688;
  wire[2:0] T689;
  wire T690;
  wire T691;
  wire T692;
  wire[3:0] T693;
  wire[3:0] T694;
  wire[3:0] T695;
  wire[10:0] T696;
  wire[10:0] T697;
  wire T698;
  wire T699;
  wire T700;
  wire[1:0] T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire[2:0] T704;
  wire[2:0] T705;
  wire T706;
  wire T707;
  wire T708;
  wire[3:0] T709;
  wire[3:0] T710;
  wire[3:0] T711;
  wire[10:0] T712;
  wire[10:0] T713;
  wire T714;
  wire T715;
  wire T716;
  wire[1:0] T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire[2:0] T720;
  wire[2:0] T721;
  wire T722;
  wire T723;
  wire T724;
  wire[3:0] T725;
  wire[3:0] T726;
  wire[3:0] T727;
  wire[10:0] T728;
  wire[10:0] T729;
  wire T730;
  wire T731;
  wire T732;
  wire[1:0] T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire[2:0] T736;
  wire[2:0] T737;
  wire T738;
  wire T739;
  wire T740;
  wire[3:0] T741;
  wire[3:0] T742;
  wire[3:0] T743;
  wire[10:0] T744;
  wire[10:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire[1:0] T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire[2:0] T752;
  wire[2:0] T753;
  wire T754;
  wire T755;
  wire T756;
  wire[3:0] T757;
  wire[3:0] T758;
  wire[3:0] T759;
  wire[10:0] T760;
  wire[10:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire[1:0] T768;
  wire[1:0] T769;
  wire T770;
  wire T771;
  wire T772;
  wire[3:0] T773;
  wire[3:0] T774;
  wire[3:0] T775;
  wire[10:0] T776;
  wire[10:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[1:0] T784;
  wire[1:0] T785;
  wire T786;
  wire T787;
  wire T788;
  wire[3:0] T789;
  wire[3:0] T790;
  wire[3:0] T791;
  wire[10:0] T792;
  wire[10:0] T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire[1:0] T800;
  wire[1:0] T801;
  wire T802;
  wire T803;
  wire T804;
  wire[3:0] T805;
  wire[3:0] T806;
  wire[3:0] T807;
  wire[9:0] T808;
  wire[9:0] T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire[1:0] T816;
  wire[1:0] T817;
  wire T818;
  wire T819;
  wire T820;
  wire[3:0] T821;
  wire[3:0] T822;
  wire[3:0] T823;
  wire[9:0] T824;
  wire[9:0] T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire[1:0] T832;
  wire[1:0] T833;
  wire T834;
  wire T835;
  wire T836;
  wire[3:0] T837;
  wire[3:0] T838;
  wire[3:0] T839;
  wire[9:0] T840;
  wire[9:0] T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire T847;
  wire[1:0] T848;
  wire[1:0] T849;
  wire T850;
  wire T851;
  wire T852;
  wire[3:0] T853;
  wire[3:0] T854;
  wire[3:0] T855;
  wire[9:0] T856;
  wire[9:0] T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire[1:0] T864;
  wire[1:0] T865;
  wire T866;
  wire T867;
  wire T868;
  wire[3:0] T869;
  wire[3:0] T870;
  wire[3:0] T871;
  wire[9:0] T872;
  wire[9:0] T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire[1:0] T880;
  wire[1:0] T881;
  wire T882;
  wire T883;
  wire T884;
  wire[3:0] T885;
  wire[3:0] T886;
  wire[3:0] T887;
  wire[9:0] T888;
  wire[9:0] T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire[1:0] T896;
  wire[1:0] T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire[1:0] T904;
  wire[1:0] T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire[1:0] T912;
  wire[1:0] T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire[1:0] T920;
  wire[1:0] T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire[1:0] T928;
  wire[1:0] T929;
  wire T930;
  wire T931;
  wire T932;
  wire[3:0] T933;
  wire[3:0] T934;
  wire[3:0] T935;
  wire[8:0] T936;
  wire[8:0] T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire[1:0] T944;
  wire[1:0] T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire[1:0] T952;
  wire[1:0] T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire[1:0] T960;
  wire[1:0] T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire T966;
  wire T967;
  wire[1:0] T968;
  wire[1:0] T969;
  wire T970;
  wire T971;
  wire T972;
  wire[3:0] T973;
  wire[3:0] T974;
  wire[3:0] T975;
  wire[8:0] T976;
  wire[8:0] T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire[1:0] T984;
  wire[1:0] T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire[1:0] T992;
  wire[1:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[1:0] T1000;
  wire[1:0] T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire T1006;
  wire T1007;
  wire[1:0] T1008;
  wire[1:0] T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire[3:0] T1013;
  wire[3:0] T1014;
  wire[3:0] T1015;
  wire[8:0] T1016;
  wire[8:0] T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[1:0] T1024;
  wire[1:0] T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire[1:0] T1032;
  wire[1:0] T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire[1:0] T1040;
  wire[1:0] T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  wire[1:0] T1048;
  wire[1:0] T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire[3:0] T1053;
  wire[3:0] T1054;
  wire[3:0] T1055;
  wire[8:0] T1056;
  wire[8:0] T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[1:0] T1064;
  wire[1:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire[1:0] T1072;
  wire[1:0] T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire T1078;
  wire T1079;
  wire[1:0] T1080;
  wire[1:0] T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire[1:0] T1088;
  wire[1:0] T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire[3:0] T1093;
  wire[3:0] T1094;
  wire[3:0] T1095;
  wire[8:0] T1096;
  wire[8:0] T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire[1:0] T1104;
  wire[1:0] T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire[1:0] T1112;
  wire[1:0] T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire[1:0] T1120;
  wire[1:0] T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire T1127;
  wire[1:0] T1128;
  wire[1:0] T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire[3:0] T1133;
  wire[3:0] T1134;
  wire[3:0] T1135;
  wire[8:0] T1136;
  wire[8:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[1:0] T1144;
  wire[1:0] T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire[1:0] T1152;
  wire[1:0] T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire[1:0] T1160;
  wire[1:0] T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire[1:0] T1168;
  wire[1:0] T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire[3:0] T1173;
  wire[3:0] T1174;
  wire[3:0] T1175;
  wire[8:0] T1176;
  wire[8:0] T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire[1:0] T1184;
  wire[1:0] T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire[1:0] T1192;
  wire[1:0] T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire[1:0] T1200;
  wire[1:0] T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[1:0] T1208;
  wire[1:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire[3:0] T1213;
  wire[3:0] T1214;
  wire[3:0] T1215;
  wire[8:0] T1216;
  wire[8:0] T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire[1:0] T1224;
  wire[1:0] T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire[1:0] T1232;
  wire[1:0] T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire[1:0] T1240;
  wire[1:0] T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire[1:0] T1248;
  wire[1:0] T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire[3:0] T1253;
  wire[3:0] T1254;
  wire[3:0] T1255;
  wire[8:0] T1256;
  wire[8:0] T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire[1:0] T1264;
  wire[1:0] T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire[1:0] T1272;
  wire[1:0] T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire T1277;
  wire T1278;
  wire T1279;
  wire[1:0] T1280;
  wire[1:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[1:0] T1288;
  wire[1:0] T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire[3:0] T1293;
  wire[3:0] T1294;
  wire[3:0] T1295;
  wire[8:0] T1296;
  wire[8:0] T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire[1:0] T1304;
  wire[1:0] T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire[1:0] T1312;
  wire[1:0] T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire[1:0] T1320;
  wire[1:0] T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire[1:0] T1328;
  wire[1:0] T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire[3:0] T1333;
  wire[3:0] T1334;
  wire[3:0] T1335;
  wire[8:0] T1336;
  wire[8:0] T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire T1343;
  wire[1:0] T1344;
  wire[1:0] T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[1:0] T1352;
  wire[1:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire T1357;
  wire T1358;
  wire T1359;
  wire[1:0] T1360;
  wire[1:0] T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  wire T1366;
  wire T1367;
  wire[1:0] T1368;
  wire[1:0] T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire[3:0] T1373;
  wire[3:0] T1374;
  wire[3:0] T1375;
  wire[8:0] T1376;
  wire[8:0] T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire[1:0] T1384;
  wire[1:0] T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire[1:0] T1392;
  wire[1:0] T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[1:0] T1400;
  wire[1:0] T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire[1:0] T1408;
  wire[1:0] T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire[3:0] T1413;
  wire[3:0] T1414;
  wire[3:0] T1415;
  wire[8:0] T1416;
  wire[8:0] T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire T1421;
  wire T1422;
  wire T1423;
  wire[1:0] T1424;
  wire[1:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[1:0] T1432;
  wire[1:0] T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire T1437;
  wire T1438;
  wire T1439;
  wire[1:0] T1440;
  wire[1:0] T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire[1:0] T1448;
  wire[1:0] T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire[3:0] T1453;
  wire[3:0] T1454;
  wire[3:0] T1455;
  wire[8:0] T1456;
  wire[8:0] T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire[1:0] T1464;
  wire[1:0] T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire[1:0] T1472;
  wire[1:0] T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire T1478;
  wire T1479;
  wire[1:0] T1480;
  wire[1:0] T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire T1485;
  wire T1486;
  wire T1487;
  wire[1:0] T1488;
  wire[1:0] T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire[3:0] T1493;
  wire[3:0] T1494;
  wire[3:0] T1495;
  wire[8:0] T1496;
  wire[8:0] T1497;
  wire[22:0] T1498;
  wire[22:0] T1499;
  wire[21:0] T1500;
  wire[21:0] T1501;
  wire[20:0] T1502;
  wire[20:0] T1503;
  wire[19:0] T1504;
  wire[19:0] T1505;
  wire[18:0] T1506;
  wire[18:0] T1507;
  wire[17:0] T1508;
  wire[17:0] T1509;
  wire[16:0] T1510;
  wire[16:0] T1511;
  wire[15:0] T1512;
  wire[15:0] T1513;
  wire[14:0] T1514;
  wire[14:0] T1515;
  wire[13:0] T1516;
  wire[13:0] T1517;
  wire[12:0] T1518;
  wire[12:0] T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[10:0] T1522;
  wire[10:0] T1523;
  wire[9:0] T1524;
  wire[9:0] T1525;
  wire[8:0] T1526;
  wire[8:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[6:0] T1530;
  wire[6:0] T1531;
  wire[5:0] T1532;
  wire[5:0] T1533;
  wire[4:0] T1534;
  wire[4:0] T1535;
  wire[3:0] T1536;
  wire[3:0] T1537;
  wire[2:0] T1538;
  wire[2:0] T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[11:0] T1660;
  wire[11:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[11:0] T1668;
  wire[11:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[11:0] T1676;
  wire[11:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[11:0] T1684;
  wire[11:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[11:0] T1692;
  wire[11:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[11:0] T1700;
  wire[11:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[11:0] T1708;
  wire[11:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[11:0] T1716;
  wire[11:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[11:0] T1724;
  wire[11:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1490, T2};
  assign T2 = T3;
  assign T3 = {T1482, T4};
  assign T4 = T5;
  assign T5 = {T1474, T6};
  assign T6 = T7;
  assign T7 = {T1466, T8};
  assign T8 = T9;
  assign T9 = {T1458, T10};
  assign T10 = T11;
  assign T11 = {T1450, T12};
  assign T12 = T13;
  assign T13 = {T1442, T14};
  assign T14 = T15;
  assign T15 = {T1434, T16};
  assign T16 = T17;
  assign T17 = {T1426, T18};
  assign T18 = T19;
  assign T19 = {T1418, T20};
  assign T20 = T21;
  assign T21 = {T1410, T22};
  assign T22 = T23;
  assign T23 = {T1402, T24};
  assign T24 = T25;
  assign T25 = {T1394, T26};
  assign T26 = T27;
  assign T27 = {T1386, T28};
  assign T28 = T29;
  assign T29 = {T1378, T30};
  assign T30 = T31;
  assign T31 = {T1370, T32};
  assign T32 = T33;
  assign T33 = {T1362, T34};
  assign T34 = T35;
  assign T35 = {T1354, T36};
  assign T36 = T37;
  assign T37 = {T1346, T38};
  assign T38 = T39;
  assign T39 = {T1338, T40};
  assign T40 = T41;
  assign T41 = {T1330, T42};
  assign T42 = T43;
  assign T43 = {T1322, T44};
  assign T44 = T45;
  assign T45 = {T1314, T46};
  assign T46 = T47;
  assign T47 = {T1306, T48};
  assign T48 = T49;
  assign T49 = {T1298, T50};
  assign T50 = T51;
  assign T51 = {T1290, T52};
  assign T52 = T53;
  assign T53 = {T1282, T54};
  assign T54 = T55;
  assign T55 = {T1274, T56};
  assign T56 = T57;
  assign T57 = {T1266, T58};
  assign T58 = T59;
  assign T59 = {T1258, T60};
  assign T60 = T61;
  assign T61 = {T1250, T62};
  assign T62 = T63;
  assign T63 = {T1242, T64};
  assign T64 = T65;
  assign T65 = {T1234, T66};
  assign T66 = T67;
  assign T67 = {T1226, T68};
  assign T68 = T69;
  assign T69 = {T1218, T70};
  assign T70 = T71;
  assign T71 = {T1210, T72};
  assign T72 = T73;
  assign T73 = {T1202, T74};
  assign T74 = T75;
  assign T75 = {T1194, T76};
  assign T76 = T77;
  assign T77 = {T1186, T78};
  assign T78 = T79;
  assign T79 = {T1178, T80};
  assign T80 = T81;
  assign T81 = {T1170, T82};
  assign T82 = T83;
  assign T83 = {T1162, T84};
  assign T84 = T85;
  assign T85 = {T1154, T86};
  assign T86 = T87;
  assign T87 = {T1146, T88};
  assign T88 = T89;
  assign T89 = {T1138, T90};
  assign T90 = T91;
  assign T91 = {T1130, T92};
  assign T92 = T93;
  assign T93 = {T1122, T94};
  assign T94 = T95;
  assign T95 = {T1114, T96};
  assign T96 = T97;
  assign T97 = {T1106, T98};
  assign T98 = T99;
  assign T99 = {T1098, T100};
  assign T100 = T101;
  assign T101 = {T1090, T102};
  assign T102 = T103;
  assign T103 = {T1082, T104};
  assign T104 = T105;
  assign T105 = {T1074, T106};
  assign T106 = T107;
  assign T107 = {T1066, T108};
  assign T108 = T109;
  assign T109 = {T1058, T110};
  assign T110 = T111;
  assign T111 = {T1050, T112};
  assign T112 = T113;
  assign T113 = {T1042, T114};
  assign T114 = T115;
  assign T115 = {T1034, T116};
  assign T116 = T117;
  assign T117 = {T1026, T118};
  assign T118 = T119;
  assign T119 = {T1018, T120};
  assign T120 = T121;
  assign T121 = {T1010, T122};
  assign T122 = T123;
  assign T123 = {T1002, T124};
  assign T124 = T125;
  assign T125 = {T994, T126};
  assign T126 = T127;
  assign T127 = {T986, T128};
  assign T128 = T129;
  assign T129 = {T978, T130};
  assign T130 = T131;
  assign T131 = {T970, T132};
  assign T132 = T133;
  assign T133 = {T962, T134};
  assign T134 = T135;
  assign T135 = {T954, T136};
  assign T136 = T137;
  assign T137 = {T946, T138};
  assign T138 = T139;
  assign T139 = {T938, T140};
  assign T140 = T141;
  assign T141 = {T930, T142};
  assign T142 = T143;
  assign T143 = {T922, T144};
  assign T144 = T145;
  assign T145 = {T914, T146};
  assign T146 = T147;
  assign T147 = {T906, T148};
  assign T148 = T149;
  assign T149 = {T898, T150};
  assign T150 = T151;
  assign T151 = {T890, T152};
  assign T152 = T153;
  assign T153 = {T882, T154};
  assign T154 = T155;
  assign T155 = {T874, T156};
  assign T156 = T157;
  assign T157 = {T866, T158};
  assign T158 = T159;
  assign T159 = {T858, T160};
  assign T160 = T161;
  assign T161 = {T850, T162};
  assign T162 = T163;
  assign T163 = {T842, T164};
  assign T164 = T165;
  assign T165 = {T834, T166};
  assign T166 = T167;
  assign T167 = {T826, T168};
  assign T168 = T169;
  assign T169 = {T818, T170};
  assign T170 = T171;
  assign T171 = {T810, T172};
  assign T172 = T173;
  assign T173 = {T802, T174};
  assign T174 = T175;
  assign T175 = {T794, T176};
  assign T176 = T177;
  assign T177 = {T786, T178};
  assign T178 = T179;
  assign T179 = {T778, T180};
  assign T180 = T181;
  assign T181 = {T770, T182};
  assign T182 = T183;
  assign T183 = {T762, T184};
  assign T184 = T185;
  assign T185 = {T754, T186};
  assign T186 = T187;
  assign T187 = {T746, T188};
  assign T188 = T189;
  assign T189 = {T738, T190};
  assign T190 = T191;
  assign T191 = {T730, T192};
  assign T192 = T193;
  assign T193 = {T722, T194};
  assign T194 = T195;
  assign T195 = {T714, T196};
  assign T196 = T197;
  assign T197 = {T706, T198};
  assign T198 = T199;
  assign T199 = {T698, T200};
  assign T200 = T201;
  assign T201 = {T690, T202};
  assign T202 = T203;
  assign T203 = {T682, T204};
  assign T204 = T205;
  assign T205 = {T674, T206};
  assign T206 = T207;
  assign T207 = {T666, T208};
  assign T208 = T209;
  assign T209 = {T658, T210};
  assign T210 = T211;
  assign T211 = {T650, T212};
  assign T212 = T213;
  assign T213 = {T642, T214};
  assign T214 = T215;
  assign T215 = {T634, T216};
  assign T216 = T217;
  assign T217 = {T626, T218};
  assign T218 = T219;
  assign T219 = {T618, T220};
  assign T220 = T221;
  assign T221 = {T610, T222};
  assign T222 = T223;
  assign T223 = {T602, T224};
  assign T224 = T225;
  assign T225 = {T594, T226};
  assign T226 = T227;
  assign T227 = {T586, T228};
  assign T228 = T229;
  assign T229 = {T578, T230};
  assign T230 = T231;
  assign T231 = {T570, T232};
  assign T232 = T233;
  assign T233 = {T562, T234};
  assign T234 = T235;
  assign T235 = {T554, T236};
  assign T236 = T237;
  assign T237 = {T546, T238};
  assign T238 = T239;
  assign T239 = {T538, T240};
  assign T240 = T241;
  assign T241 = {T530, T242};
  assign T242 = T243;
  assign T243 = {T522, T244};
  assign T244 = T245;
  assign T245 = {T514, T246};
  assign T246 = T247;
  assign T247 = {T506, T248};
  assign T248 = T249;
  assign T249 = {T498, T250};
  assign T250 = T251;
  assign T251 = {T490, T252};
  assign T252 = T253;
  assign T253 = {T482, T254};
  assign T254 = T255;
  assign T255 = {T474, T256};
  assign T256 = T257;
  assign T257 = {T466, T258};
  assign T258 = T259;
  assign T259 = {T458, T260};
  assign T260 = T261;
  assign T261 = {T450, T262};
  assign T262 = T263;
  assign T263 = {T442, T264};
  assign T264 = T265;
  assign T265 = {T434, T266};
  assign T266 = T267;
  assign T267 = {T426, T268};
  assign T268 = T269;
  assign T269 = {T418, T270};
  assign T270 = T271;
  assign T271 = {T410, T272};
  assign T272 = T273;
  assign T273 = {T402, T274};
  assign T274 = T275;
  assign T275 = {T394, T276};
  assign T276 = T277;
  assign T277 = {T386, T278};
  assign T278 = T279;
  assign T279 = {T378, T280};
  assign T280 = T281;
  assign T281 = {T370, T282};
  assign T282 = T283;
  assign T283 = {T362, T284};
  assign T284 = T285;
  assign T285 = {T354, T286};
  assign T286 = T287;
  assign T287 = {T346, T288};
  assign T288 = T289;
  assign T289 = {T338, T290};
  assign T290 = T291;
  assign T291 = {T330, T292};
  assign T292 = T293;
  assign T293 = {T322, T294};
  assign T294 = T295;
  assign T295 = {T314, T296};
  assign T296 = T297;
  assign T297 = {T306, T298};
  assign T298 = T299;
  assign T299 = T300;
  assign T300 = T304[T301];
  assign T301 = T302;
  assign T302 = T303;
  assign T303 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T304 = T305;
  assign T305 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T306 = T307;
  assign T307 = T308;
  assign T308 = T312[T309];
  assign T309 = T310;
  assign T310 = T311;
  assign T311 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T312 = T313;
  assign T313 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T314 = T315;
  assign T315 = T316;
  assign T316 = T320[T317];
  assign T317 = T318;
  assign T318 = T319;
  assign T319 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T320 = T321;
  assign T321 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T322 = T323;
  assign T323 = T324;
  assign T324 = T328[T325];
  assign T325 = T326;
  assign T326 = T327;
  assign T327 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T328 = T329;
  assign T329 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T330 = T331;
  assign T331 = T332;
  assign T332 = T336[T333];
  assign T333 = T334;
  assign T334 = T335;
  assign T335 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T336 = T337;
  assign T337 = io_chanxy_in[4'he/* 14*/:4'hc/* 12*/];
  assign T338 = T339;
  assign T339 = T340;
  assign T340 = T344[T341];
  assign T341 = T342;
  assign T342 = T343;
  assign T343 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T344 = T345;
  assign T345 = io_chanxy_in[5'h11/* 17*/:4'hf/* 15*/];
  assign T346 = T347;
  assign T347 = T348;
  assign T348 = T352[T349];
  assign T349 = T350;
  assign T350 = T351;
  assign T351 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T352 = T353;
  assign T353 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T354 = T355;
  assign T355 = T356;
  assign T356 = T360[T357];
  assign T357 = T358;
  assign T358 = T359;
  assign T359 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T360 = T361;
  assign T361 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T362 = T363;
  assign T363 = T364;
  assign T364 = T368[T365];
  assign T365 = T366;
  assign T366 = T367;
  assign T367 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T368 = T369;
  assign T369 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T370 = T371;
  assign T371 = T372;
  assign T372 = T376[T373];
  assign T373 = T374;
  assign T374 = T375;
  assign T375 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T376 = T377;
  assign T377 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T378 = T379;
  assign T379 = T380;
  assign T380 = T384[T381];
  assign T381 = T382;
  assign T382 = T383;
  assign T383 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T384 = T385;
  assign T385 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T386 = T387;
  assign T387 = T388;
  assign T388 = T392[T389];
  assign T389 = T390;
  assign T390 = T391;
  assign T391 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T392 = T393;
  assign T393 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T394 = T395;
  assign T395 = T396;
  assign T396 = T400[T397];
  assign T397 = T398;
  assign T398 = T399;
  assign T399 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T400 = T401;
  assign T401 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T402 = T403;
  assign T403 = T404;
  assign T404 = T408[T405];
  assign T405 = T406;
  assign T406 = T407;
  assign T407 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T408 = T409;
  assign T409 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T410 = T411;
  assign T411 = T412;
  assign T412 = T416[T413];
  assign T413 = T414;
  assign T414 = T415;
  assign T415 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T416 = T417;
  assign T417 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T418 = T419;
  assign T419 = T420;
  assign T420 = T424[T421];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = io_chanxy_config[5'h16/* 22*/:5'h15/* 21*/];
  assign T424 = T425;
  assign T425 = io_chanxy_in[6'h26/* 38*/:6'h24/* 36*/];
  assign T426 = T427;
  assign T427 = T428;
  assign T428 = T432[T429];
  assign T429 = T430;
  assign T430 = T431;
  assign T431 = io_chanxy_config[5'h18/* 24*/:5'h17/* 23*/];
  assign T432 = T433;
  assign T433 = io_chanxy_in[6'h29/* 41*/:6'h27/* 39*/];
  assign T434 = T435;
  assign T435 = T436;
  assign T436 = T440[T437];
  assign T437 = T438;
  assign T438 = T439;
  assign T439 = io_chanxy_config[5'h1a/* 26*/:5'h19/* 25*/];
  assign T440 = T441;
  assign T441 = io_chanxy_in[6'h2c/* 44*/:6'h2a/* 42*/];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = T448[T445];
  assign T445 = T446;
  assign T446 = T447;
  assign T447 = io_chanxy_config[5'h1c/* 28*/:5'h1b/* 27*/];
  assign T448 = T449;
  assign T449 = io_chanxy_in[6'h2f/* 47*/:6'h2d/* 45*/];
  assign T450 = T451;
  assign T451 = T452;
  assign T452 = T456[T453];
  assign T453 = T454;
  assign T454 = T455;
  assign T455 = io_chanxy_config[5'h1e/* 30*/:5'h1d/* 29*/];
  assign T456 = T457;
  assign T457 = io_chanxy_in[6'h32/* 50*/:6'h30/* 48*/];
  assign T458 = T459;
  assign T459 = T460;
  assign T460 = T464[T461];
  assign T461 = T462;
  assign T462 = T463;
  assign T463 = io_chanxy_config[6'h20/* 32*/:5'h1f/* 31*/];
  assign T464 = T465;
  assign T465 = io_chanxy_in[6'h35/* 53*/:6'h33/* 51*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T472[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T472 = T473;
  assign T473 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T474 = T475;
  assign T475 = T476;
  assign T476 = T480[T477];
  assign T477 = T478;
  assign T478 = T479;
  assign T479 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T480 = T481;
  assign T481 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T482 = T483;
  assign T483 = T484;
  assign T484 = T488[T485];
  assign T485 = T486;
  assign T486 = T487;
  assign T487 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T488 = T489;
  assign T489 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T490 = T491;
  assign T491 = T492;
  assign T492 = T496[T493];
  assign T493 = T494;
  assign T494 = T495;
  assign T495 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T496 = T497;
  assign T497 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T498 = T499;
  assign T499 = T500;
  assign T500 = T504[T501];
  assign T501 = T502;
  assign T502 = T503;
  assign T503 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T504 = T505;
  assign T505 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T506 = T507;
  assign T507 = T508;
  assign T508 = T512[T509];
  assign T509 = T510;
  assign T510 = T511;
  assign T511 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T512 = T513;
  assign T513 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T514 = T515;
  assign T515 = T516;
  assign T516 = T520[T517];
  assign T517 = T518;
  assign T518 = T519;
  assign T519 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T520 = T521;
  assign T521 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T522 = T523;
  assign T523 = T524;
  assign T524 = T528[T525];
  assign T525 = T526;
  assign T526 = T527;
  assign T527 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T528 = T529;
  assign T529 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T530 = T531;
  assign T531 = T532;
  assign T532 = T536[T533];
  assign T533 = T534;
  assign T534 = T535;
  assign T535 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T536 = T537;
  assign T537 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T538 = T539;
  assign T539 = T540;
  assign T540 = T544[T541];
  assign T541 = T542;
  assign T542 = T543;
  assign T543 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T544 = T545;
  assign T545 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T546 = T547;
  assign T547 = T548;
  assign T548 = T552[T549];
  assign T549 = T550;
  assign T550 = T551;
  assign T551 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T552 = T553;
  assign T553 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T554 = T555;
  assign T555 = T556;
  assign T556 = T560[T557];
  assign T557 = T558;
  assign T558 = T559;
  assign T559 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T560 = T561;
  assign T561 = io_chanxy_in[7'h50/* 80*/:7'h4e/* 78*/];
  assign T562 = T563;
  assign T563 = T564;
  assign T564 = T568[T565];
  assign T565 = T566;
  assign T566 = T567;
  assign T567 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T568 = T569;
  assign T569 = io_chanxy_in[7'h53/* 83*/:7'h51/* 81*/];
  assign T570 = T571;
  assign T571 = T572;
  assign T572 = T576[T573];
  assign T573 = T574;
  assign T574 = T575;
  assign T575 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T576 = T577;
  assign T577 = io_chanxy_in[7'h56/* 86*/:7'h54/* 84*/];
  assign T578 = T579;
  assign T579 = T580;
  assign T580 = T584[T581];
  assign T581 = T582;
  assign T582 = T583;
  assign T583 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T584 = T585;
  assign T585 = io_chanxy_in[7'h59/* 89*/:7'h57/* 87*/];
  assign T586 = T587;
  assign T587 = T588;
  assign T588 = T592[T589];
  assign T589 = T590;
  assign T590 = T591;
  assign T591 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T592 = T593;
  assign T593 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T594 = T595;
  assign T595 = T596;
  assign T596 = T600[T597];
  assign T597 = T598;
  assign T598 = T599;
  assign T599 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T600 = T601;
  assign T601 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T602 = T603;
  assign T603 = T604;
  assign T604 = T608[T605];
  assign T605 = T606;
  assign T606 = T607;
  assign T607 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T608 = T609;
  assign T609 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T610 = T611;
  assign T611 = T612;
  assign T612 = T616[T613];
  assign T613 = T614;
  assign T614 = T615;
  assign T615 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T616 = T617;
  assign T617 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T618 = T619;
  assign T619 = T620;
  assign T620 = T624[T621];
  assign T621 = T622;
  assign T622 = T623;
  assign T623 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T624 = T625;
  assign T625 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T626 = T627;
  assign T627 = T628;
  assign T628 = T632[T629];
  assign T629 = T630;
  assign T630 = T631;
  assign T631 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T632 = T633;
  assign T633 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T634 = T635;
  assign T635 = T636;
  assign T636 = T640[T637];
  assign T637 = T638;
  assign T638 = T639;
  assign T639 = io_chanxy_config[6'h3c/* 60*/:6'h3c/* 60*/];
  assign T640 = T641;
  assign T641 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T642 = T643;
  assign T643 = T644;
  assign T644 = T648[T645];
  assign T645 = T646;
  assign T646 = T647;
  assign T647 = io_chanxy_config[6'h3d/* 61*/:6'h3d/* 61*/];
  assign T648 = T649;
  assign T649 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T650 = T651;
  assign T651 = T652;
  assign T652 = T656[T653];
  assign T653 = T654;
  assign T654 = T655;
  assign T655 = io_chanxy_config[6'h3e/* 62*/:6'h3e/* 62*/];
  assign T656 = T657;
  assign T657 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T658 = T659;
  assign T659 = T660;
  assign T660 = T664[T661];
  assign T661 = T662;
  assign T662 = T663;
  assign T663 = io_chanxy_config[7'h42/* 66*/:6'h3f/* 63*/];
  assign T664 = T665;
  assign T665 = io_chanxy_in[7'h76/* 118*/:7'h6c/* 108*/];
  assign T666 = T667;
  assign T667 = T668;
  assign T668 = T672[T669];
  assign T669 = T670;
  assign T670 = T671;
  assign T671 = io_chanxy_config[7'h44/* 68*/:7'h43/* 67*/];
  assign T672 = T673;
  assign T673 = io_chanxy_in[7'h79/* 121*/:7'h77/* 119*/];
  assign T674 = T675;
  assign T675 = T676;
  assign T676 = T680[T677];
  assign T677 = T678;
  assign T678 = T679;
  assign T679 = io_chanxy_config[7'h48/* 72*/:7'h45/* 69*/];
  assign T680 = T681;
  assign T681 = io_chanxy_in[8'h84/* 132*/:7'h7a/* 122*/];
  assign T682 = T683;
  assign T683 = T684;
  assign T684 = T688[T685];
  assign T685 = T686;
  assign T686 = T687;
  assign T687 = io_chanxy_config[7'h4a/* 74*/:7'h49/* 73*/];
  assign T688 = T689;
  assign T689 = io_chanxy_in[8'h87/* 135*/:8'h85/* 133*/];
  assign T690 = T691;
  assign T691 = T692;
  assign T692 = T696[T693];
  assign T693 = T694;
  assign T694 = T695;
  assign T695 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T696 = T697;
  assign T697 = io_chanxy_in[8'h92/* 146*/:8'h88/* 136*/];
  assign T698 = T699;
  assign T699 = T700;
  assign T700 = T704[T701];
  assign T701 = T702;
  assign T702 = T703;
  assign T703 = io_chanxy_config[7'h50/* 80*/:7'h4f/* 79*/];
  assign T704 = T705;
  assign T705 = io_chanxy_in[8'h95/* 149*/:8'h93/* 147*/];
  assign T706 = T707;
  assign T707 = T708;
  assign T708 = T712[T709];
  assign T709 = T710;
  assign T710 = T711;
  assign T711 = io_chanxy_config[7'h54/* 84*/:7'h51/* 81*/];
  assign T712 = T713;
  assign T713 = io_chanxy_in[8'ha0/* 160*/:8'h96/* 150*/];
  assign T714 = T715;
  assign T715 = T716;
  assign T716 = T720[T717];
  assign T717 = T718;
  assign T718 = T719;
  assign T719 = io_chanxy_config[7'h56/* 86*/:7'h55/* 85*/];
  assign T720 = T721;
  assign T721 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T722 = T723;
  assign T723 = T724;
  assign T724 = T728[T725];
  assign T725 = T726;
  assign T726 = T727;
  assign T727 = io_chanxy_config[7'h5a/* 90*/:7'h57/* 87*/];
  assign T728 = T729;
  assign T729 = io_chanxy_in[8'hae/* 174*/:8'ha4/* 164*/];
  assign T730 = T731;
  assign T731 = T732;
  assign T732 = T736[T733];
  assign T733 = T734;
  assign T734 = T735;
  assign T735 = io_chanxy_config[7'h5c/* 92*/:7'h5b/* 91*/];
  assign T736 = T737;
  assign T737 = io_chanxy_in[8'hb1/* 177*/:8'haf/* 175*/];
  assign T738 = T739;
  assign T739 = T740;
  assign T740 = T744[T741];
  assign T741 = T742;
  assign T742 = T743;
  assign T743 = io_chanxy_config[7'h60/* 96*/:7'h5d/* 93*/];
  assign T744 = T745;
  assign T745 = io_chanxy_in[8'hbc/* 188*/:8'hb2/* 178*/];
  assign T746 = T747;
  assign T747 = T748;
  assign T748 = T752[T749];
  assign T749 = T750;
  assign T750 = T751;
  assign T751 = io_chanxy_config[7'h62/* 98*/:7'h61/* 97*/];
  assign T752 = T753;
  assign T753 = io_chanxy_in[8'hbf/* 191*/:8'hbd/* 189*/];
  assign T754 = T755;
  assign T755 = T756;
  assign T756 = T760[T757];
  assign T757 = T758;
  assign T758 = T759;
  assign T759 = io_chanxy_config[7'h66/* 102*/:7'h63/* 99*/];
  assign T760 = T761;
  assign T761 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T762 = T763;
  assign T763 = T764;
  assign T764 = T768[T765];
  assign T765 = T766;
  assign T766 = T767;
  assign T767 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T768 = T769;
  assign T769 = io_chanxy_in[8'hcc/* 204*/:8'hcb/* 203*/];
  assign T770 = T771;
  assign T771 = T772;
  assign T772 = T776[T773];
  assign T773 = T774;
  assign T774 = T775;
  assign T775 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T776 = T777;
  assign T777 = io_chanxy_in[8'hd7/* 215*/:8'hcd/* 205*/];
  assign T778 = T779;
  assign T779 = T780;
  assign T780 = T784[T781];
  assign T781 = T782;
  assign T782 = T783;
  assign T783 = io_chanxy_config[7'h6c/* 108*/:7'h6c/* 108*/];
  assign T784 = T785;
  assign T785 = io_chanxy_in[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T786 = T787;
  assign T787 = T788;
  assign T788 = T792[T789];
  assign T789 = T790;
  assign T790 = T791;
  assign T791 = io_chanxy_config[7'h70/* 112*/:7'h6d/* 109*/];
  assign T792 = T793;
  assign T793 = io_chanxy_in[8'he4/* 228*/:8'hda/* 218*/];
  assign T794 = T795;
  assign T795 = T796;
  assign T796 = T800[T797];
  assign T797 = T798;
  assign T798 = T799;
  assign T799 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T800 = T801;
  assign T801 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T802 = T803;
  assign T803 = T804;
  assign T804 = T808[T805];
  assign T805 = T806;
  assign T806 = T807;
  assign T807 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T808 = T809;
  assign T809 = io_chanxy_in[8'hf0/* 240*/:8'he7/* 231*/];
  assign T810 = T811;
  assign T811 = T812;
  assign T812 = T816[T813];
  assign T813 = T814;
  assign T814 = T815;
  assign T815 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T816 = T817;
  assign T817 = io_chanxy_in[8'hf2/* 242*/:8'hf1/* 241*/];
  assign T818 = T819;
  assign T819 = T820;
  assign T820 = T824[T821];
  assign T821 = T822;
  assign T822 = T823;
  assign T823 = io_chanxy_config[7'h7a/* 122*/:7'h77/* 119*/];
  assign T824 = T825;
  assign T825 = io_chanxy_in[8'hfc/* 252*/:8'hf3/* 243*/];
  assign T826 = T827;
  assign T827 = T828;
  assign T828 = T832[T829];
  assign T829 = T830;
  assign T830 = T831;
  assign T831 = io_chanxy_config[7'h7b/* 123*/:7'h7b/* 123*/];
  assign T832 = T833;
  assign T833 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T834 = T835;
  assign T835 = T836;
  assign T836 = T840[T837];
  assign T837 = T838;
  assign T838 = T839;
  assign T839 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T840 = T841;
  assign T841 = io_chanxy_in[9'h108/* 264*/:8'hff/* 255*/];
  assign T842 = T843;
  assign T843 = T844;
  assign T844 = T848[T845];
  assign T845 = T846;
  assign T846 = T847;
  assign T847 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T848 = T849;
  assign T849 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T850 = T851;
  assign T851 = T852;
  assign T852 = T856[T853];
  assign T853 = T854;
  assign T854 = T855;
  assign T855 = io_chanxy_config[8'h84/* 132*/:8'h81/* 129*/];
  assign T856 = T857;
  assign T857 = io_chanxy_in[9'h114/* 276*/:9'h10b/* 267*/];
  assign T858 = T859;
  assign T859 = T860;
  assign T860 = T864[T861];
  assign T861 = T862;
  assign T862 = T863;
  assign T863 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T864 = T865;
  assign T865 = io_chanxy_in[9'h116/* 278*/:9'h115/* 277*/];
  assign T866 = T867;
  assign T867 = T868;
  assign T868 = T872[T869];
  assign T869 = T870;
  assign T870 = T871;
  assign T871 = io_chanxy_config[8'h89/* 137*/:8'h86/* 134*/];
  assign T872 = T873;
  assign T873 = io_chanxy_in[9'h120/* 288*/:9'h117/* 279*/];
  assign T874 = T875;
  assign T875 = T876;
  assign T876 = T880[T877];
  assign T877 = T878;
  assign T878 = T879;
  assign T879 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T880 = T881;
  assign T881 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T882 = T883;
  assign T883 = T884;
  assign T884 = T888[T885];
  assign T885 = T886;
  assign T886 = T887;
  assign T887 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T888 = T889;
  assign T889 = io_chanxy_in[9'h12c/* 300*/:9'h123/* 291*/];
  assign T890 = T891;
  assign T891 = T892;
  assign T892 = T896[T893];
  assign T893 = T894;
  assign T894 = T895;
  assign T895 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T896 = T897;
  assign T897 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T898 = T899;
  assign T899 = T900;
  assign T900 = T904[T901];
  assign T901 = T902;
  assign T902 = T903;
  assign T903 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T904 = T905;
  assign T905 = io_chanxy_in[9'h130/* 304*/:9'h12f/* 303*/];
  assign T906 = T907;
  assign T907 = T908;
  assign T908 = T912[T909];
  assign T909 = T910;
  assign T910 = T911;
  assign T911 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T912 = T913;
  assign T913 = io_chanxy_in[9'h132/* 306*/:9'h131/* 305*/];
  assign T914 = T915;
  assign T915 = T916;
  assign T916 = T920[T917];
  assign T917 = T918;
  assign T918 = T919;
  assign T919 = io_chanxy_config[8'h92/* 146*/:8'h92/* 146*/];
  assign T920 = T921;
  assign T921 = io_chanxy_in[9'h134/* 308*/:9'h133/* 307*/];
  assign T922 = T923;
  assign T923 = T924;
  assign T924 = T928[T925];
  assign T925 = T926;
  assign T926 = T927;
  assign T927 = io_chanxy_config[8'h93/* 147*/:8'h93/* 147*/];
  assign T928 = T929;
  assign T929 = io_chanxy_in[9'h136/* 310*/:9'h135/* 309*/];
  assign T930 = T931;
  assign T931 = T932;
  assign T932 = T936[T933];
  assign T933 = T934;
  assign T934 = T935;
  assign T935 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T936 = T937;
  assign T937 = io_chanxy_in[9'h13f/* 319*/:9'h137/* 311*/];
  assign T938 = T939;
  assign T939 = T940;
  assign T940 = T944[T941];
  assign T941 = T942;
  assign T942 = T943;
  assign T943 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T944 = T945;
  assign T945 = io_chanxy_in[9'h141/* 321*/:9'h140/* 320*/];
  assign T946 = T947;
  assign T947 = T948;
  assign T948 = T952[T949];
  assign T949 = T950;
  assign T950 = T951;
  assign T951 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T952 = T953;
  assign T953 = io_chanxy_in[9'h143/* 323*/:9'h142/* 322*/];
  assign T954 = T955;
  assign T955 = T956;
  assign T956 = T960[T957];
  assign T957 = T958;
  assign T958 = T959;
  assign T959 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T960 = T961;
  assign T961 = io_chanxy_in[9'h145/* 325*/:9'h144/* 324*/];
  assign T962 = T963;
  assign T963 = T964;
  assign T964 = T968[T965];
  assign T965 = T966;
  assign T966 = T967;
  assign T967 = io_chanxy_config[8'h9b/* 155*/:8'h9b/* 155*/];
  assign T968 = T969;
  assign T969 = io_chanxy_in[9'h147/* 327*/:9'h146/* 326*/];
  assign T970 = T971;
  assign T971 = T972;
  assign T972 = T976[T973];
  assign T973 = T974;
  assign T974 = T975;
  assign T975 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T976 = T977;
  assign T977 = io_chanxy_in[9'h150/* 336*/:9'h148/* 328*/];
  assign T978 = T979;
  assign T979 = T980;
  assign T980 = T984[T981];
  assign T981 = T982;
  assign T982 = T983;
  assign T983 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T984 = T985;
  assign T985 = io_chanxy_in[9'h152/* 338*/:9'h151/* 337*/];
  assign T986 = T987;
  assign T987 = T988;
  assign T988 = T992[T989];
  assign T989 = T990;
  assign T990 = T991;
  assign T991 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T992 = T993;
  assign T993 = io_chanxy_in[9'h154/* 340*/:9'h153/* 339*/];
  assign T994 = T995;
  assign T995 = T996;
  assign T996 = T1000[T997];
  assign T997 = T998;
  assign T998 = T999;
  assign T999 = io_chanxy_config[8'ha2/* 162*/:8'ha2/* 162*/];
  assign T1000 = T1001;
  assign T1001 = io_chanxy_in[9'h156/* 342*/:9'h155/* 341*/];
  assign T1002 = T1003;
  assign T1003 = T1004;
  assign T1004 = T1008[T1005];
  assign T1005 = T1006;
  assign T1006 = T1007;
  assign T1007 = io_chanxy_config[8'ha3/* 163*/:8'ha3/* 163*/];
  assign T1008 = T1009;
  assign T1009 = io_chanxy_in[9'h158/* 344*/:9'h157/* 343*/];
  assign T1010 = T1011;
  assign T1011 = T1012;
  assign T1012 = T1016[T1013];
  assign T1013 = T1014;
  assign T1014 = T1015;
  assign T1015 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T1016 = T1017;
  assign T1017 = io_chanxy_in[9'h161/* 353*/:9'h159/* 345*/];
  assign T1018 = T1019;
  assign T1019 = T1020;
  assign T1020 = T1024[T1021];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T1024 = T1025;
  assign T1025 = io_chanxy_in[9'h163/* 355*/:9'h162/* 354*/];
  assign T1026 = T1027;
  assign T1027 = T1028;
  assign T1028 = T1032[T1029];
  assign T1029 = T1030;
  assign T1030 = T1031;
  assign T1031 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T1032 = T1033;
  assign T1033 = io_chanxy_in[9'h165/* 357*/:9'h164/* 356*/];
  assign T1034 = T1035;
  assign T1035 = T1036;
  assign T1036 = T1040[T1037];
  assign T1037 = T1038;
  assign T1038 = T1039;
  assign T1039 = io_chanxy_config[8'haa/* 170*/:8'haa/* 170*/];
  assign T1040 = T1041;
  assign T1041 = io_chanxy_in[9'h167/* 359*/:9'h166/* 358*/];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = T1048[T1045];
  assign T1045 = T1046;
  assign T1046 = T1047;
  assign T1047 = io_chanxy_config[8'hab/* 171*/:8'hab/* 171*/];
  assign T1048 = T1049;
  assign T1049 = io_chanxy_in[9'h169/* 361*/:9'h168/* 360*/];
  assign T1050 = T1051;
  assign T1051 = T1052;
  assign T1052 = T1056[T1053];
  assign T1053 = T1054;
  assign T1054 = T1055;
  assign T1055 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T1056 = T1057;
  assign T1057 = io_chanxy_in[9'h172/* 370*/:9'h16a/* 362*/];
  assign T1058 = T1059;
  assign T1059 = T1060;
  assign T1060 = T1064[T1061];
  assign T1061 = T1062;
  assign T1062 = T1063;
  assign T1063 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T1064 = T1065;
  assign T1065 = io_chanxy_in[9'h174/* 372*/:9'h173/* 371*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1072[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T1072 = T1073;
  assign T1073 = io_chanxy_in[9'h176/* 374*/:9'h175/* 373*/];
  assign T1074 = T1075;
  assign T1075 = T1076;
  assign T1076 = T1080[T1077];
  assign T1077 = T1078;
  assign T1078 = T1079;
  assign T1079 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T1080 = T1081;
  assign T1081 = io_chanxy_in[9'h178/* 376*/:9'h177/* 375*/];
  assign T1082 = T1083;
  assign T1083 = T1084;
  assign T1084 = T1088[T1085];
  assign T1085 = T1086;
  assign T1086 = T1087;
  assign T1087 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1088 = T1089;
  assign T1089 = io_chanxy_in[9'h17a/* 378*/:9'h179/* 377*/];
  assign T1090 = T1091;
  assign T1091 = T1092;
  assign T1092 = T1096[T1093];
  assign T1093 = T1094;
  assign T1094 = T1095;
  assign T1095 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T1096 = T1097;
  assign T1097 = io_chanxy_in[9'h183/* 387*/:9'h17b/* 379*/];
  assign T1098 = T1099;
  assign T1099 = T1100;
  assign T1100 = T1104[T1101];
  assign T1101 = T1102;
  assign T1102 = T1103;
  assign T1103 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1104 = T1105;
  assign T1105 = io_chanxy_in[9'h185/* 389*/:9'h184/* 388*/];
  assign T1106 = T1107;
  assign T1107 = T1108;
  assign T1108 = T1112[T1109];
  assign T1109 = T1110;
  assign T1110 = T1111;
  assign T1111 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T1112 = T1113;
  assign T1113 = io_chanxy_in[9'h187/* 391*/:9'h186/* 390*/];
  assign T1114 = T1115;
  assign T1115 = T1116;
  assign T1116 = T1120[T1117];
  assign T1117 = T1118;
  assign T1118 = T1119;
  assign T1119 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T1120 = T1121;
  assign T1121 = io_chanxy_in[9'h189/* 393*/:9'h188/* 392*/];
  assign T1122 = T1123;
  assign T1123 = T1124;
  assign T1124 = T1128[T1125];
  assign T1125 = T1126;
  assign T1126 = T1127;
  assign T1127 = io_chanxy_config[8'hbb/* 187*/:8'hbb/* 187*/];
  assign T1128 = T1129;
  assign T1129 = io_chanxy_in[9'h18b/* 395*/:9'h18a/* 394*/];
  assign T1130 = T1131;
  assign T1131 = T1132;
  assign T1132 = T1136[T1133];
  assign T1133 = T1134;
  assign T1134 = T1135;
  assign T1135 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T1136 = T1137;
  assign T1137 = io_chanxy_in[9'h194/* 404*/:9'h18c/* 396*/];
  assign T1138 = T1139;
  assign T1139 = T1140;
  assign T1140 = T1144[T1141];
  assign T1141 = T1142;
  assign T1142 = T1143;
  assign T1143 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1144 = T1145;
  assign T1145 = io_chanxy_in[9'h196/* 406*/:9'h195/* 405*/];
  assign T1146 = T1147;
  assign T1147 = T1148;
  assign T1148 = T1152[T1149];
  assign T1149 = T1150;
  assign T1150 = T1151;
  assign T1151 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T1152 = T1153;
  assign T1153 = io_chanxy_in[9'h198/* 408*/:9'h197/* 407*/];
  assign T1154 = T1155;
  assign T1155 = T1156;
  assign T1156 = T1160[T1157];
  assign T1157 = T1158;
  assign T1158 = T1159;
  assign T1159 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1160 = T1161;
  assign T1161 = io_chanxy_in[9'h19a/* 410*/:9'h199/* 409*/];
  assign T1162 = T1163;
  assign T1163 = T1164;
  assign T1164 = T1168[T1165];
  assign T1165 = T1166;
  assign T1166 = T1167;
  assign T1167 = io_chanxy_config[8'hc3/* 195*/:8'hc3/* 195*/];
  assign T1168 = T1169;
  assign T1169 = io_chanxy_in[9'h19c/* 412*/:9'h19b/* 411*/];
  assign T1170 = T1171;
  assign T1171 = T1172;
  assign T1172 = T1176[T1173];
  assign T1173 = T1174;
  assign T1174 = T1175;
  assign T1175 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T1176 = T1177;
  assign T1177 = io_chanxy_in[9'h1a5/* 421*/:9'h19d/* 413*/];
  assign T1178 = T1179;
  assign T1179 = T1180;
  assign T1180 = T1184[T1181];
  assign T1181 = T1182;
  assign T1182 = T1183;
  assign T1183 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T1184 = T1185;
  assign T1185 = io_chanxy_in[9'h1a7/* 423*/:9'h1a6/* 422*/];
  assign T1186 = T1187;
  assign T1187 = T1188;
  assign T1188 = T1192[T1189];
  assign T1189 = T1190;
  assign T1190 = T1191;
  assign T1191 = io_chanxy_config[8'hc9/* 201*/:8'hc9/* 201*/];
  assign T1192 = T1193;
  assign T1193 = io_chanxy_in[9'h1a9/* 425*/:9'h1a8/* 424*/];
  assign T1194 = T1195;
  assign T1195 = T1196;
  assign T1196 = T1200[T1197];
  assign T1197 = T1198;
  assign T1198 = T1199;
  assign T1199 = io_chanxy_config[8'hca/* 202*/:8'hca/* 202*/];
  assign T1200 = T1201;
  assign T1201 = io_chanxy_in[9'h1ab/* 427*/:9'h1aa/* 426*/];
  assign T1202 = T1203;
  assign T1203 = T1204;
  assign T1204 = T1208[T1205];
  assign T1205 = T1206;
  assign T1206 = T1207;
  assign T1207 = io_chanxy_config[8'hcb/* 203*/:8'hcb/* 203*/];
  assign T1208 = T1209;
  assign T1209 = io_chanxy_in[9'h1ad/* 429*/:9'h1ac/* 428*/];
  assign T1210 = T1211;
  assign T1211 = T1212;
  assign T1212 = T1216[T1213];
  assign T1213 = T1214;
  assign T1214 = T1215;
  assign T1215 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T1216 = T1217;
  assign T1217 = io_chanxy_in[9'h1b6/* 438*/:9'h1ae/* 430*/];
  assign T1218 = T1219;
  assign T1219 = T1220;
  assign T1220 = T1224[T1221];
  assign T1221 = T1222;
  assign T1222 = T1223;
  assign T1223 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T1224 = T1225;
  assign T1225 = io_chanxy_in[9'h1b8/* 440*/:9'h1b7/* 439*/];
  assign T1226 = T1227;
  assign T1227 = T1228;
  assign T1228 = T1232[T1229];
  assign T1229 = T1230;
  assign T1230 = T1231;
  assign T1231 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T1232 = T1233;
  assign T1233 = io_chanxy_in[9'h1ba/* 442*/:9'h1b9/* 441*/];
  assign T1234 = T1235;
  assign T1235 = T1236;
  assign T1236 = T1240[T1237];
  assign T1237 = T1238;
  assign T1238 = T1239;
  assign T1239 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T1240 = T1241;
  assign T1241 = io_chanxy_in[9'h1bc/* 444*/:9'h1bb/* 443*/];
  assign T1242 = T1243;
  assign T1243 = T1244;
  assign T1244 = T1248[T1245];
  assign T1245 = T1246;
  assign T1246 = T1247;
  assign T1247 = io_chanxy_config[8'hd3/* 211*/:8'hd3/* 211*/];
  assign T1248 = T1249;
  assign T1249 = io_chanxy_in[9'h1be/* 446*/:9'h1bd/* 445*/];
  assign T1250 = T1251;
  assign T1251 = T1252;
  assign T1252 = T1256[T1253];
  assign T1253 = T1254;
  assign T1254 = T1255;
  assign T1255 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T1256 = T1257;
  assign T1257 = io_chanxy_in[9'h1c7/* 455*/:9'h1bf/* 447*/];
  assign T1258 = T1259;
  assign T1259 = T1260;
  assign T1260 = T1264[T1261];
  assign T1261 = T1262;
  assign T1262 = T1263;
  assign T1263 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T1264 = T1265;
  assign T1265 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T1266 = T1267;
  assign T1267 = T1268;
  assign T1268 = T1272[T1269];
  assign T1269 = T1270;
  assign T1270 = T1271;
  assign T1271 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T1272 = T1273;
  assign T1273 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T1274 = T1275;
  assign T1275 = T1276;
  assign T1276 = T1280[T1277];
  assign T1277 = T1278;
  assign T1278 = T1279;
  assign T1279 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T1280 = T1281;
  assign T1281 = io_chanxy_in[9'h1cd/* 461*/:9'h1cc/* 460*/];
  assign T1282 = T1283;
  assign T1283 = T1284;
  assign T1284 = T1288[T1285];
  assign T1285 = T1286;
  assign T1286 = T1287;
  assign T1287 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T1288 = T1289;
  assign T1289 = io_chanxy_in[9'h1cf/* 463*/:9'h1ce/* 462*/];
  assign T1290 = T1291;
  assign T1291 = T1292;
  assign T1292 = T1296[T1293];
  assign T1293 = T1294;
  assign T1294 = T1295;
  assign T1295 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1296 = T1297;
  assign T1297 = io_chanxy_in[9'h1d8/* 472*/:9'h1d0/* 464*/];
  assign T1298 = T1299;
  assign T1299 = T1300;
  assign T1300 = T1304[T1301];
  assign T1301 = T1302;
  assign T1302 = T1303;
  assign T1303 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T1304 = T1305;
  assign T1305 = io_chanxy_in[9'h1da/* 474*/:9'h1d9/* 473*/];
  assign T1306 = T1307;
  assign T1307 = T1308;
  assign T1308 = T1312[T1309];
  assign T1309 = T1310;
  assign T1310 = T1311;
  assign T1311 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T1312 = T1313;
  assign T1313 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T1314 = T1315;
  assign T1315 = T1316;
  assign T1316 = T1320[T1317];
  assign T1317 = T1318;
  assign T1318 = T1319;
  assign T1319 = io_chanxy_config[8'he2/* 226*/:8'he2/* 226*/];
  assign T1320 = T1321;
  assign T1321 = io_chanxy_in[9'h1de/* 478*/:9'h1dd/* 477*/];
  assign T1322 = T1323;
  assign T1323 = T1324;
  assign T1324 = T1328[T1325];
  assign T1325 = T1326;
  assign T1326 = T1327;
  assign T1327 = io_chanxy_config[8'he3/* 227*/:8'he3/* 227*/];
  assign T1328 = T1329;
  assign T1329 = io_chanxy_in[9'h1e0/* 480*/:9'h1df/* 479*/];
  assign T1330 = T1331;
  assign T1331 = T1332;
  assign T1332 = T1336[T1333];
  assign T1333 = T1334;
  assign T1334 = T1335;
  assign T1335 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T1336 = T1337;
  assign T1337 = io_chanxy_in[9'h1e9/* 489*/:9'h1e1/* 481*/];
  assign T1338 = T1339;
  assign T1339 = T1340;
  assign T1340 = T1344[T1341];
  assign T1341 = T1342;
  assign T1342 = T1343;
  assign T1343 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T1344 = T1345;
  assign T1345 = io_chanxy_in[9'h1eb/* 491*/:9'h1ea/* 490*/];
  assign T1346 = T1347;
  assign T1347 = T1348;
  assign T1348 = T1352[T1349];
  assign T1349 = T1350;
  assign T1350 = T1351;
  assign T1351 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T1352 = T1353;
  assign T1353 = io_chanxy_in[9'h1ed/* 493*/:9'h1ec/* 492*/];
  assign T1354 = T1355;
  assign T1355 = T1356;
  assign T1356 = T1360[T1357];
  assign T1357 = T1358;
  assign T1358 = T1359;
  assign T1359 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T1360 = T1361;
  assign T1361 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T1362 = T1363;
  assign T1363 = T1364;
  assign T1364 = T1368[T1365];
  assign T1365 = T1366;
  assign T1366 = T1367;
  assign T1367 = io_chanxy_config[8'heb/* 235*/:8'heb/* 235*/];
  assign T1368 = T1369;
  assign T1369 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T1370 = T1371;
  assign T1371 = T1372;
  assign T1372 = T1376[T1373];
  assign T1373 = T1374;
  assign T1374 = T1375;
  assign T1375 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T1376 = T1377;
  assign T1377 = io_chanxy_in[9'h1fa/* 506*/:9'h1f2/* 498*/];
  assign T1378 = T1379;
  assign T1379 = T1380;
  assign T1380 = T1384[T1381];
  assign T1381 = T1382;
  assign T1382 = T1383;
  assign T1383 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T1384 = T1385;
  assign T1385 = io_chanxy_in[9'h1fc/* 508*/:9'h1fb/* 507*/];
  assign T1386 = T1387;
  assign T1387 = T1388;
  assign T1388 = T1392[T1389];
  assign T1389 = T1390;
  assign T1390 = T1391;
  assign T1391 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T1392 = T1393;
  assign T1393 = io_chanxy_in[9'h1fe/* 510*/:9'h1fd/* 509*/];
  assign T1394 = T1395;
  assign T1395 = T1396;
  assign T1396 = T1400[T1397];
  assign T1397 = T1398;
  assign T1398 = T1399;
  assign T1399 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1400 = T1401;
  assign T1401 = io_chanxy_in[10'h200/* 512*/:9'h1ff/* 511*/];
  assign T1402 = T1403;
  assign T1403 = T1404;
  assign T1404 = T1408[T1405];
  assign T1405 = T1406;
  assign T1406 = T1407;
  assign T1407 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T1408 = T1409;
  assign T1409 = io_chanxy_in[10'h202/* 514*/:10'h201/* 513*/];
  assign T1410 = T1411;
  assign T1411 = T1412;
  assign T1412 = T1416[T1413];
  assign T1413 = T1414;
  assign T1414 = T1415;
  assign T1415 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1416 = T1417;
  assign T1417 = io_chanxy_in[10'h20b/* 523*/:10'h203/* 515*/];
  assign T1418 = T1419;
  assign T1419 = T1420;
  assign T1420 = T1424[T1421];
  assign T1421 = T1422;
  assign T1422 = T1423;
  assign T1423 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1424 = T1425;
  assign T1425 = io_chanxy_in[10'h20d/* 525*/:10'h20c/* 524*/];
  assign T1426 = T1427;
  assign T1427 = T1428;
  assign T1428 = T1432[T1429];
  assign T1429 = T1430;
  assign T1430 = T1431;
  assign T1431 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T1432 = T1433;
  assign T1433 = io_chanxy_in[10'h20f/* 527*/:10'h20e/* 526*/];
  assign T1434 = T1435;
  assign T1435 = T1436;
  assign T1436 = T1440[T1437];
  assign T1437 = T1438;
  assign T1438 = T1439;
  assign T1439 = io_chanxy_config[8'hfa/* 250*/:8'hfa/* 250*/];
  assign T1440 = T1441;
  assign T1441 = io_chanxy_in[10'h211/* 529*/:10'h210/* 528*/];
  assign T1442 = T1443;
  assign T1443 = T1444;
  assign T1444 = T1448[T1445];
  assign T1445 = T1446;
  assign T1446 = T1447;
  assign T1447 = io_chanxy_config[8'hfb/* 251*/:8'hfb/* 251*/];
  assign T1448 = T1449;
  assign T1449 = io_chanxy_in[10'h213/* 531*/:10'h212/* 530*/];
  assign T1450 = T1451;
  assign T1451 = T1452;
  assign T1452 = T1456[T1453];
  assign T1453 = T1454;
  assign T1454 = T1455;
  assign T1455 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1456 = T1457;
  assign T1457 = io_chanxy_in[10'h21c/* 540*/:10'h214/* 532*/];
  assign T1458 = T1459;
  assign T1459 = T1460;
  assign T1460 = T1464[T1461];
  assign T1461 = T1462;
  assign T1462 = T1463;
  assign T1463 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1464 = T1465;
  assign T1465 = io_chanxy_in[10'h21e/* 542*/:10'h21d/* 541*/];
  assign T1466 = T1467;
  assign T1467 = T1468;
  assign T1468 = T1472[T1469];
  assign T1469 = T1470;
  assign T1470 = T1471;
  assign T1471 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1472 = T1473;
  assign T1473 = io_chanxy_in[10'h220/* 544*/:10'h21f/* 543*/];
  assign T1474 = T1475;
  assign T1475 = T1476;
  assign T1476 = T1480[T1477];
  assign T1477 = T1478;
  assign T1478 = T1479;
  assign T1479 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1480 = T1481;
  assign T1481 = io_chanxy_in[10'h222/* 546*/:10'h221/* 545*/];
  assign T1482 = T1483;
  assign T1483 = T1484;
  assign T1484 = T1488[T1485];
  assign T1485 = T1486;
  assign T1486 = T1487;
  assign T1487 = io_chanxy_config[9'h103/* 259*/:9'h103/* 259*/];
  assign T1488 = T1489;
  assign T1489 = io_chanxy_in[10'h224/* 548*/:10'h223/* 547*/];
  assign T1490 = T1491;
  assign T1491 = T1492;
  assign T1492 = T1496[T1493];
  assign T1493 = T1494;
  assign T1494 = T1495;
  assign T1495 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1496 = T1497;
  assign T1497 = io_chanxy_in[10'h22d/* 557*/:10'h225/* 549*/];
  assign io_ipin_out = T1498;
  assign T1498 = T1499;
  assign T1499 = {T1718, T1500};
  assign T1500 = T1501;
  assign T1501 = {T1710, T1502};
  assign T1502 = T1503;
  assign T1503 = {T1702, T1504};
  assign T1504 = T1505;
  assign T1505 = {T1694, T1506};
  assign T1506 = T1507;
  assign T1507 = {T1686, T1508};
  assign T1508 = T1509;
  assign T1509 = {T1678, T1510};
  assign T1510 = T1511;
  assign T1511 = {T1670, T1512};
  assign T1512 = T1513;
  assign T1513 = {T1662, T1514};
  assign T1514 = T1515;
  assign T1515 = {T1654, T1516};
  assign T1516 = T1517;
  assign T1517 = {T1646, T1518};
  assign T1518 = T1519;
  assign T1519 = {T1638, T1520};
  assign T1520 = T1521;
  assign T1521 = {T1630, T1522};
  assign T1522 = T1523;
  assign T1523 = {T1622, T1524};
  assign T1524 = T1525;
  assign T1525 = {T1614, T1526};
  assign T1526 = T1527;
  assign T1527 = {T1606, T1528};
  assign T1528 = T1529;
  assign T1529 = {T1598, T1530};
  assign T1530 = T1531;
  assign T1531 = {T1590, T1532};
  assign T1532 = T1533;
  assign T1533 = {T1582, T1534};
  assign T1534 = T1535;
  assign T1535 = {T1574, T1536};
  assign T1536 = T1537;
  assign T1537 = {T1566, T1538};
  assign T1538 = T1539;
  assign T1539 = {T1558, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1550, T1542};
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_10(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [557:0] io_chanxy_in,
    output[149:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[149:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_6 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_7(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [572:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[1:0] T211;
  wire[1:0] T212;
  wire[1:0] T213;
  wire[2:0] T214;
  wire[2:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[1:0] T219;
  wire[1:0] T220;
  wire[1:0] T221;
  wire[2:0] T222;
  wire[2:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[1:0] T227;
  wire[1:0] T228;
  wire[1:0] T229;
  wire[2:0] T230;
  wire[2:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[1:0] T236;
  wire[1:0] T237;
  wire[2:0] T238;
  wire[2:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire[1:0] T244;
  wire[1:0] T245;
  wire[2:0] T246;
  wire[2:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[1:0] T251;
  wire[1:0] T252;
  wire[1:0] T253;
  wire[2:0] T254;
  wire[2:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire[1:0] T262;
  wire[1:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire[1:0] T270;
  wire[1:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire[1:0] T278;
  wire[1:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire[1:0] T286;
  wire[1:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire[1:0] T294;
  wire[1:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire[1:0] T302;
  wire[1:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire[1:0] T310;
  wire[1:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire[1:0] T318;
  wire[1:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire[1:0] T326;
  wire[1:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[1:0] T331;
  wire[1:0] T332;
  wire[1:0] T333;
  wire[2:0] T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[1:0] T339;
  wire[1:0] T340;
  wire[1:0] T341;
  wire[2:0] T342;
  wire[2:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[1:0] T347;
  wire[1:0] T348;
  wire[1:0] T349;
  wire[2:0] T350;
  wire[2:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[1:0] T355;
  wire[1:0] T356;
  wire[1:0] T357;
  wire[2:0] T358;
  wire[2:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[1:0] T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[2:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[1:0] T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire[2:0] T374;
  wire[2:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire[1:0] T382;
  wire[1:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire[1:0] T390;
  wire[1:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire[1:0] T398;
  wire[1:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire[1:0] T406;
  wire[1:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire[1:0] T414;
  wire[1:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire[1:0] T422;
  wire[1:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire[1:0] T430;
  wire[1:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire[1:0] T438;
  wire[1:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire[1:0] T446;
  wire[1:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[1:0] T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[1:0] T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire[2:0] T470;
  wire[2:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[1:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[2:0] T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[1:0] T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire[2:0] T486;
  wire[2:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[3:0] T571;
  wire[3:0] T572;
  wire[3:0] T573;
  wire[10:0] T574;
  wire[10:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[2:0] T582;
  wire[2:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[3:0] T587;
  wire[3:0] T588;
  wire[3:0] T589;
  wire[10:0] T590;
  wire[10:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire[2:0] T598;
  wire[2:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[3:0] T603;
  wire[3:0] T604;
  wire[3:0] T605;
  wire[10:0] T606;
  wire[10:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[3:0] T619;
  wire[3:0] T620;
  wire[3:0] T621;
  wire[10:0] T622;
  wire[10:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[1:0] T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire[2:0] T630;
  wire[2:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[3:0] T635;
  wire[3:0] T636;
  wire[3:0] T637;
  wire[10:0] T638;
  wire[10:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[1:0] T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire[2:0] T646;
  wire[2:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire[3:0] T651;
  wire[3:0] T652;
  wire[3:0] T653;
  wire[10:0] T654;
  wire[10:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[1:0] T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire[2:0] T662;
  wire[2:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[3:0] T667;
  wire[3:0] T668;
  wire[3:0] T669;
  wire[10:0] T670;
  wire[10:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[1:0] T678;
  wire[1:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[3:0] T683;
  wire[3:0] T684;
  wire[3:0] T685;
  wire[10:0] T686;
  wire[10:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire[3:0] T699;
  wire[3:0] T700;
  wire[3:0] T701;
  wire[10:0] T702;
  wire[10:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire[3:0] T715;
  wire[3:0] T716;
  wire[3:0] T717;
  wire[9:0] T718;
  wire[9:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire[3:0] T731;
  wire[3:0] T732;
  wire[3:0] T733;
  wire[9:0] T734;
  wire[9:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire[3:0] T747;
  wire[3:0] T748;
  wire[3:0] T749;
  wire[9:0] T750;
  wire[9:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire[3:0] T763;
  wire[3:0] T764;
  wire[3:0] T765;
  wire[9:0] T766;
  wire[9:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire[3:0] T779;
  wire[3:0] T780;
  wire[3:0] T781;
  wire[9:0] T782;
  wire[9:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire[3:0] T795;
  wire[3:0] T796;
  wire[3:0] T797;
  wire[9:0] T798;
  wire[9:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[8:0] T814;
  wire[8:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[8:0] T822;
  wire[8:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[8:0] T830;
  wire[8:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[8:0] T838;
  wire[8:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[8:0] T846;
  wire[8:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[3:0] T851;
  wire[3:0] T852;
  wire[3:0] T853;
  wire[8:0] T854;
  wire[8:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[8:0] T862;
  wire[8:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[8:0] T870;
  wire[8:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[8:0] T878;
  wire[8:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[8:0] T886;
  wire[8:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[8:0] T894;
  wire[8:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[8:0] T902;
  wire[8:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[8:0] T910;
  wire[8:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[8:0] T918;
  wire[8:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[8:0] T926;
  wire[8:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire[3:0] T931;
  wire[3:0] T932;
  wire[3:0] T933;
  wire[8:0] T934;
  wire[8:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[8:0] T942;
  wire[8:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[8:0] T950;
  wire[8:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[8:0] T958;
  wire[8:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[8:0] T966;
  wire[8:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[8:0] T974;
  wire[8:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[8:0] T982;
  wire[8:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[8:0] T990;
  wire[8:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[8:0] T998;
  wire[8:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[8:0] T1006;
  wire[8:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire[3:0] T1011;
  wire[3:0] T1012;
  wire[3:0] T1013;
  wire[8:0] T1014;
  wire[8:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[8:0] T1022;
  wire[8:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[8:0] T1030;
  wire[8:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[8:0] T1038;
  wire[8:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[8:0] T1046;
  wire[8:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[4'he/* 14*/:4'hc/* 12*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[5'h11/* 17*/:4'hf/* 15*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[5'h16/* 22*/:5'h15/* 21*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[6'h26/* 38*/:6'h24/* 36*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[5'h18/* 24*/:5'h17/* 23*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[6'h29/* 41*/:6'h27/* 39*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[5'h1a/* 26*/:5'h19/* 25*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[6'h2c/* 44*/:6'h2a/* 42*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[5'h1c/* 28*/:5'h1b/* 27*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[6'h2f/* 47*/:6'h2d/* 45*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[5'h1e/* 30*/:5'h1d/* 29*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[6'h32/* 50*/:6'h30/* 48*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[6'h20/* 32*/:5'h1f/* 31*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[6'h35/* 53*/:6'h33/* 51*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[7'h50/* 80*/:7'h4e/* 78*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[7'h53/* 83*/:7'h51/* 81*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[7'h56/* 86*/:7'h54/* 84*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[7'h59/* 89*/:7'h57/* 87*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[6'h3c/* 60*/:6'h3c/* 60*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[6'h3d/* 61*/:6'h3d/* 61*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[6'h3e/* 62*/:6'h3e/* 62*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[7'h42/* 66*/:6'h3f/* 63*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[7'h76/* 118*/:7'h6c/* 108*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[7'h44/* 68*/:7'h43/* 67*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[7'h79/* 121*/:7'h77/* 119*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[7'h48/* 72*/:7'h45/* 69*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[8'h84/* 132*/:7'h7a/* 122*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[7'h4a/* 74*/:7'h49/* 73*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[8'h87/* 135*/:8'h85/* 133*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[8'h92/* 146*/:8'h88/* 136*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[7'h50/* 80*/:7'h4f/* 79*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[8'h95/* 149*/:8'h93/* 147*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[7'h54/* 84*/:7'h51/* 81*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[8'ha0/* 160*/:8'h96/* 150*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[7'h56/* 86*/:7'h55/* 85*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[7'h5a/* 90*/:7'h57/* 87*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[8'hae/* 174*/:8'ha4/* 164*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[7'h5c/* 92*/:7'h5b/* 91*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[8'hb1/* 177*/:8'haf/* 175*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[7'h60/* 96*/:7'h5d/* 93*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[8'hbc/* 188*/:8'hb2/* 178*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[7'h62/* 98*/:7'h61/* 97*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[8'hbf/* 191*/:8'hbd/* 189*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[7'h66/* 102*/:7'h63/* 99*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[8'hcc/* 204*/:8'hcb/* 203*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[8'hd7/* 215*/:8'hcd/* 205*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[7'h6c/* 108*/:7'h6c/* 108*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[7'h70/* 112*/:7'h6d/* 109*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[8'he4/* 228*/:8'hda/* 218*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[8'he6/* 230*/:8'he5/* 229*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[8'hf0/* 240*/:8'he7/* 231*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[7'h76/* 118*/:7'h76/* 118*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[8'hf2/* 242*/:8'hf1/* 241*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[7'h7a/* 122*/:7'h77/* 119*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[8'hfc/* 252*/:8'hf3/* 243*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[7'h7b/* 123*/:7'h7b/* 123*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h108/* 264*/:8'hff/* 255*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'h84/* 132*/:8'h81/* 129*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h114/* 276*/:9'h10b/* 267*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h116/* 278*/:9'h115/* 277*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'h89/* 137*/:8'h86/* 134*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h120/* 288*/:9'h117/* 279*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h12c/* 300*/:9'h123/* 291*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h137/* 311*/:9'h12f/* 303*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h140/* 320*/:9'h138/* 312*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h149/* 329*/:9'h141/* 321*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h152/* 338*/:9'h14a/* 330*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h15b/* 347*/:9'h153/* 339*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h164/* 356*/:9'h15c/* 348*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h16d/* 365*/:9'h165/* 357*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h176/* 374*/:9'h16e/* 366*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h17f/* 383*/:9'h177/* 375*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h188/* 392*/:9'h180/* 384*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h191/* 401*/:9'h189/* 393*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h19a/* 410*/:9'h192/* 402*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1a3/* 419*/:9'h19b/* 411*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1ac/* 428*/:9'h1a4/* 420*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1b5/* 437*/:9'h1ad/* 429*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1be/* 446*/:9'h1b6/* 438*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1c7/* 455*/:9'h1bf/* 447*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1d0/* 464*/:9'h1c8/* 456*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1d9/* 473*/:9'h1d1/* 465*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[9'h1e2/* 482*/:9'h1da/* 474*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[9'h1eb/* 491*/:9'h1e3/* 483*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[9'h1f4/* 500*/:9'h1ec/* 492*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[9'h1fd/* 509*/:9'h1f5/* 501*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h206/* 518*/:9'h1fe/* 510*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h20f/* 527*/:10'h207/* 519*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h218/* 536*/:10'h210/* 528*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h221/* 545*/:10'h219/* 537*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h22a/* 554*/:10'h222/* 546*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h233/* 563*/:10'h22b/* 555*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h23c/* 572*/:10'h234/* 564*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_11(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_12(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_13(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_14(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_15(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_16(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_17(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_18(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


module sbcb_sp_8(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [509:0] io_chanxy_in,
    input [239:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[149:0] io_chanxy_out);

  wire[149:0] T0;
  wire[149:0] T1;
  wire[148:0] T2;
  wire[148:0] T3;
  wire[147:0] T4;
  wire[147:0] T5;
  wire[146:0] T6;
  wire[146:0] T7;
  wire[145:0] T8;
  wire[145:0] T9;
  wire[144:0] T10;
  wire[144:0] T11;
  wire[143:0] T12;
  wire[143:0] T13;
  wire[142:0] T14;
  wire[142:0] T15;
  wire[141:0] T16;
  wire[141:0] T17;
  wire[140:0] T18;
  wire[140:0] T19;
  wire[139:0] T20;
  wire[139:0] T21;
  wire[138:0] T22;
  wire[138:0] T23;
  wire[137:0] T24;
  wire[137:0] T25;
  wire[136:0] T26;
  wire[136:0] T27;
  wire[135:0] T28;
  wire[135:0] T29;
  wire[134:0] T30;
  wire[134:0] T31;
  wire[133:0] T32;
  wire[133:0] T33;
  wire[132:0] T34;
  wire[132:0] T35;
  wire[131:0] T36;
  wire[131:0] T37;
  wire[130:0] T38;
  wire[130:0] T39;
  wire[129:0] T40;
  wire[129:0] T41;
  wire[128:0] T42;
  wire[128:0] T43;
  wire[127:0] T44;
  wire[127:0] T45;
  wire[126:0] T46;
  wire[126:0] T47;
  wire[125:0] T48;
  wire[125:0] T49;
  wire[124:0] T50;
  wire[124:0] T51;
  wire[123:0] T52;
  wire[123:0] T53;
  wire[122:0] T54;
  wire[122:0] T55;
  wire[121:0] T56;
  wire[121:0] T57;
  wire[120:0] T58;
  wire[120:0] T59;
  wire[119:0] T60;
  wire[119:0] T61;
  wire[118:0] T62;
  wire[118:0] T63;
  wire[117:0] T64;
  wire[117:0] T65;
  wire[116:0] T66;
  wire[116:0] T67;
  wire[115:0] T68;
  wire[115:0] T69;
  wire[114:0] T70;
  wire[114:0] T71;
  wire[113:0] T72;
  wire[113:0] T73;
  wire[112:0] T74;
  wire[112:0] T75;
  wire[111:0] T76;
  wire[111:0] T77;
  wire[110:0] T78;
  wire[110:0] T79;
  wire[109:0] T80;
  wire[109:0] T81;
  wire[108:0] T82;
  wire[108:0] T83;
  wire[107:0] T84;
  wire[107:0] T85;
  wire[106:0] T86;
  wire[106:0] T87;
  wire[105:0] T88;
  wire[105:0] T89;
  wire[104:0] T90;
  wire[104:0] T91;
  wire[103:0] T92;
  wire[103:0] T93;
  wire[102:0] T94;
  wire[102:0] T95;
  wire[101:0] T96;
  wire[101:0] T97;
  wire[100:0] T98;
  wire[100:0] T99;
  wire[99:0] T100;
  wire[99:0] T101;
  wire[98:0] T102;
  wire[98:0] T103;
  wire[97:0] T104;
  wire[97:0] T105;
  wire[96:0] T106;
  wire[96:0] T107;
  wire[95:0] T108;
  wire[95:0] T109;
  wire[94:0] T110;
  wire[94:0] T111;
  wire[93:0] T112;
  wire[93:0] T113;
  wire[92:0] T114;
  wire[92:0] T115;
  wire[91:0] T116;
  wire[91:0] T117;
  wire[90:0] T118;
  wire[90:0] T119;
  wire[89:0] T120;
  wire[89:0] T121;
  wire[88:0] T122;
  wire[88:0] T123;
  wire[87:0] T124;
  wire[87:0] T125;
  wire[86:0] T126;
  wire[86:0] T127;
  wire[85:0] T128;
  wire[85:0] T129;
  wire[84:0] T130;
  wire[84:0] T131;
  wire[83:0] T132;
  wire[83:0] T133;
  wire[82:0] T134;
  wire[82:0] T135;
  wire[81:0] T136;
  wire[81:0] T137;
  wire[80:0] T138;
  wire[80:0] T139;
  wire[79:0] T140;
  wire[79:0] T141;
  wire[78:0] T142;
  wire[78:0] T143;
  wire[77:0] T144;
  wire[77:0] T145;
  wire[76:0] T146;
  wire[76:0] T147;
  wire[75:0] T148;
  wire[75:0] T149;
  wire[74:0] T150;
  wire[74:0] T151;
  wire[73:0] T152;
  wire[73:0] T153;
  wire[72:0] T154;
  wire[72:0] T155;
  wire[71:0] T156;
  wire[71:0] T157;
  wire[70:0] T158;
  wire[70:0] T159;
  wire[69:0] T160;
  wire[69:0] T161;
  wire[68:0] T162;
  wire[68:0] T163;
  wire[67:0] T164;
  wire[67:0] T165;
  wire[66:0] T166;
  wire[66:0] T167;
  wire[65:0] T168;
  wire[65:0] T169;
  wire[64:0] T170;
  wire[64:0] T171;
  wire[63:0] T172;
  wire[63:0] T173;
  wire[62:0] T174;
  wire[62:0] T175;
  wire[61:0] T176;
  wire[61:0] T177;
  wire[60:0] T178;
  wire[60:0] T179;
  wire[59:0] T180;
  wire[59:0] T181;
  wire[58:0] T182;
  wire[58:0] T183;
  wire[57:0] T184;
  wire[57:0] T185;
  wire[56:0] T186;
  wire[56:0] T187;
  wire[55:0] T188;
  wire[55:0] T189;
  wire[54:0] T190;
  wire[54:0] T191;
  wire[53:0] T192;
  wire[53:0] T193;
  wire[52:0] T194;
  wire[52:0] T195;
  wire[51:0] T196;
  wire[51:0] T197;
  wire[50:0] T198;
  wire[50:0] T199;
  wire[49:0] T200;
  wire[49:0] T201;
  wire[48:0] T202;
  wire[48:0] T203;
  wire[47:0] T204;
  wire[47:0] T205;
  wire[46:0] T206;
  wire[46:0] T207;
  wire[45:0] T208;
  wire[45:0] T209;
  wire[44:0] T210;
  wire[44:0] T211;
  wire[43:0] T212;
  wire[43:0] T213;
  wire[42:0] T214;
  wire[42:0] T215;
  wire[41:0] T216;
  wire[41:0] T217;
  wire[40:0] T218;
  wire[40:0] T219;
  wire[39:0] T220;
  wire[39:0] T221;
  wire[38:0] T222;
  wire[38:0] T223;
  wire[37:0] T224;
  wire[37:0] T225;
  wire[36:0] T226;
  wire[36:0] T227;
  wire[35:0] T228;
  wire[35:0] T229;
  wire[34:0] T230;
  wire[34:0] T231;
  wire[33:0] T232;
  wire[33:0] T233;
  wire[32:0] T234;
  wire[32:0] T235;
  wire[31:0] T236;
  wire[31:0] T237;
  wire[30:0] T238;
  wire[30:0] T239;
  wire[29:0] T240;
  wire[29:0] T241;
  wire[28:0] T242;
  wire[28:0] T243;
  wire[27:0] T244;
  wire[27:0] T245;
  wire[26:0] T246;
  wire[26:0] T247;
  wire[25:0] T248;
  wire[25:0] T249;
  wire[24:0] T250;
  wire[24:0] T251;
  wire[23:0] T252;
  wire[23:0] T253;
  wire[22:0] T254;
  wire[22:0] T255;
  wire[21:0] T256;
  wire[21:0] T257;
  wire[20:0] T258;
  wire[20:0] T259;
  wire[19:0] T260;
  wire[19:0] T261;
  wire[18:0] T262;
  wire[18:0] T263;
  wire[17:0] T264;
  wire[17:0] T265;
  wire[16:0] T266;
  wire[16:0] T267;
  wire[15:0] T268;
  wire[15:0] T269;
  wire[14:0] T270;
  wire[14:0] T271;
  wire[13:0] T272;
  wire[13:0] T273;
  wire[12:0] T274;
  wire[12:0] T275;
  wire[11:0] T276;
  wire[11:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire[9:0] T280;
  wire[9:0] T281;
  wire[8:0] T282;
  wire[8:0] T283;
  wire[7:0] T284;
  wire[7:0] T285;
  wire[6:0] T286;
  wire[6:0] T287;
  wire[5:0] T288;
  wire[5:0] T289;
  wire[4:0] T290;
  wire[4:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[2:0] T294;
  wire[2:0] T295;
  wire[1:0] T296;
  wire[1:0] T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire[1:0] T304;
  wire[1:0] T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  wire[1:0] T312;
  wire[1:0] T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  wire[1:0] T320;
  wire[1:0] T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire[1:0] T328;
  wire[1:0] T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  wire[1:0] T336;
  wire[1:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[1:0] T344;
  wire[1:0] T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  wire[1:0] T352;
  wire[1:0] T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire[1:0] T360;
  wire[1:0] T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire[1:0] T368;
  wire[1:0] T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire[1:0] T376;
  wire[1:0] T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire[1:0] T384;
  wire[1:0] T385;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire[1:0] T393;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire[1:0] T401;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire[1:0] T408;
  wire[1:0] T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire[1:0] T416;
  wire[1:0] T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[1:0] T424;
  wire[1:0] T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire[1:0] T432;
  wire[1:0] T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire[1:0] T440;
  wire[1:0] T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire[1:0] T448;
  wire[1:0] T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire[1:0] T456;
  wire[1:0] T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire[1:0] T464;
  wire[1:0] T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire T470;
  wire T471;
  wire[1:0] T472;
  wire[1:0] T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire[1:0] T480;
  wire[1:0] T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[1:0] T488;
  wire[1:0] T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire[1:0] T496;
  wire[1:0] T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire T502;
  wire T503;
  wire[1:0] T504;
  wire[1:0] T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire[1:0] T512;
  wire[1:0] T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire[1:0] T520;
  wire[1:0] T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire[1:0] T528;
  wire[1:0] T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire[1:0] T536;
  wire[1:0] T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire[1:0] T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire[1:0] T552;
  wire[1:0] T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire[1:0] T560;
  wire[1:0] T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire[1:0] T568;
  wire[1:0] T569;
  wire T570;
  wire T571;
  wire T572;
  wire T573;
  wire T574;
  wire T575;
  wire[1:0] T576;
  wire[1:0] T577;
  wire T578;
  wire T579;
  wire T580;
  wire T581;
  wire T582;
  wire T583;
  wire[1:0] T584;
  wire[1:0] T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire[1:0] T592;
  wire[1:0] T593;
  wire T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire[1:0] T600;
  wire[1:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire[1:0] T608;
  wire[1:0] T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire[1:0] T616;
  wire[1:0] T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire[1:0] T624;
  wire[1:0] T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[1:0] T632;
  wire[1:0] T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire[1:0] T640;
  wire[1:0] T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire[1:0] T648;
  wire[1:0] T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire[1:0] T656;
  wire[1:0] T657;
  wire T658;
  wire T659;
  wire T660;
  wire[3:0] T661;
  wire[3:0] T662;
  wire[3:0] T663;
  wire[8:0] T664;
  wire[8:0] T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire[1:0] T672;
  wire[1:0] T673;
  wire T674;
  wire T675;
  wire T676;
  wire[3:0] T677;
  wire[3:0] T678;
  wire[3:0] T679;
  wire[8:0] T680;
  wire[8:0] T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire[1:0] T688;
  wire[1:0] T689;
  wire T690;
  wire T691;
  wire T692;
  wire[3:0] T693;
  wire[3:0] T694;
  wire[3:0] T695;
  wire[8:0] T696;
  wire[8:0] T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire T702;
  wire T703;
  wire[1:0] T704;
  wire[1:0] T705;
  wire T706;
  wire T707;
  wire T708;
  wire[3:0] T709;
  wire[3:0] T710;
  wire[3:0] T711;
  wire[8:0] T712;
  wire[8:0] T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire T718;
  wire T719;
  wire[1:0] T720;
  wire[1:0] T721;
  wire T722;
  wire T723;
  wire T724;
  wire[3:0] T725;
  wire[3:0] T726;
  wire[3:0] T727;
  wire[8:0] T728;
  wire[8:0] T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire[1:0] T736;
  wire[1:0] T737;
  wire T738;
  wire T739;
  wire T740;
  wire[3:0] T741;
  wire[3:0] T742;
  wire[3:0] T743;
  wire[8:0] T744;
  wire[8:0] T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire[1:0] T752;
  wire[1:0] T753;
  wire T754;
  wire T755;
  wire T756;
  wire[3:0] T757;
  wire[3:0] T758;
  wire[3:0] T759;
  wire[8:0] T760;
  wire[8:0] T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire[1:0] T768;
  wire[1:0] T769;
  wire T770;
  wire T771;
  wire T772;
  wire[3:0] T773;
  wire[3:0] T774;
  wire[3:0] T775;
  wire[8:0] T776;
  wire[8:0] T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire[1:0] T784;
  wire[1:0] T785;
  wire T786;
  wire T787;
  wire T788;
  wire[3:0] T789;
  wire[3:0] T790;
  wire[3:0] T791;
  wire[8:0] T792;
  wire[8:0] T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire[1:0] T800;
  wire[1:0] T801;
  wire T802;
  wire T803;
  wire T804;
  wire[3:0] T805;
  wire[3:0] T806;
  wire[3:0] T807;
  wire[8:0] T808;
  wire[8:0] T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire[1:0] T816;
  wire[1:0] T817;
  wire T818;
  wire T819;
  wire T820;
  wire[3:0] T821;
  wire[3:0] T822;
  wire[3:0] T823;
  wire[8:0] T824;
  wire[8:0] T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire[1:0] T832;
  wire[1:0] T833;
  wire T834;
  wire T835;
  wire T836;
  wire[3:0] T837;
  wire[3:0] T838;
  wire[3:0] T839;
  wire[8:0] T840;
  wire[8:0] T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire T846;
  wire T847;
  wire[1:0] T848;
  wire[1:0] T849;
  wire T850;
  wire T851;
  wire T852;
  wire[3:0] T853;
  wire[3:0] T854;
  wire[3:0] T855;
  wire[8:0] T856;
  wire[8:0] T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire T862;
  wire T863;
  wire[1:0] T864;
  wire[1:0] T865;
  wire T866;
  wire T867;
  wire T868;
  wire[3:0] T869;
  wire[3:0] T870;
  wire[3:0] T871;
  wire[8:0] T872;
  wire[8:0] T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire[1:0] T880;
  wire[1:0] T881;
  wire T882;
  wire T883;
  wire T884;
  wire[3:0] T885;
  wire[3:0] T886;
  wire[3:0] T887;
  wire[8:0] T888;
  wire[8:0] T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire[1:0] T896;
  wire[1:0] T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire[1:0] T904;
  wire[1:0] T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T911;
  wire[1:0] T912;
  wire[1:0] T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire[1:0] T920;
  wire[1:0] T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire T926;
  wire T927;
  wire[1:0] T928;
  wire[1:0] T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire T934;
  wire T935;
  wire[1:0] T936;
  wire[1:0] T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire[1:0] T944;
  wire[1:0] T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire[1:0] T952;
  wire[1:0] T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire[1:0] T960;
  wire[1:0] T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire T966;
  wire T967;
  wire[1:0] T968;
  wire[1:0] T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire[1:0] T976;
  wire[1:0] T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire T982;
  wire T983;
  wire[1:0] T984;
  wire[1:0] T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire T990;
  wire T991;
  wire[1:0] T992;
  wire[1:0] T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[1:0] T1000;
  wire[1:0] T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire T1006;
  wire T1007;
  wire[1:0] T1008;
  wire[1:0] T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire T1014;
  wire T1015;
  wire[1:0] T1016;
  wire[1:0] T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire[1:0] T1024;
  wire[1:0] T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire[1:0] T1032;
  wire[1:0] T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire[1:0] T1040;
  wire[1:0] T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire T1046;
  wire T1047;
  wire[1:0] T1048;
  wire[1:0] T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire T1055;
  wire[1:0] T1056;
  wire[1:0] T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[1:0] T1064;
  wire[1:0] T1065;
  wire T1066;
  wire T1067;
  wire T1068;
  wire T1069;
  wire T1070;
  wire T1071;
  wire[1:0] T1072;
  wire[1:0] T1073;
  wire T1074;
  wire T1075;
  wire T1076;
  wire T1077;
  wire T1078;
  wire T1079;
  wire[1:0] T1080;
  wire[1:0] T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire[1:0] T1088;
  wire[1:0] T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire[1:0] T1096;
  wire[1:0] T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire[1:0] T1104;
  wire[1:0] T1105;
  wire T1106;
  wire T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire T1111;
  wire[1:0] T1112;
  wire[1:0] T1113;
  wire T1114;
  wire T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire[1:0] T1120;
  wire[1:0] T1121;
  wire T1122;
  wire T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire T1127;
  wire[1:0] T1128;
  wire[1:0] T1129;
  wire T1130;
  wire T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire T1135;
  wire[1:0] T1136;
  wire[1:0] T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[1:0] T1144;
  wire[1:0] T1145;
  wire T1146;
  wire T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire T1151;
  wire[1:0] T1152;
  wire[1:0] T1153;
  wire T1154;
  wire T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire T1159;
  wire[1:0] T1160;
  wire[1:0] T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire[1:0] T1168;
  wire[1:0] T1169;
  wire T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire[1:0] T1176;
  wire[1:0] T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire[1:0] T1184;
  wire[1:0] T1185;
  wire T1186;
  wire T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire T1191;
  wire[1:0] T1192;
  wire[1:0] T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire T1199;
  wire[1:0] T1200;
  wire[1:0] T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[1:0] T1208;
  wire[1:0] T1209;
  wire T1210;
  wire T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire T1215;
  wire[1:0] T1216;
  wire[1:0] T1217;
  wire T1218;
  wire T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire T1223;
  wire[1:0] T1224;
  wire[1:0] T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire[1:0] T1232;
  wire[1:0] T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire[1:0] T1240;
  wire[1:0] T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire[1:0] T1248;
  wire[1:0] T1249;
  wire T1250;
  wire T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire T1255;
  wire[1:0] T1256;
  wire[1:0] T1257;
  wire T1258;
  wire T1259;
  wire T1260;
  wire[3:0] T1261;
  wire[3:0] T1262;
  wire[3:0] T1263;
  wire[8:0] T1264;
  wire[8:0] T1265;
  wire T1266;
  wire T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire T1271;
  wire[1:0] T1272;
  wire[1:0] T1273;
  wire T1274;
  wire T1275;
  wire T1276;
  wire[3:0] T1277;
  wire[3:0] T1278;
  wire[3:0] T1279;
  wire[8:0] T1280;
  wire[8:0] T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[1:0] T1288;
  wire[1:0] T1289;
  wire T1290;
  wire T1291;
  wire T1292;
  wire[3:0] T1293;
  wire[3:0] T1294;
  wire[3:0] T1295;
  wire[8:0] T1296;
  wire[8:0] T1297;
  wire T1298;
  wire T1299;
  wire T1300;
  wire T1301;
  wire T1302;
  wire T1303;
  wire[1:0] T1304;
  wire[1:0] T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire[3:0] T1309;
  wire[3:0] T1310;
  wire[3:0] T1311;
  wire[8:0] T1312;
  wire[8:0] T1313;
  wire T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire[1:0] T1320;
  wire[1:0] T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire[3:0] T1325;
  wire[3:0] T1326;
  wire[3:0] T1327;
  wire[8:0] T1328;
  wire[8:0] T1329;
  wire T1330;
  wire T1331;
  wire T1332;
  wire T1333;
  wire T1334;
  wire T1335;
  wire[1:0] T1336;
  wire[1:0] T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire[3:0] T1341;
  wire[3:0] T1342;
  wire[3:0] T1343;
  wire[8:0] T1344;
  wire[8:0] T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[1:0] T1352;
  wire[1:0] T1353;
  wire T1354;
  wire T1355;
  wire T1356;
  wire[3:0] T1357;
  wire[3:0] T1358;
  wire[3:0] T1359;
  wire[8:0] T1360;
  wire[8:0] T1361;
  wire T1362;
  wire T1363;
  wire T1364;
  wire T1365;
  wire T1366;
  wire T1367;
  wire[1:0] T1368;
  wire[1:0] T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire[3:0] T1373;
  wire[3:0] T1374;
  wire[3:0] T1375;
  wire[8:0] T1376;
  wire[8:0] T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire[1:0] T1384;
  wire[1:0] T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire[3:0] T1389;
  wire[3:0] T1390;
  wire[3:0] T1391;
  wire[8:0] T1392;
  wire[8:0] T1393;
  wire T1394;
  wire T1395;
  wire T1396;
  wire T1397;
  wire T1398;
  wire T1399;
  wire[1:0] T1400;
  wire[1:0] T1401;
  wire T1402;
  wire T1403;
  wire T1404;
  wire[3:0] T1405;
  wire[3:0] T1406;
  wire[3:0] T1407;
  wire[8:0] T1408;
  wire[8:0] T1409;
  wire T1410;
  wire T1411;
  wire T1412;
  wire T1413;
  wire T1414;
  wire T1415;
  wire[1:0] T1416;
  wire[1:0] T1417;
  wire T1418;
  wire T1419;
  wire T1420;
  wire[3:0] T1421;
  wire[3:0] T1422;
  wire[3:0] T1423;
  wire[8:0] T1424;
  wire[8:0] T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[1:0] T1432;
  wire[1:0] T1433;
  wire T1434;
  wire T1435;
  wire T1436;
  wire[3:0] T1437;
  wire[3:0] T1438;
  wire[3:0] T1439;
  wire[8:0] T1440;
  wire[8:0] T1441;
  wire T1442;
  wire T1443;
  wire T1444;
  wire T1445;
  wire T1446;
  wire T1447;
  wire[1:0] T1448;
  wire[1:0] T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire[3:0] T1453;
  wire[3:0] T1454;
  wire[3:0] T1455;
  wire[8:0] T1456;
  wire[8:0] T1457;
  wire T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire[1:0] T1464;
  wire[1:0] T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire[3:0] T1469;
  wire[3:0] T1470;
  wire[3:0] T1471;
  wire[8:0] T1472;
  wire[8:0] T1473;
  wire T1474;
  wire T1475;
  wire T1476;
  wire T1477;
  wire T1478;
  wire T1479;
  wire[1:0] T1480;
  wire[1:0] T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire[3:0] T1485;
  wire[3:0] T1486;
  wire[3:0] T1487;
  wire[8:0] T1488;
  wire[8:0] T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[1:0] T1496;
  wire[1:0] T1497;
  wire[22:0] T1498;
  wire[22:0] T1499;
  wire[21:0] T1500;
  wire[21:0] T1501;
  wire[20:0] T1502;
  wire[20:0] T1503;
  wire[19:0] T1504;
  wire[19:0] T1505;
  wire[18:0] T1506;
  wire[18:0] T1507;
  wire[17:0] T1508;
  wire[17:0] T1509;
  wire[16:0] T1510;
  wire[16:0] T1511;
  wire[15:0] T1512;
  wire[15:0] T1513;
  wire[14:0] T1514;
  wire[14:0] T1515;
  wire[13:0] T1516;
  wire[13:0] T1517;
  wire[12:0] T1518;
  wire[12:0] T1519;
  wire[11:0] T1520;
  wire[11:0] T1521;
  wire[10:0] T1522;
  wire[10:0] T1523;
  wire[9:0] T1524;
  wire[9:0] T1525;
  wire[8:0] T1526;
  wire[8:0] T1527;
  wire[7:0] T1528;
  wire[7:0] T1529;
  wire[6:0] T1530;
  wire[6:0] T1531;
  wire[5:0] T1532;
  wire[5:0] T1533;
  wire[4:0] T1534;
  wire[4:0] T1535;
  wire[3:0] T1536;
  wire[3:0] T1537;
  wire[2:0] T1538;
  wire[2:0] T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[11:0] T1548;
  wire[11:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[11:0] T1556;
  wire[11:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[11:0] T1564;
  wire[11:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[11:0] T1572;
  wire[11:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[11:0] T1580;
  wire[11:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[11:0] T1588;
  wire[11:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[11:0] T1596;
  wire[11:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[11:0] T1604;
  wire[11:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[11:0] T1612;
  wire[11:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[11:0] T1620;
  wire[11:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[11:0] T1628;
  wire[11:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[11:0] T1636;
  wire[11:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[11:0] T1644;
  wire[11:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[11:0] T1652;
  wire[11:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[11:0] T1660;
  wire[11:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[11:0] T1668;
  wire[11:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[11:0] T1676;
  wire[11:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[11:0] T1684;
  wire[11:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[11:0] T1692;
  wire[11:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[11:0] T1700;
  wire[11:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[11:0] T1708;
  wire[11:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[11:0] T1716;
  wire[11:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[11:0] T1724;
  wire[11:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1490, T2};
  assign T2 = T3;
  assign T3 = {T1482, T4};
  assign T4 = T5;
  assign T5 = {T1474, T6};
  assign T6 = T7;
  assign T7 = {T1466, T8};
  assign T8 = T9;
  assign T9 = {T1458, T10};
  assign T10 = T11;
  assign T11 = {T1450, T12};
  assign T12 = T13;
  assign T13 = {T1442, T14};
  assign T14 = T15;
  assign T15 = {T1434, T16};
  assign T16 = T17;
  assign T17 = {T1426, T18};
  assign T18 = T19;
  assign T19 = {T1418, T20};
  assign T20 = T21;
  assign T21 = {T1410, T22};
  assign T22 = T23;
  assign T23 = {T1402, T24};
  assign T24 = T25;
  assign T25 = {T1394, T26};
  assign T26 = T27;
  assign T27 = {T1386, T28};
  assign T28 = T29;
  assign T29 = {T1378, T30};
  assign T30 = T31;
  assign T31 = {T1370, T32};
  assign T32 = T33;
  assign T33 = {T1362, T34};
  assign T34 = T35;
  assign T35 = {T1354, T36};
  assign T36 = T37;
  assign T37 = {T1346, T38};
  assign T38 = T39;
  assign T39 = {T1338, T40};
  assign T40 = T41;
  assign T41 = {T1330, T42};
  assign T42 = T43;
  assign T43 = {T1322, T44};
  assign T44 = T45;
  assign T45 = {T1314, T46};
  assign T46 = T47;
  assign T47 = {T1306, T48};
  assign T48 = T49;
  assign T49 = {T1298, T50};
  assign T50 = T51;
  assign T51 = {T1290, T52};
  assign T52 = T53;
  assign T53 = {T1282, T54};
  assign T54 = T55;
  assign T55 = {T1274, T56};
  assign T56 = T57;
  assign T57 = {T1266, T58};
  assign T58 = T59;
  assign T59 = {T1258, T60};
  assign T60 = T61;
  assign T61 = {T1250, T62};
  assign T62 = T63;
  assign T63 = {T1242, T64};
  assign T64 = T65;
  assign T65 = {T1234, T66};
  assign T66 = T67;
  assign T67 = {T1226, T68};
  assign T68 = T69;
  assign T69 = {T1218, T70};
  assign T70 = T71;
  assign T71 = {T1210, T72};
  assign T72 = T73;
  assign T73 = {T1202, T74};
  assign T74 = T75;
  assign T75 = {T1194, T76};
  assign T76 = T77;
  assign T77 = {T1186, T78};
  assign T78 = T79;
  assign T79 = {T1178, T80};
  assign T80 = T81;
  assign T81 = {T1170, T82};
  assign T82 = T83;
  assign T83 = {T1162, T84};
  assign T84 = T85;
  assign T85 = {T1154, T86};
  assign T86 = T87;
  assign T87 = {T1146, T88};
  assign T88 = T89;
  assign T89 = {T1138, T90};
  assign T90 = T91;
  assign T91 = {T1130, T92};
  assign T92 = T93;
  assign T93 = {T1122, T94};
  assign T94 = T95;
  assign T95 = {T1114, T96};
  assign T96 = T97;
  assign T97 = {T1106, T98};
  assign T98 = T99;
  assign T99 = {T1098, T100};
  assign T100 = T101;
  assign T101 = {T1090, T102};
  assign T102 = T103;
  assign T103 = {T1082, T104};
  assign T104 = T105;
  assign T105 = {T1074, T106};
  assign T106 = T107;
  assign T107 = {T1066, T108};
  assign T108 = T109;
  assign T109 = {T1058, T110};
  assign T110 = T111;
  assign T111 = {T1050, T112};
  assign T112 = T113;
  assign T113 = {T1042, T114};
  assign T114 = T115;
  assign T115 = {T1034, T116};
  assign T116 = T117;
  assign T117 = {T1026, T118};
  assign T118 = T119;
  assign T119 = {T1018, T120};
  assign T120 = T121;
  assign T121 = {T1010, T122};
  assign T122 = T123;
  assign T123 = {T1002, T124};
  assign T124 = T125;
  assign T125 = {T994, T126};
  assign T126 = T127;
  assign T127 = {T986, T128};
  assign T128 = T129;
  assign T129 = {T978, T130};
  assign T130 = T131;
  assign T131 = {T970, T132};
  assign T132 = T133;
  assign T133 = {T962, T134};
  assign T134 = T135;
  assign T135 = {T954, T136};
  assign T136 = T137;
  assign T137 = {T946, T138};
  assign T138 = T139;
  assign T139 = {T938, T140};
  assign T140 = T141;
  assign T141 = {T930, T142};
  assign T142 = T143;
  assign T143 = {T922, T144};
  assign T144 = T145;
  assign T145 = {T914, T146};
  assign T146 = T147;
  assign T147 = {T906, T148};
  assign T148 = T149;
  assign T149 = {T898, T150};
  assign T150 = T151;
  assign T151 = {T890, T152};
  assign T152 = T153;
  assign T153 = {T882, T154};
  assign T154 = T155;
  assign T155 = {T874, T156};
  assign T156 = T157;
  assign T157 = {T866, T158};
  assign T158 = T159;
  assign T159 = {T858, T160};
  assign T160 = T161;
  assign T161 = {T850, T162};
  assign T162 = T163;
  assign T163 = {T842, T164};
  assign T164 = T165;
  assign T165 = {T834, T166};
  assign T166 = T167;
  assign T167 = {T826, T168};
  assign T168 = T169;
  assign T169 = {T818, T170};
  assign T170 = T171;
  assign T171 = {T810, T172};
  assign T172 = T173;
  assign T173 = {T802, T174};
  assign T174 = T175;
  assign T175 = {T794, T176};
  assign T176 = T177;
  assign T177 = {T786, T178};
  assign T178 = T179;
  assign T179 = {T778, T180};
  assign T180 = T181;
  assign T181 = {T770, T182};
  assign T182 = T183;
  assign T183 = {T762, T184};
  assign T184 = T185;
  assign T185 = {T754, T186};
  assign T186 = T187;
  assign T187 = {T746, T188};
  assign T188 = T189;
  assign T189 = {T738, T190};
  assign T190 = T191;
  assign T191 = {T730, T192};
  assign T192 = T193;
  assign T193 = {T722, T194};
  assign T194 = T195;
  assign T195 = {T714, T196};
  assign T196 = T197;
  assign T197 = {T706, T198};
  assign T198 = T199;
  assign T199 = {T698, T200};
  assign T200 = T201;
  assign T201 = {T690, T202};
  assign T202 = T203;
  assign T203 = {T682, T204};
  assign T204 = T205;
  assign T205 = {T674, T206};
  assign T206 = T207;
  assign T207 = {T666, T208};
  assign T208 = T209;
  assign T209 = {T658, T210};
  assign T210 = T211;
  assign T211 = {T650, T212};
  assign T212 = T213;
  assign T213 = {T642, T214};
  assign T214 = T215;
  assign T215 = {T634, T216};
  assign T216 = T217;
  assign T217 = {T626, T218};
  assign T218 = T219;
  assign T219 = {T618, T220};
  assign T220 = T221;
  assign T221 = {T610, T222};
  assign T222 = T223;
  assign T223 = {T602, T224};
  assign T224 = T225;
  assign T225 = {T594, T226};
  assign T226 = T227;
  assign T227 = {T586, T228};
  assign T228 = T229;
  assign T229 = {T578, T230};
  assign T230 = T231;
  assign T231 = {T570, T232};
  assign T232 = T233;
  assign T233 = {T562, T234};
  assign T234 = T235;
  assign T235 = {T554, T236};
  assign T236 = T237;
  assign T237 = {T546, T238};
  assign T238 = T239;
  assign T239 = {T538, T240};
  assign T240 = T241;
  assign T241 = {T530, T242};
  assign T242 = T243;
  assign T243 = {T522, T244};
  assign T244 = T245;
  assign T245 = {T514, T246};
  assign T246 = T247;
  assign T247 = {T506, T248};
  assign T248 = T249;
  assign T249 = {T498, T250};
  assign T250 = T251;
  assign T251 = {T490, T252};
  assign T252 = T253;
  assign T253 = {T482, T254};
  assign T254 = T255;
  assign T255 = {T474, T256};
  assign T256 = T257;
  assign T257 = {T466, T258};
  assign T258 = T259;
  assign T259 = {T458, T260};
  assign T260 = T261;
  assign T261 = {T450, T262};
  assign T262 = T263;
  assign T263 = {T442, T264};
  assign T264 = T265;
  assign T265 = {T434, T266};
  assign T266 = T267;
  assign T267 = {T426, T268};
  assign T268 = T269;
  assign T269 = {T418, T270};
  assign T270 = T271;
  assign T271 = {T410, T272};
  assign T272 = T273;
  assign T273 = {T402, T274};
  assign T274 = T275;
  assign T275 = {T394, T276};
  assign T276 = T277;
  assign T277 = {T386, T278};
  assign T278 = T279;
  assign T279 = {T378, T280};
  assign T280 = T281;
  assign T281 = {T370, T282};
  assign T282 = T283;
  assign T283 = {T362, T284};
  assign T284 = T285;
  assign T285 = {T354, T286};
  assign T286 = T287;
  assign T287 = {T346, T288};
  assign T288 = T289;
  assign T289 = {T338, T290};
  assign T290 = T291;
  assign T291 = {T330, T292};
  assign T292 = T293;
  assign T293 = {T322, T294};
  assign T294 = T295;
  assign T295 = {T314, T296};
  assign T296 = T297;
  assign T297 = {T306, T298};
  assign T298 = T299;
  assign T299 = T300;
  assign T300 = T304[T301];
  assign T301 = T302;
  assign T302 = T303;
  assign T303 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T304 = T305;
  assign T305 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T306 = T307;
  assign T307 = T308;
  assign T308 = T312[T309];
  assign T309 = T310;
  assign T310 = T311;
  assign T311 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T312 = T313;
  assign T313 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T314 = T315;
  assign T315 = T316;
  assign T316 = T320[T317];
  assign T317 = T318;
  assign T318 = T319;
  assign T319 = io_chanxy_config[2'h2/* 2*/:2'h2/* 2*/];
  assign T320 = T321;
  assign T321 = io_chanxy_in[3'h5/* 5*/:3'h4/* 4*/];
  assign T322 = T323;
  assign T323 = T324;
  assign T324 = T328[T325];
  assign T325 = T326;
  assign T326 = T327;
  assign T327 = io_chanxy_config[2'h3/* 3*/:2'h3/* 3*/];
  assign T328 = T329;
  assign T329 = io_chanxy_in[3'h7/* 7*/:3'h6/* 6*/];
  assign T330 = T331;
  assign T331 = T332;
  assign T332 = T336[T333];
  assign T333 = T334;
  assign T334 = T335;
  assign T335 = io_chanxy_config[3'h4/* 4*/:3'h4/* 4*/];
  assign T336 = T337;
  assign T337 = io_chanxy_in[4'h9/* 9*/:4'h8/* 8*/];
  assign T338 = T339;
  assign T339 = T340;
  assign T340 = T344[T341];
  assign T341 = T342;
  assign T342 = T343;
  assign T343 = io_chanxy_config[3'h5/* 5*/:3'h5/* 5*/];
  assign T344 = T345;
  assign T345 = io_chanxy_in[4'hb/* 11*/:4'ha/* 10*/];
  assign T346 = T347;
  assign T347 = T348;
  assign T348 = T352[T349];
  assign T349 = T350;
  assign T350 = T351;
  assign T351 = io_chanxy_config[3'h6/* 6*/:3'h6/* 6*/];
  assign T352 = T353;
  assign T353 = io_chanxy_in[4'hd/* 13*/:4'hc/* 12*/];
  assign T354 = T355;
  assign T355 = T356;
  assign T356 = T360[T357];
  assign T357 = T358;
  assign T358 = T359;
  assign T359 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T360 = T361;
  assign T361 = io_chanxy_in[4'hf/* 15*/:4'he/* 14*/];
  assign T362 = T363;
  assign T363 = T364;
  assign T364 = T368[T365];
  assign T365 = T366;
  assign T366 = T367;
  assign T367 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T368 = T369;
  assign T369 = io_chanxy_in[5'h11/* 17*/:5'h10/* 16*/];
  assign T370 = T371;
  assign T371 = T372;
  assign T372 = T376[T373];
  assign T373 = T374;
  assign T374 = T375;
  assign T375 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T376 = T377;
  assign T377 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T378 = T379;
  assign T379 = T380;
  assign T380 = T384[T381];
  assign T381 = T382;
  assign T382 = T383;
  assign T383 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T384 = T385;
  assign T385 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T386 = T387;
  assign T387 = T388;
  assign T388 = T392[T389];
  assign T389 = T390;
  assign T390 = T391;
  assign T391 = io_chanxy_config[4'hb/* 11*/:4'hb/* 11*/];
  assign T392 = T393;
  assign T393 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T394 = T395;
  assign T395 = T396;
  assign T396 = T400[T397];
  assign T397 = T398;
  assign T398 = T399;
  assign T399 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T400 = T401;
  assign T401 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T402 = T403;
  assign T403 = T404;
  assign T404 = T408[T405];
  assign T405 = T406;
  assign T406 = T407;
  assign T407 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T408 = T409;
  assign T409 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T410 = T411;
  assign T411 = T412;
  assign T412 = T416[T413];
  assign T413 = T414;
  assign T414 = T415;
  assign T415 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T416 = T417;
  assign T417 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T418 = T419;
  assign T419 = T420;
  assign T420 = T424[T421];
  assign T421 = T422;
  assign T422 = T423;
  assign T423 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T424 = T425;
  assign T425 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T426 = T427;
  assign T427 = T428;
  assign T428 = T432[T429];
  assign T429 = T430;
  assign T430 = T431;
  assign T431 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T432 = T433;
  assign T433 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T434 = T435;
  assign T435 = T436;
  assign T436 = T440[T437];
  assign T437 = T438;
  assign T438 = T439;
  assign T439 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T440 = T441;
  assign T441 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T442 = T443;
  assign T443 = T444;
  assign T444 = T448[T445];
  assign T445 = T446;
  assign T446 = T447;
  assign T447 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T448 = T449;
  assign T449 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T450 = T451;
  assign T451 = T452;
  assign T452 = T456[T453];
  assign T453 = T454;
  assign T454 = T455;
  assign T455 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T456 = T457;
  assign T457 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T458 = T459;
  assign T459 = T460;
  assign T460 = T464[T461];
  assign T461 = T462;
  assign T462 = T463;
  assign T463 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T464 = T465;
  assign T465 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T466 = T467;
  assign T467 = T468;
  assign T468 = T472[T469];
  assign T469 = T470;
  assign T470 = T471;
  assign T471 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T472 = T473;
  assign T473 = io_chanxy_in[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T474 = T475;
  assign T475 = T476;
  assign T476 = T480[T477];
  assign T477 = T478;
  assign T478 = T479;
  assign T479 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T480 = T481;
  assign T481 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T482 = T483;
  assign T483 = T484;
  assign T484 = T488[T485];
  assign T485 = T486;
  assign T486 = T487;
  assign T487 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T488 = T489;
  assign T489 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T490 = T491;
  assign T491 = T492;
  assign T492 = T496[T493];
  assign T493 = T494;
  assign T494 = T495;
  assign T495 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T496 = T497;
  assign T497 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T498 = T499;
  assign T499 = T500;
  assign T500 = T504[T501];
  assign T501 = T502;
  assign T502 = T503;
  assign T503 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T504 = T505;
  assign T505 = io_chanxy_in[6'h33/* 51*/:6'h32/* 50*/];
  assign T506 = T507;
  assign T507 = T508;
  assign T508 = T512[T509];
  assign T509 = T510;
  assign T510 = T511;
  assign T511 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T512 = T513;
  assign T513 = io_chanxy_in[6'h35/* 53*/:6'h34/* 52*/];
  assign T514 = T515;
  assign T515 = T516;
  assign T516 = T520[T517];
  assign T517 = T518;
  assign T518 = T519;
  assign T519 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T520 = T521;
  assign T521 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T522 = T523;
  assign T523 = T524;
  assign T524 = T528[T525];
  assign T525 = T526;
  assign T526 = T527;
  assign T527 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T528 = T529;
  assign T529 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T530 = T531;
  assign T531 = T532;
  assign T532 = T536[T533];
  assign T533 = T534;
  assign T534 = T535;
  assign T535 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T536 = T537;
  assign T537 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T538 = T539;
  assign T539 = T540;
  assign T540 = T544[T541];
  assign T541 = T542;
  assign T542 = T543;
  assign T543 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T544 = T545;
  assign T545 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T546 = T547;
  assign T547 = T548;
  assign T548 = T552[T549];
  assign T549 = T550;
  assign T550 = T551;
  assign T551 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T552 = T553;
  assign T553 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T554 = T555;
  assign T555 = T556;
  assign T556 = T560[T557];
  assign T557 = T558;
  assign T558 = T559;
  assign T559 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T560 = T561;
  assign T561 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T562 = T563;
  assign T563 = T564;
  assign T564 = T568[T565];
  assign T565 = T566;
  assign T566 = T567;
  assign T567 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T568 = T569;
  assign T569 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T570 = T571;
  assign T571 = T572;
  assign T572 = T576[T573];
  assign T573 = T574;
  assign T574 = T575;
  assign T575 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T576 = T577;
  assign T577 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T578 = T579;
  assign T579 = T580;
  assign T580 = T584[T581];
  assign T581 = T582;
  assign T582 = T583;
  assign T583 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T584 = T585;
  assign T585 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T586 = T587;
  assign T587 = T588;
  assign T588 = T592[T589];
  assign T589 = T590;
  assign T590 = T591;
  assign T591 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T592 = T593;
  assign T593 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T594 = T595;
  assign T595 = T596;
  assign T596 = T600[T597];
  assign T597 = T598;
  assign T598 = T599;
  assign T599 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T600 = T601;
  assign T601 = io_chanxy_in[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T602 = T603;
  assign T603 = T604;
  assign T604 = T608[T605];
  assign T605 = T606;
  assign T606 = T607;
  assign T607 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T608 = T609;
  assign T609 = io_chanxy_in[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T610 = T611;
  assign T611 = T612;
  assign T612 = T616[T613];
  assign T613 = T614;
  assign T614 = T615;
  assign T615 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T616 = T617;
  assign T617 = io_chanxy_in[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T618 = T619;
  assign T619 = T620;
  assign T620 = T624[T621];
  assign T621 = T622;
  assign T622 = T623;
  assign T623 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T624 = T625;
  assign T625 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T626 = T627;
  assign T627 = T628;
  assign T628 = T632[T629];
  assign T629 = T630;
  assign T630 = T631;
  assign T631 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T632 = T633;
  assign T633 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T634 = T635;
  assign T635 = T636;
  assign T636 = T640[T637];
  assign T637 = T638;
  assign T638 = T639;
  assign T639 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T640 = T641;
  assign T641 = io_chanxy_in[7'h55/* 85*/:7'h54/* 84*/];
  assign T642 = T643;
  assign T643 = T644;
  assign T644 = T648[T645];
  assign T645 = T646;
  assign T646 = T647;
  assign T647 = io_chanxy_config[6'h2b/* 43*/:6'h2b/* 43*/];
  assign T648 = T649;
  assign T649 = io_chanxy_in[7'h57/* 87*/:7'h56/* 86*/];
  assign T650 = T651;
  assign T651 = T652;
  assign T652 = T656[T653];
  assign T653 = T654;
  assign T654 = T655;
  assign T655 = io_chanxy_config[6'h2c/* 44*/:6'h2c/* 44*/];
  assign T656 = T657;
  assign T657 = io_chanxy_in[7'h59/* 89*/:7'h58/* 88*/];
  assign T658 = T659;
  assign T659 = T660;
  assign T660 = T664[T661];
  assign T661 = T662;
  assign T662 = T663;
  assign T663 = io_chanxy_config[6'h30/* 48*/:6'h2d/* 45*/];
  assign T664 = T665;
  assign T665 = io_chanxy_in[7'h62/* 98*/:7'h5a/* 90*/];
  assign T666 = T667;
  assign T667 = T668;
  assign T668 = T672[T669];
  assign T669 = T670;
  assign T670 = T671;
  assign T671 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T672 = T673;
  assign T673 = io_chanxy_in[7'h64/* 100*/:7'h63/* 99*/];
  assign T674 = T675;
  assign T675 = T676;
  assign T676 = T680[T677];
  assign T677 = T678;
  assign T678 = T679;
  assign T679 = io_chanxy_config[6'h35/* 53*/:6'h32/* 50*/];
  assign T680 = T681;
  assign T681 = io_chanxy_in[7'h6d/* 109*/:7'h65/* 101*/];
  assign T682 = T683;
  assign T683 = T684;
  assign T684 = T688[T685];
  assign T685 = T686;
  assign T686 = T687;
  assign T687 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T688 = T689;
  assign T689 = io_chanxy_in[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T690 = T691;
  assign T691 = T692;
  assign T692 = T696[T693];
  assign T693 = T694;
  assign T694 = T695;
  assign T695 = io_chanxy_config[6'h3a/* 58*/:6'h37/* 55*/];
  assign T696 = T697;
  assign T697 = io_chanxy_in[7'h78/* 120*/:7'h70/* 112*/];
  assign T698 = T699;
  assign T699 = T700;
  assign T700 = T704[T701];
  assign T701 = T702;
  assign T702 = T703;
  assign T703 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T704 = T705;
  assign T705 = io_chanxy_in[7'h7a/* 122*/:7'h79/* 121*/];
  assign T706 = T707;
  assign T707 = T708;
  assign T708 = T712[T709];
  assign T709 = T710;
  assign T710 = T711;
  assign T711 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T712 = T713;
  assign T713 = io_chanxy_in[8'h83/* 131*/:7'h7b/* 123*/];
  assign T714 = T715;
  assign T715 = T716;
  assign T716 = T720[T717];
  assign T717 = T718;
  assign T718 = T719;
  assign T719 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T720 = T721;
  assign T721 = io_chanxy_in[8'h85/* 133*/:8'h84/* 132*/];
  assign T722 = T723;
  assign T723 = T724;
  assign T724 = T728[T725];
  assign T725 = T726;
  assign T726 = T727;
  assign T727 = io_chanxy_config[7'h44/* 68*/:7'h41/* 65*/];
  assign T728 = T729;
  assign T729 = io_chanxy_in[8'h8e/* 142*/:8'h86/* 134*/];
  assign T730 = T731;
  assign T731 = T732;
  assign T732 = T736[T733];
  assign T733 = T734;
  assign T734 = T735;
  assign T735 = io_chanxy_config[7'h45/* 69*/:7'h45/* 69*/];
  assign T736 = T737;
  assign T737 = io_chanxy_in[8'h90/* 144*/:8'h8f/* 143*/];
  assign T738 = T739;
  assign T739 = T740;
  assign T740 = T744[T741];
  assign T741 = T742;
  assign T742 = T743;
  assign T743 = io_chanxy_config[7'h49/* 73*/:7'h46/* 70*/];
  assign T744 = T745;
  assign T745 = io_chanxy_in[8'h99/* 153*/:8'h91/* 145*/];
  assign T746 = T747;
  assign T747 = T748;
  assign T748 = T752[T749];
  assign T749 = T750;
  assign T750 = T751;
  assign T751 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T752 = T753;
  assign T753 = io_chanxy_in[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T754 = T755;
  assign T755 = T756;
  assign T756 = T760[T757];
  assign T757 = T758;
  assign T758 = T759;
  assign T759 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T760 = T761;
  assign T761 = io_chanxy_in[8'ha4/* 164*/:8'h9c/* 156*/];
  assign T762 = T763;
  assign T763 = T764;
  assign T764 = T768[T765];
  assign T765 = T766;
  assign T766 = T767;
  assign T767 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T768 = T769;
  assign T769 = io_chanxy_in[8'ha6/* 166*/:8'ha5/* 165*/];
  assign T770 = T771;
  assign T771 = T772;
  assign T772 = T776[T773];
  assign T773 = T774;
  assign T774 = T775;
  assign T775 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T776 = T777;
  assign T777 = io_chanxy_in[8'haf/* 175*/:8'ha7/* 167*/];
  assign T778 = T779;
  assign T779 = T780;
  assign T780 = T784[T781];
  assign T781 = T782;
  assign T782 = T783;
  assign T783 = io_chanxy_config[7'h54/* 84*/:7'h54/* 84*/];
  assign T784 = T785;
  assign T785 = io_chanxy_in[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T786 = T787;
  assign T787 = T788;
  assign T788 = T792[T789];
  assign T789 = T790;
  assign T790 = T791;
  assign T791 = io_chanxy_config[7'h58/* 88*/:7'h55/* 85*/];
  assign T792 = T793;
  assign T793 = io_chanxy_in[8'hba/* 186*/:8'hb2/* 178*/];
  assign T794 = T795;
  assign T795 = T796;
  assign T796 = T800[T797];
  assign T797 = T798;
  assign T798 = T799;
  assign T799 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T800 = T801;
  assign T801 = io_chanxy_in[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T802 = T803;
  assign T803 = T804;
  assign T804 = T808[T805];
  assign T805 = T806;
  assign T806 = T807;
  assign T807 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T808 = T809;
  assign T809 = io_chanxy_in[8'hc5/* 197*/:8'hbd/* 189*/];
  assign T810 = T811;
  assign T811 = T812;
  assign T812 = T816[T813];
  assign T813 = T814;
  assign T814 = T815;
  assign T815 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T816 = T817;
  assign T817 = io_chanxy_in[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T818 = T819;
  assign T819 = T820;
  assign T820 = T824[T821];
  assign T821 = T822;
  assign T822 = T823;
  assign T823 = io_chanxy_config[7'h62/* 98*/:7'h5f/* 95*/];
  assign T824 = T825;
  assign T825 = io_chanxy_in[8'hd0/* 208*/:8'hc8/* 200*/];
  assign T826 = T827;
  assign T827 = T828;
  assign T828 = T832[T829];
  assign T829 = T830;
  assign T830 = T831;
  assign T831 = io_chanxy_config[7'h63/* 99*/:7'h63/* 99*/];
  assign T832 = T833;
  assign T833 = io_chanxy_in[8'hd2/* 210*/:8'hd1/* 209*/];
  assign T834 = T835;
  assign T835 = T836;
  assign T836 = T840[T837];
  assign T837 = T838;
  assign T838 = T839;
  assign T839 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T840 = T841;
  assign T841 = io_chanxy_in[8'hdb/* 219*/:8'hd3/* 211*/];
  assign T842 = T843;
  assign T843 = T844;
  assign T844 = T848[T845];
  assign T845 = T846;
  assign T846 = T847;
  assign T847 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T848 = T849;
  assign T849 = io_chanxy_in[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T850 = T851;
  assign T851 = T852;
  assign T852 = T856[T853];
  assign T853 = T854;
  assign T854 = T855;
  assign T855 = io_chanxy_config[7'h6c/* 108*/:7'h69/* 105*/];
  assign T856 = T857;
  assign T857 = io_chanxy_in[8'he6/* 230*/:8'hde/* 222*/];
  assign T858 = T859;
  assign T859 = T860;
  assign T860 = T864[T861];
  assign T861 = T862;
  assign T862 = T863;
  assign T863 = io_chanxy_config[7'h6d/* 109*/:7'h6d/* 109*/];
  assign T864 = T865;
  assign T865 = io_chanxy_in[8'he8/* 232*/:8'he7/* 231*/];
  assign T866 = T867;
  assign T867 = T868;
  assign T868 = T872[T869];
  assign T869 = T870;
  assign T870 = T871;
  assign T871 = io_chanxy_config[7'h71/* 113*/:7'h6e/* 110*/];
  assign T872 = T873;
  assign T873 = io_chanxy_in[8'hf1/* 241*/:8'he9/* 233*/];
  assign T874 = T875;
  assign T875 = T876;
  assign T876 = T880[T877];
  assign T877 = T878;
  assign T878 = T879;
  assign T879 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T880 = T881;
  assign T881 = io_chanxy_in[8'hf3/* 243*/:8'hf2/* 242*/];
  assign T882 = T883;
  assign T883 = T884;
  assign T884 = T888[T885];
  assign T885 = T886;
  assign T886 = T887;
  assign T887 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T888 = T889;
  assign T889 = io_chanxy_in[8'hfc/* 252*/:8'hf4/* 244*/];
  assign T890 = T891;
  assign T891 = T892;
  assign T892 = T896[T893];
  assign T893 = T894;
  assign T894 = T895;
  assign T895 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T896 = T897;
  assign T897 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T898 = T899;
  assign T899 = T900;
  assign T900 = T904[T901];
  assign T901 = T902;
  assign T902 = T903;
  assign T903 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T904 = T905;
  assign T905 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T906 = T907;
  assign T907 = T908;
  assign T908 = T912[T909];
  assign T909 = T910;
  assign T910 = T911;
  assign T911 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T912 = T913;
  assign T913 = io_chanxy_in[9'h102/* 258*/:9'h101/* 257*/];
  assign T914 = T915;
  assign T915 = T916;
  assign T916 = T920[T917];
  assign T917 = T918;
  assign T918 = T919;
  assign T919 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T920 = T921;
  assign T921 = io_chanxy_in[9'h104/* 260*/:9'h103/* 259*/];
  assign T922 = T923;
  assign T923 = T924;
  assign T924 = T928[T925];
  assign T925 = T926;
  assign T926 = T927;
  assign T927 = io_chanxy_config[7'h7b/* 123*/:7'h7b/* 123*/];
  assign T928 = T929;
  assign T929 = io_chanxy_in[9'h106/* 262*/:9'h105/* 261*/];
  assign T930 = T931;
  assign T931 = T932;
  assign T932 = T936[T933];
  assign T933 = T934;
  assign T934 = T935;
  assign T935 = io_chanxy_config[7'h7c/* 124*/:7'h7c/* 124*/];
  assign T936 = T937;
  assign T937 = io_chanxy_in[9'h108/* 264*/:9'h107/* 263*/];
  assign T938 = T939;
  assign T939 = T940;
  assign T940 = T944[T941];
  assign T941 = T942;
  assign T942 = T943;
  assign T943 = io_chanxy_config[7'h7d/* 125*/:7'h7d/* 125*/];
  assign T944 = T945;
  assign T945 = io_chanxy_in[9'h10a/* 266*/:9'h109/* 265*/];
  assign T946 = T947;
  assign T947 = T948;
  assign T948 = T952[T949];
  assign T949 = T950;
  assign T950 = T951;
  assign T951 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T952 = T953;
  assign T953 = io_chanxy_in[9'h10c/* 268*/:9'h10b/* 267*/];
  assign T954 = T955;
  assign T955 = T956;
  assign T956 = T960[T957];
  assign T957 = T958;
  assign T958 = T959;
  assign T959 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T960 = T961;
  assign T961 = io_chanxy_in[9'h10e/* 270*/:9'h10d/* 269*/];
  assign T962 = T963;
  assign T963 = T964;
  assign T964 = T968[T965];
  assign T965 = T966;
  assign T966 = T967;
  assign T967 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T968 = T969;
  assign T969 = io_chanxy_in[9'h110/* 272*/:9'h10f/* 271*/];
  assign T970 = T971;
  assign T971 = T972;
  assign T972 = T976[T973];
  assign T973 = T974;
  assign T974 = T975;
  assign T975 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T976 = T977;
  assign T977 = io_chanxy_in[9'h112/* 274*/:9'h111/* 273*/];
  assign T978 = T979;
  assign T979 = T980;
  assign T980 = T984[T981];
  assign T981 = T982;
  assign T982 = T983;
  assign T983 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T984 = T985;
  assign T985 = io_chanxy_in[9'h114/* 276*/:9'h113/* 275*/];
  assign T986 = T987;
  assign T987 = T988;
  assign T988 = T992[T989];
  assign T989 = T990;
  assign T990 = T991;
  assign T991 = io_chanxy_config[8'h83/* 131*/:8'h83/* 131*/];
  assign T992 = T993;
  assign T993 = io_chanxy_in[9'h116/* 278*/:9'h115/* 277*/];
  assign T994 = T995;
  assign T995 = T996;
  assign T996 = T1000[T997];
  assign T997 = T998;
  assign T998 = T999;
  assign T999 = io_chanxy_config[8'h84/* 132*/:8'h84/* 132*/];
  assign T1000 = T1001;
  assign T1001 = io_chanxy_in[9'h118/* 280*/:9'h117/* 279*/];
  assign T1002 = T1003;
  assign T1003 = T1004;
  assign T1004 = T1008[T1005];
  assign T1005 = T1006;
  assign T1006 = T1007;
  assign T1007 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T1008 = T1009;
  assign T1009 = io_chanxy_in[9'h11a/* 282*/:9'h119/* 281*/];
  assign T1010 = T1011;
  assign T1011 = T1012;
  assign T1012 = T1016[T1013];
  assign T1013 = T1014;
  assign T1014 = T1015;
  assign T1015 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T1016 = T1017;
  assign T1017 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T1018 = T1019;
  assign T1019 = T1020;
  assign T1020 = T1024[T1021];
  assign T1021 = T1022;
  assign T1022 = T1023;
  assign T1023 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T1024 = T1025;
  assign T1025 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T1026 = T1027;
  assign T1027 = T1028;
  assign T1028 = T1032[T1029];
  assign T1029 = T1030;
  assign T1030 = T1031;
  assign T1031 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T1032 = T1033;
  assign T1033 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T1034 = T1035;
  assign T1035 = T1036;
  assign T1036 = T1040[T1037];
  assign T1037 = T1038;
  assign T1038 = T1039;
  assign T1039 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T1040 = T1041;
  assign T1041 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T1042 = T1043;
  assign T1043 = T1044;
  assign T1044 = T1048[T1045];
  assign T1045 = T1046;
  assign T1046 = T1047;
  assign T1047 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T1048 = T1049;
  assign T1049 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T1050 = T1051;
  assign T1051 = T1052;
  assign T1052 = T1056[T1053];
  assign T1053 = T1054;
  assign T1054 = T1055;
  assign T1055 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T1056 = T1057;
  assign T1057 = io_chanxy_in[9'h126/* 294*/:9'h125/* 293*/];
  assign T1058 = T1059;
  assign T1059 = T1060;
  assign T1060 = T1064[T1061];
  assign T1061 = T1062;
  assign T1062 = T1063;
  assign T1063 = io_chanxy_config[8'h8c/* 140*/:8'h8c/* 140*/];
  assign T1064 = T1065;
  assign T1065 = io_chanxy_in[9'h128/* 296*/:9'h127/* 295*/];
  assign T1066 = T1067;
  assign T1067 = T1068;
  assign T1068 = T1072[T1069];
  assign T1069 = T1070;
  assign T1070 = T1071;
  assign T1071 = io_chanxy_config[8'h8d/* 141*/:8'h8d/* 141*/];
  assign T1072 = T1073;
  assign T1073 = io_chanxy_in[9'h12a/* 298*/:9'h129/* 297*/];
  assign T1074 = T1075;
  assign T1075 = T1076;
  assign T1076 = T1080[T1077];
  assign T1077 = T1078;
  assign T1078 = T1079;
  assign T1079 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T1080 = T1081;
  assign T1081 = io_chanxy_in[9'h12c/* 300*/:9'h12b/* 299*/];
  assign T1082 = T1083;
  assign T1083 = T1084;
  assign T1084 = T1088[T1085];
  assign T1085 = T1086;
  assign T1086 = T1087;
  assign T1087 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T1088 = T1089;
  assign T1089 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T1090 = T1091;
  assign T1091 = T1092;
  assign T1092 = T1096[T1093];
  assign T1093 = T1094;
  assign T1094 = T1095;
  assign T1095 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T1096 = T1097;
  assign T1097 = io_chanxy_in[9'h130/* 304*/:9'h12f/* 303*/];
  assign T1098 = T1099;
  assign T1099 = T1100;
  assign T1100 = T1104[T1101];
  assign T1101 = T1102;
  assign T1102 = T1103;
  assign T1103 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T1104 = T1105;
  assign T1105 = io_chanxy_in[9'h132/* 306*/:9'h131/* 305*/];
  assign T1106 = T1107;
  assign T1107 = T1108;
  assign T1108 = T1112[T1109];
  assign T1109 = T1110;
  assign T1110 = T1111;
  assign T1111 = io_chanxy_config[8'h92/* 146*/:8'h92/* 146*/];
  assign T1112 = T1113;
  assign T1113 = io_chanxy_in[9'h134/* 308*/:9'h133/* 307*/];
  assign T1114 = T1115;
  assign T1115 = T1116;
  assign T1116 = T1120[T1117];
  assign T1117 = T1118;
  assign T1118 = T1119;
  assign T1119 = io_chanxy_config[8'h93/* 147*/:8'h93/* 147*/];
  assign T1120 = T1121;
  assign T1121 = io_chanxy_in[9'h136/* 310*/:9'h135/* 309*/];
  assign T1122 = T1123;
  assign T1123 = T1124;
  assign T1124 = T1128[T1125];
  assign T1125 = T1126;
  assign T1126 = T1127;
  assign T1127 = io_chanxy_config[8'h94/* 148*/:8'h94/* 148*/];
  assign T1128 = T1129;
  assign T1129 = io_chanxy_in[9'h138/* 312*/:9'h137/* 311*/];
  assign T1130 = T1131;
  assign T1131 = T1132;
  assign T1132 = T1136[T1133];
  assign T1133 = T1134;
  assign T1134 = T1135;
  assign T1135 = io_chanxy_config[8'h95/* 149*/:8'h95/* 149*/];
  assign T1136 = T1137;
  assign T1137 = io_chanxy_in[9'h13a/* 314*/:9'h139/* 313*/];
  assign T1138 = T1139;
  assign T1139 = T1140;
  assign T1140 = T1144[T1141];
  assign T1141 = T1142;
  assign T1142 = T1143;
  assign T1143 = io_chanxy_config[8'h96/* 150*/:8'h96/* 150*/];
  assign T1144 = T1145;
  assign T1145 = io_chanxy_in[9'h13c/* 316*/:9'h13b/* 315*/];
  assign T1146 = T1147;
  assign T1147 = T1148;
  assign T1148 = T1152[T1149];
  assign T1149 = T1150;
  assign T1150 = T1151;
  assign T1151 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T1152 = T1153;
  assign T1153 = io_chanxy_in[9'h13e/* 318*/:9'h13d/* 317*/];
  assign T1154 = T1155;
  assign T1155 = T1156;
  assign T1156 = T1160[T1157];
  assign T1157 = T1158;
  assign T1158 = T1159;
  assign T1159 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T1160 = T1161;
  assign T1161 = io_chanxy_in[9'h140/* 320*/:9'h13f/* 319*/];
  assign T1162 = T1163;
  assign T1163 = T1164;
  assign T1164 = T1168[T1165];
  assign T1165 = T1166;
  assign T1166 = T1167;
  assign T1167 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T1168 = T1169;
  assign T1169 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T1170 = T1171;
  assign T1171 = T1172;
  assign T1172 = T1176[T1173];
  assign T1173 = T1174;
  assign T1174 = T1175;
  assign T1175 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T1176 = T1177;
  assign T1177 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T1178 = T1179;
  assign T1179 = T1180;
  assign T1180 = T1184[T1181];
  assign T1181 = T1182;
  assign T1182 = T1183;
  assign T1183 = io_chanxy_config[8'h9b/* 155*/:8'h9b/* 155*/];
  assign T1184 = T1185;
  assign T1185 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T1186 = T1187;
  assign T1187 = T1188;
  assign T1188 = T1192[T1189];
  assign T1189 = T1190;
  assign T1190 = T1191;
  assign T1191 = io_chanxy_config[8'h9c/* 156*/:8'h9c/* 156*/];
  assign T1192 = T1193;
  assign T1193 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T1194 = T1195;
  assign T1195 = T1196;
  assign T1196 = T1200[T1197];
  assign T1197 = T1198;
  assign T1198 = T1199;
  assign T1199 = io_chanxy_config[8'h9d/* 157*/:8'h9d/* 157*/];
  assign T1200 = T1201;
  assign T1201 = io_chanxy_in[9'h14a/* 330*/:9'h149/* 329*/];
  assign T1202 = T1203;
  assign T1203 = T1204;
  assign T1204 = T1208[T1205];
  assign T1205 = T1206;
  assign T1206 = T1207;
  assign T1207 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T1208 = T1209;
  assign T1209 = io_chanxy_in[9'h14c/* 332*/:9'h14b/* 331*/];
  assign T1210 = T1211;
  assign T1211 = T1212;
  assign T1212 = T1216[T1213];
  assign T1213 = T1214;
  assign T1214 = T1215;
  assign T1215 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T1216 = T1217;
  assign T1217 = io_chanxy_in[9'h14e/* 334*/:9'h14d/* 333*/];
  assign T1218 = T1219;
  assign T1219 = T1220;
  assign T1220 = T1224[T1221];
  assign T1221 = T1222;
  assign T1222 = T1223;
  assign T1223 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T1224 = T1225;
  assign T1225 = io_chanxy_in[9'h150/* 336*/:9'h14f/* 335*/];
  assign T1226 = T1227;
  assign T1227 = T1228;
  assign T1228 = T1232[T1229];
  assign T1229 = T1230;
  assign T1230 = T1231;
  assign T1231 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T1232 = T1233;
  assign T1233 = io_chanxy_in[9'h152/* 338*/:9'h151/* 337*/];
  assign T1234 = T1235;
  assign T1235 = T1236;
  assign T1236 = T1240[T1237];
  assign T1237 = T1238;
  assign T1238 = T1239;
  assign T1239 = io_chanxy_config[8'ha2/* 162*/:8'ha2/* 162*/];
  assign T1240 = T1241;
  assign T1241 = io_chanxy_in[9'h154/* 340*/:9'h153/* 339*/];
  assign T1242 = T1243;
  assign T1243 = T1244;
  assign T1244 = T1248[T1245];
  assign T1245 = T1246;
  assign T1246 = T1247;
  assign T1247 = io_chanxy_config[8'ha3/* 163*/:8'ha3/* 163*/];
  assign T1248 = T1249;
  assign T1249 = io_chanxy_in[9'h156/* 342*/:9'h155/* 341*/];
  assign T1250 = T1251;
  assign T1251 = T1252;
  assign T1252 = T1256[T1253];
  assign T1253 = T1254;
  assign T1254 = T1255;
  assign T1255 = io_chanxy_config[8'ha4/* 164*/:8'ha4/* 164*/];
  assign T1256 = T1257;
  assign T1257 = io_chanxy_in[9'h158/* 344*/:9'h157/* 343*/];
  assign T1258 = T1259;
  assign T1259 = T1260;
  assign T1260 = T1264[T1261];
  assign T1261 = T1262;
  assign T1262 = T1263;
  assign T1263 = io_chanxy_config[8'ha8/* 168*/:8'ha5/* 165*/];
  assign T1264 = T1265;
  assign T1265 = io_chanxy_in[9'h161/* 353*/:9'h159/* 345*/];
  assign T1266 = T1267;
  assign T1267 = T1268;
  assign T1268 = T1272[T1269];
  assign T1269 = T1270;
  assign T1270 = T1271;
  assign T1271 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T1272 = T1273;
  assign T1273 = io_chanxy_in[9'h163/* 355*/:9'h162/* 354*/];
  assign T1274 = T1275;
  assign T1275 = T1276;
  assign T1276 = T1280[T1277];
  assign T1277 = T1278;
  assign T1278 = T1279;
  assign T1279 = io_chanxy_config[8'had/* 173*/:8'haa/* 170*/];
  assign T1280 = T1281;
  assign T1281 = io_chanxy_in[9'h16c/* 364*/:9'h164/* 356*/];
  assign T1282 = T1283;
  assign T1283 = T1284;
  assign T1284 = T1288[T1285];
  assign T1285 = T1286;
  assign T1286 = T1287;
  assign T1287 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T1288 = T1289;
  assign T1289 = io_chanxy_in[9'h16e/* 366*/:9'h16d/* 365*/];
  assign T1290 = T1291;
  assign T1291 = T1292;
  assign T1292 = T1296[T1293];
  assign T1293 = T1294;
  assign T1294 = T1295;
  assign T1295 = io_chanxy_config[8'hb2/* 178*/:8'haf/* 175*/];
  assign T1296 = T1297;
  assign T1297 = io_chanxy_in[9'h177/* 375*/:9'h16f/* 367*/];
  assign T1298 = T1299;
  assign T1299 = T1300;
  assign T1300 = T1304[T1301];
  assign T1301 = T1302;
  assign T1302 = T1303;
  assign T1303 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1304 = T1305;
  assign T1305 = io_chanxy_in[9'h179/* 377*/:9'h178/* 376*/];
  assign T1306 = T1307;
  assign T1307 = T1308;
  assign T1308 = T1312[T1309];
  assign T1309 = T1310;
  assign T1310 = T1311;
  assign T1311 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T1312 = T1313;
  assign T1313 = io_chanxy_in[9'h182/* 386*/:9'h17a/* 378*/];
  assign T1314 = T1315;
  assign T1315 = T1316;
  assign T1316 = T1320[T1317];
  assign T1317 = T1318;
  assign T1318 = T1319;
  assign T1319 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1320 = T1321;
  assign T1321 = io_chanxy_in[9'h184/* 388*/:9'h183/* 387*/];
  assign T1322 = T1323;
  assign T1323 = T1324;
  assign T1324 = T1328[T1325];
  assign T1325 = T1326;
  assign T1326 = T1327;
  assign T1327 = io_chanxy_config[8'hbc/* 188*/:8'hb9/* 185*/];
  assign T1328 = T1329;
  assign T1329 = io_chanxy_in[9'h18d/* 397*/:9'h185/* 389*/];
  assign T1330 = T1331;
  assign T1331 = T1332;
  assign T1332 = T1336[T1333];
  assign T1333 = T1334;
  assign T1334 = T1335;
  assign T1335 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1336 = T1337;
  assign T1337 = io_chanxy_in[9'h18f/* 399*/:9'h18e/* 398*/];
  assign T1338 = T1339;
  assign T1339 = T1340;
  assign T1340 = T1344[T1341];
  assign T1341 = T1342;
  assign T1342 = T1343;
  assign T1343 = io_chanxy_config[8'hc1/* 193*/:8'hbe/* 190*/];
  assign T1344 = T1345;
  assign T1345 = io_chanxy_in[9'h198/* 408*/:9'h190/* 400*/];
  assign T1346 = T1347;
  assign T1347 = T1348;
  assign T1348 = T1352[T1349];
  assign T1349 = T1350;
  assign T1350 = T1351;
  assign T1351 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1352 = T1353;
  assign T1353 = io_chanxy_in[9'h19a/* 410*/:9'h199/* 409*/];
  assign T1354 = T1355;
  assign T1355 = T1356;
  assign T1356 = T1360[T1357];
  assign T1357 = T1358;
  assign T1358 = T1359;
  assign T1359 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T1360 = T1361;
  assign T1361 = io_chanxy_in[9'h1a3/* 419*/:9'h19b/* 411*/];
  assign T1362 = T1363;
  assign T1363 = T1364;
  assign T1364 = T1368[T1365];
  assign T1365 = T1366;
  assign T1366 = T1367;
  assign T1367 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1368 = T1369;
  assign T1369 = io_chanxy_in[9'h1a5/* 421*/:9'h1a4/* 420*/];
  assign T1370 = T1371;
  assign T1371 = T1372;
  assign T1372 = T1376[T1373];
  assign T1373 = T1374;
  assign T1374 = T1375;
  assign T1375 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T1376 = T1377;
  assign T1377 = io_chanxy_in[9'h1ae/* 430*/:9'h1a6/* 422*/];
  assign T1378 = T1379;
  assign T1379 = T1380;
  assign T1380 = T1384[T1381];
  assign T1381 = T1382;
  assign T1382 = T1383;
  assign T1383 = io_chanxy_config[8'hcc/* 204*/:8'hcc/* 204*/];
  assign T1384 = T1385;
  assign T1385 = io_chanxy_in[9'h1b0/* 432*/:9'h1af/* 431*/];
  assign T1386 = T1387;
  assign T1387 = T1388;
  assign T1388 = T1392[T1389];
  assign T1389 = T1390;
  assign T1390 = T1391;
  assign T1391 = io_chanxy_config[8'hd0/* 208*/:8'hcd/* 205*/];
  assign T1392 = T1393;
  assign T1393 = io_chanxy_in[9'h1b9/* 441*/:9'h1b1/* 433*/];
  assign T1394 = T1395;
  assign T1395 = T1396;
  assign T1396 = T1400[T1397];
  assign T1397 = T1398;
  assign T1398 = T1399;
  assign T1399 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T1400 = T1401;
  assign T1401 = io_chanxy_in[9'h1bb/* 443*/:9'h1ba/* 442*/];
  assign T1402 = T1403;
  assign T1403 = T1404;
  assign T1404 = T1408[T1405];
  assign T1405 = T1406;
  assign T1406 = T1407;
  assign T1407 = io_chanxy_config[8'hd5/* 213*/:8'hd2/* 210*/];
  assign T1408 = T1409;
  assign T1409 = io_chanxy_in[9'h1c4/* 452*/:9'h1bc/* 444*/];
  assign T1410 = T1411;
  assign T1411 = T1412;
  assign T1412 = T1416[T1413];
  assign T1413 = T1414;
  assign T1414 = T1415;
  assign T1415 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T1416 = T1417;
  assign T1417 = io_chanxy_in[9'h1c6/* 454*/:9'h1c5/* 453*/];
  assign T1418 = T1419;
  assign T1419 = T1420;
  assign T1420 = T1424[T1421];
  assign T1421 = T1422;
  assign T1422 = T1423;
  assign T1423 = io_chanxy_config[8'hda/* 218*/:8'hd7/* 215*/];
  assign T1424 = T1425;
  assign T1425 = io_chanxy_in[9'h1cf/* 463*/:9'h1c7/* 455*/];
  assign T1426 = T1427;
  assign T1427 = T1428;
  assign T1428 = T1432[T1429];
  assign T1429 = T1430;
  assign T1430 = T1431;
  assign T1431 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T1432 = T1433;
  assign T1433 = io_chanxy_in[9'h1d1/* 465*/:9'h1d0/* 464*/];
  assign T1434 = T1435;
  assign T1435 = T1436;
  assign T1436 = T1440[T1437];
  assign T1437 = T1438;
  assign T1438 = T1439;
  assign T1439 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1440 = T1441;
  assign T1441 = io_chanxy_in[9'h1da/* 474*/:9'h1d2/* 466*/];
  assign T1442 = T1443;
  assign T1443 = T1444;
  assign T1444 = T1448[T1445];
  assign T1445 = T1446;
  assign T1446 = T1447;
  assign T1447 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T1448 = T1449;
  assign T1449 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T1450 = T1451;
  assign T1451 = T1452;
  assign T1452 = T1456[T1453];
  assign T1453 = T1454;
  assign T1454 = T1455;
  assign T1455 = io_chanxy_config[8'he4/* 228*/:8'he1/* 225*/];
  assign T1456 = T1457;
  assign T1457 = io_chanxy_in[9'h1e5/* 485*/:9'h1dd/* 477*/];
  assign T1458 = T1459;
  assign T1459 = T1460;
  assign T1460 = T1464[T1461];
  assign T1461 = T1462;
  assign T1462 = T1463;
  assign T1463 = io_chanxy_config[8'he5/* 229*/:8'he5/* 229*/];
  assign T1464 = T1465;
  assign T1465 = io_chanxy_in[9'h1e7/* 487*/:9'h1e6/* 486*/];
  assign T1466 = T1467;
  assign T1467 = T1468;
  assign T1468 = T1472[T1469];
  assign T1469 = T1470;
  assign T1470 = T1471;
  assign T1471 = io_chanxy_config[8'he9/* 233*/:8'he6/* 230*/];
  assign T1472 = T1473;
  assign T1473 = io_chanxy_in[9'h1f0/* 496*/:9'h1e8/* 488*/];
  assign T1474 = T1475;
  assign T1475 = T1476;
  assign T1476 = T1480[T1477];
  assign T1477 = T1478;
  assign T1478 = T1479;
  assign T1479 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T1480 = T1481;
  assign T1481 = io_chanxy_in[9'h1f2/* 498*/:9'h1f1/* 497*/];
  assign T1482 = T1483;
  assign T1483 = T1484;
  assign T1484 = T1488[T1485];
  assign T1485 = T1486;
  assign T1486 = T1487;
  assign T1487 = io_chanxy_config[8'hee/* 238*/:8'heb/* 235*/];
  assign T1488 = T1489;
  assign T1489 = io_chanxy_in[9'h1fb/* 507*/:9'h1f3/* 499*/];
  assign T1490 = T1491;
  assign T1491 = T1492;
  assign T1492 = T1496[T1493];
  assign T1493 = T1494;
  assign T1494 = T1495;
  assign T1495 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T1496 = T1497;
  assign T1497 = io_chanxy_in[9'h1fd/* 509*/:9'h1fc/* 508*/];
  assign io_ipin_out = T1498;
  assign T1498 = T1499;
  assign T1499 = {T1718, T1500};
  assign T1500 = T1501;
  assign T1501 = {T1710, T1502};
  assign T1502 = T1503;
  assign T1503 = {T1702, T1504};
  assign T1504 = T1505;
  assign T1505 = {T1694, T1506};
  assign T1506 = T1507;
  assign T1507 = {T1686, T1508};
  assign T1508 = T1509;
  assign T1509 = {T1678, T1510};
  assign T1510 = T1511;
  assign T1511 = {T1670, T1512};
  assign T1512 = T1513;
  assign T1513 = {T1662, T1514};
  assign T1514 = T1515;
  assign T1515 = {T1654, T1516};
  assign T1516 = T1517;
  assign T1517 = {T1646, T1518};
  assign T1518 = T1519;
  assign T1519 = {T1638, T1520};
  assign T1520 = T1521;
  assign T1521 = {T1630, T1522};
  assign T1522 = T1523;
  assign T1523 = {T1622, T1524};
  assign T1524 = T1525;
  assign T1525 = {T1614, T1526};
  assign T1526 = T1527;
  assign T1527 = {T1606, T1528};
  assign T1528 = T1529;
  assign T1529 = {T1598, T1530};
  assign T1530 = T1531;
  assign T1531 = {T1590, T1532};
  assign T1532 = T1533;
  assign T1533 = {T1582, T1534};
  assign T1534 = T1535;
  assign T1535 = {T1574, T1536};
  assign T1536 = T1537;
  assign T1537 = {T1566, T1538};
  assign T1538 = T1539;
  assign T1539 = {T1558, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1550, T1542};
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_19(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [24:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [509:0] io_chanxy_in,
    output[149:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[239:0] T0;
  wire[799:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[149:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h31b/* 795*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_25 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_8 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_9(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[10:0] T214;
  wire[10:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[10:0] T222;
  wire[10:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[10:0] T230;
  wire[10:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[10:0] T238;
  wire[10:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[10:0] T246;
  wire[10:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] T253;
  wire[10:0] T254;
  wire[10:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[10:0] T262;
  wire[10:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[9:0] T286;
  wire[9:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[9:0] T294;
  wire[9:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[9:0] T302;
  wire[9:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[9:0] T310;
  wire[9:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[9:0] T318;
  wire[9:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[9:0] T326;
  wire[9:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[3:0] T331;
  wire[3:0] T332;
  wire[3:0] T333;
  wire[10:0] T334;
  wire[10:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[10:0] T342;
  wire[10:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[10:0] T350;
  wire[10:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[10:0] T358;
  wire[10:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[10:0] T366;
  wire[10:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[3:0] T373;
  wire[10:0] T374;
  wire[10:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[10:0] T382;
  wire[10:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[10:0] T390;
  wire[10:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[10:0] T398;
  wire[10:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[9:0] T406;
  wire[9:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[9:0] T414;
  wire[9:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[9:0] T422;
  wire[9:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[9:0] T430;
  wire[9:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[9:0] T438;
  wire[9:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[9:0] T446;
  wire[9:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[1:0] T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[1:0] T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire[2:0] T470;
  wire[2:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[1:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[2:0] T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[3:0] T483;
  wire[3:0] T484;
  wire[3:0] T485;
  wire[10:0] T486;
  wire[10:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire[1:0] T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire[2:0] T502;
  wire[2:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[1:0] T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire[2:0] T510;
  wire[2:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire[1:0] T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire[3:0] T523;
  wire[3:0] T524;
  wire[3:0] T525;
  wire[10:0] T526;
  wire[10:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire[1:0] T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire[2:0] T534;
  wire[2:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire[1:0] T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire[2:0] T542;
  wire[2:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire[1:0] T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire[2:0] T550;
  wire[2:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire[1:0] T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire[2:0] T558;
  wire[2:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[3:0] T563;
  wire[3:0] T564;
  wire[3:0] T565;
  wire[10:0] T566;
  wire[10:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire[2:0] T574;
  wire[2:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[2:0] T582;
  wire[2:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[2:0] T590;
  wire[2:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire[2:0] T598;
  wire[2:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[3:0] T603;
  wire[3:0] T604;
  wire[3:0] T605;
  wire[10:0] T606;
  wire[10:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[1:0] T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire[2:0] T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[1:0] T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire[2:0] T630;
  wire[2:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[1:0] T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire[2:0] T638;
  wire[2:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[3:0] T643;
  wire[3:0] T644;
  wire[3:0] T645;
  wire[10:0] T646;
  wire[10:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire[1:0] T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire[2:0] T654;
  wire[2:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[1:0] T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire[2:0] T662;
  wire[2:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[1:0] T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire[2:0] T670;
  wire[2:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire[1:0] T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire[2:0] T678;
  wire[2:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[3:0] T683;
  wire[3:0] T684;
  wire[3:0] T685;
  wire[10:0] T686;
  wire[10:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire[3:0] T723;
  wire[3:0] T724;
  wire[3:0] T725;
  wire[10:0] T726;
  wire[10:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire[3:0] T763;
  wire[3:0] T764;
  wire[3:0] T765;
  wire[10:0] T766;
  wire[10:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire[3:0] T803;
  wire[3:0] T804;
  wire[3:0] T805;
  wire[10:0] T806;
  wire[10:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[1:0] T814;
  wire[1:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire[1:0] T822;
  wire[1:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire[1:0] T830;
  wire[1:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire[1:0] T838;
  wire[1:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[9:0] T846;
  wire[9:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire[1:0] T854;
  wire[1:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire[1:0] T862;
  wire[1:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire[1:0] T870;
  wire[1:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire[1:0] T878;
  wire[1:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[3:0] T883;
  wire[3:0] T884;
  wire[3:0] T885;
  wire[9:0] T886;
  wire[9:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire[1:0] T894;
  wire[1:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire[1:0] T910;
  wire[1:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[9:0] T926;
  wire[9:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire[1:0] T942;
  wire[1:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire[1:0] T950;
  wire[1:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire[1:0] T958;
  wire[1:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire[3:0] T963;
  wire[3:0] T964;
  wire[3:0] T965;
  wire[9:0] T966;
  wire[9:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire[1:0] T974;
  wire[1:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire[1:0] T982;
  wire[1:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire[1:0] T990;
  wire[1:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire[1:0] T998;
  wire[1:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire[1:0] T1022;
  wire[1:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire[1:0] T1038;
  wire[1:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire[3:0] T1045;
  wire[9:0] T1046;
  wire[9:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[7'h6c/* 108*/:7'h63/* 99*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[7'h76/* 118*/:7'h6d/* 109*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[8'h80/* 128*/:7'h77/* 119*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[8'h8a/* 138*/:8'h81/* 129*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[8'h94/* 148*/:8'h8b/* 139*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[8'h9e/* 158*/:8'h95/* 149*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[8'ha9/* 169*/:8'h9f/* 159*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[8'hb4/* 180*/:8'haa/* 170*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[8'hbf/* 191*/:8'hb5/* 181*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[8'hd5/* 213*/:8'hcb/* 203*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[8'he0/* 224*/:8'hd6/* 214*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[8'heb/* 235*/:8'he1/* 225*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[8'hf6/* 246*/:8'hec/* 236*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[9'h101/* 257*/:8'hf7/* 247*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[9'h10b/* 267*/:9'h102/* 258*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[9'h115/* 277*/:9'h10c/* 268*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[9'h11f/* 287*/:9'h116/* 278*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[9'h129/* 297*/:9'h120/* 288*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[9'h133/* 307*/:9'h12a/* 298*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[9'h13d/* 317*/:9'h134/* 308*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[9'h140/* 320*/:9'h13e/* 318*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[9'h143/* 323*/:9'h141/* 321*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[9'h146/* 326*/:9'h144/* 324*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h7f/* 127*/:7'h7e/* 126*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[9'h149/* 329*/:9'h147/* 327*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[9'h154/* 340*/:9'h14a/* 330*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[8'h85/* 133*/:8'h84/* 132*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[9'h157/* 343*/:9'h155/* 341*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[8'h87/* 135*/:8'h86/* 134*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[9'h15a/* 346*/:9'h158/* 344*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[8'h89/* 137*/:8'h88/* 136*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[9'h15d/* 349*/:9'h15b/* 347*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[9'h160/* 352*/:9'h15e/* 350*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[9'h16b/* 363*/:9'h161/* 353*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[8'h91/* 145*/:8'h90/* 144*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[9'h16e/* 366*/:9'h16c/* 364*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[8'h93/* 147*/:8'h92/* 146*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[9'h171/* 369*/:9'h16f/* 367*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[8'h95/* 149*/:8'h94/* 148*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[9'h174/* 372*/:9'h172/* 370*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[8'h97/* 151*/:8'h96/* 150*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[9'h177/* 375*/:9'h175/* 373*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[9'h182/* 386*/:9'h178/* 376*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[8'h9d/* 157*/:8'h9c/* 156*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[9'h185/* 389*/:9'h183/* 387*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[8'h9f/* 159*/:8'h9e/* 158*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[9'h188/* 392*/:9'h186/* 390*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[9'h18b/* 395*/:9'h189/* 393*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[9'h18e/* 398*/:9'h18c/* 396*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[9'h199/* 409*/:9'h18f/* 399*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[9'h19c/* 412*/:9'h19a/* 410*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[9'h19f/* 415*/:9'h19d/* 413*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[9'h1a2/* 418*/:9'h1a0/* 416*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[9'h1a5/* 421*/:9'h1a3/* 419*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[9'h1b0/* 432*/:9'h1a6/* 422*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[9'h1b3/* 435*/:9'h1b1/* 433*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[9'h1b6/* 438*/:9'h1b4/* 436*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[9'h1b9/* 441*/:9'h1b7/* 439*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[8'hbb/* 187*/:8'hba/* 186*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[9'h1bc/* 444*/:9'h1ba/* 442*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[9'h1c7/* 455*/:9'h1bd/* 445*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h1cd/* 461*/:9'h1cc/* 460*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[8'hc3/* 195*/:8'hc3/* 195*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h1cf/* 463*/:9'h1ce/* 462*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h1da/* 474*/:9'h1d0/* 464*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'hc9/* 201*/:8'hc9/* 201*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h1de/* 478*/:9'h1dd/* 477*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'hca/* 202*/:8'hca/* 202*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h1e0/* 480*/:9'h1df/* 479*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'hcb/* 203*/:8'hcb/* 203*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h1e2/* 482*/:9'h1e1/* 481*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h1ed/* 493*/:9'h1e3/* 483*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h1f3/* 499*/:9'h1f2/* 498*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'hd3/* 211*/:8'hd3/* 211*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h1f5/* 501*/:9'h1f4/* 500*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[10'h200/* 512*/:9'h1f6/* 502*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[10'h202/* 514*/:10'h201/* 513*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[10'h204/* 516*/:10'h203/* 515*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[10'h206/* 518*/:10'h205/* 517*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[10'h208/* 520*/:10'h207/* 519*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[10'h212/* 530*/:10'h209/* 521*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[10'h214/* 532*/:10'h213/* 531*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[10'h216/* 534*/:10'h215/* 533*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'he2/* 226*/:8'he2/* 226*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[10'h218/* 536*/:10'h217/* 535*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'he3/* 227*/:8'he3/* 227*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[10'h21a/* 538*/:10'h219/* 537*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[10'h224/* 548*/:10'h21b/* 539*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[10'h226/* 550*/:10'h225/* 549*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[10'h228/* 552*/:10'h227/* 551*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[10'h22a/* 554*/:10'h229/* 553*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'heb/* 235*/:8'heb/* 235*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[10'h22c/* 556*/:10'h22b/* 555*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[10'h236/* 566*/:10'h22d/* 557*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[10'h238/* 568*/:10'h237/* 567*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[10'h23a/* 570*/:10'h239/* 569*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[10'h23c/* 572*/:10'h23b/* 571*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[10'h23e/* 574*/:10'h23d/* 573*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h248/* 584*/:10'h23f/* 575*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h24a/* 586*/:10'h249/* 585*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h24c/* 588*/:10'h24b/* 587*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'hfa/* 250*/:8'hfa/* 250*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h24e/* 590*/:10'h24d/* 589*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hfb/* 251*/:8'hfb/* 251*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h250/* 592*/:10'h24f/* 591*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h25a/* 602*/:10'h251/* 593*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h25c/* 604*/:10'h25b/* 603*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h25e/* 606*/:10'h25d/* 605*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h260/* 608*/:10'h25f/* 607*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h103/* 259*/:9'h103/* 259*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h262/* 610*/:10'h261/* 609*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h263/* 611*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_20(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_9 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_10(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[10:0] T214;
  wire[10:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[10:0] T222;
  wire[10:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[10:0] T230;
  wire[10:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[10:0] T238;
  wire[10:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[10:0] T246;
  wire[10:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] T253;
  wire[10:0] T254;
  wire[10:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[10:0] T262;
  wire[10:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[9:0] T286;
  wire[9:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[9:0] T294;
  wire[9:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[9:0] T302;
  wire[9:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[9:0] T310;
  wire[9:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[9:0] T318;
  wire[9:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[9:0] T326;
  wire[9:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[3:0] T331;
  wire[3:0] T332;
  wire[3:0] T333;
  wire[10:0] T334;
  wire[10:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[10:0] T342;
  wire[10:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[10:0] T350;
  wire[10:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[10:0] T358;
  wire[10:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[10:0] T366;
  wire[10:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[3:0] T373;
  wire[10:0] T374;
  wire[10:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[10:0] T382;
  wire[10:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[10:0] T390;
  wire[10:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[10:0] T398;
  wire[10:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[9:0] T406;
  wire[9:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[9:0] T414;
  wire[9:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[9:0] T422;
  wire[9:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[9:0] T430;
  wire[9:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[9:0] T438;
  wire[9:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[9:0] T446;
  wire[9:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[3:0] T459;
  wire[3:0] T460;
  wire[3:0] T461;
  wire[10:0] T462;
  wire[10:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[1:0] T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire[2:0] T470;
  wire[2:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[1:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[2:0] T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[1:0] T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire[2:0] T486;
  wire[2:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire[3:0] T499;
  wire[3:0] T500;
  wire[3:0] T501;
  wire[10:0] T502;
  wire[10:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[1:0] T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire[2:0] T510;
  wire[2:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire[1:0] T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire[1:0] T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[2:0] T526;
  wire[2:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire[1:0] T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire[2:0] T534;
  wire[2:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire[3:0] T539;
  wire[3:0] T540;
  wire[3:0] T541;
  wire[10:0] T542;
  wire[10:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire[1:0] T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire[2:0] T550;
  wire[2:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire[1:0] T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire[2:0] T558;
  wire[2:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[1:0] T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire[2:0] T566;
  wire[2:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire[2:0] T574;
  wire[2:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[3:0] T579;
  wire[3:0] T580;
  wire[3:0] T581;
  wire[10:0] T582;
  wire[10:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[2:0] T590;
  wire[2:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire[2:0] T598;
  wire[2:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[1:0] T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire[2:0] T606;
  wire[2:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[3:0] T619;
  wire[3:0] T620;
  wire[3:0] T621;
  wire[10:0] T622;
  wire[10:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[1:0] T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire[2:0] T630;
  wire[2:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[1:0] T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire[2:0] T638;
  wire[2:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[1:0] T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire[2:0] T646;
  wire[2:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire[1:0] T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire[2:0] T654;
  wire[2:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[3:0] T659;
  wire[3:0] T660;
  wire[3:0] T661;
  wire[10:0] T662;
  wire[10:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[1:0] T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire[2:0] T670;
  wire[2:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire[1:0] T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire[2:0] T678;
  wire[2:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[1:0] T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire[2:0] T686;
  wire[2:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire[3:0] T699;
  wire[3:0] T700;
  wire[3:0] T701;
  wire[10:0] T702;
  wire[10:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire[3:0] T739;
  wire[3:0] T740;
  wire[3:0] T741;
  wire[10:0] T742;
  wire[10:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire[3:0] T779;
  wire[3:0] T780;
  wire[3:0] T781;
  wire[10:0] T782;
  wire[10:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[1:0] T814;
  wire[1:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[3:0] T819;
  wire[3:0] T820;
  wire[3:0] T821;
  wire[9:0] T822;
  wire[9:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire[1:0] T830;
  wire[1:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire[1:0] T838;
  wire[1:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire[1:0] T846;
  wire[1:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire[1:0] T854;
  wire[1:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[9:0] T862;
  wire[9:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire[1:0] T870;
  wire[1:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire[1:0] T878;
  wire[1:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire[1:0] T886;
  wire[1:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire[1:0] T894;
  wire[1:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire[3:0] T901;
  wire[9:0] T902;
  wire[9:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire[1:0] T910;
  wire[1:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire[1:0] T926;
  wire[1:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[9:0] T942;
  wire[9:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire[1:0] T950;
  wire[1:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire[1:0] T958;
  wire[1:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire[1:0] T966;
  wire[1:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire[1:0] T974;
  wire[1:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire[3:0] T979;
  wire[3:0] T980;
  wire[3:0] T981;
  wire[9:0] T982;
  wire[9:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire[1:0] T990;
  wire[1:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire[1:0] T998;
  wire[1:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire[1:0] T1006;
  wire[1:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire[1:0] T1038;
  wire[1:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire[1:0] T1046;
  wire[1:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[7'h6c/* 108*/:7'h63/* 99*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[7'h76/* 118*/:7'h6d/* 109*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[8'h80/* 128*/:7'h77/* 119*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[8'h8a/* 138*/:8'h81/* 129*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[8'h94/* 148*/:8'h8b/* 139*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[8'h9e/* 158*/:8'h95/* 149*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[8'ha9/* 169*/:8'h9f/* 159*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[8'hb4/* 180*/:8'haa/* 170*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[8'hbf/* 191*/:8'hb5/* 181*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[8'hd5/* 213*/:8'hcb/* 203*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[8'he0/* 224*/:8'hd6/* 214*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[8'heb/* 235*/:8'he1/* 225*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[8'hf6/* 246*/:8'hec/* 236*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[9'h101/* 257*/:8'hf7/* 247*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[9'h10b/* 267*/:9'h102/* 258*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[9'h115/* 277*/:9'h10c/* 268*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[9'h11f/* 287*/:9'h116/* 278*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[9'h129/* 297*/:9'h120/* 288*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[9'h133/* 307*/:9'h12a/* 298*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[9'h13d/* 317*/:9'h134/* 308*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[9'h140/* 320*/:9'h13e/* 318*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h7d/* 125*/:7'h7a/* 122*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[9'h14b/* 331*/:9'h141/* 321*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h7f/* 127*/:7'h7e/* 126*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[9'h14e/* 334*/:9'h14c/* 332*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[8'h81/* 129*/:8'h80/* 128*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[9'h151/* 337*/:9'h14f/* 335*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[9'h154/* 340*/:9'h152/* 338*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[8'h85/* 133*/:8'h84/* 132*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[9'h157/* 343*/:9'h155/* 341*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[8'h89/* 137*/:8'h86/* 134*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[9'h162/* 354*/:9'h158/* 344*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[9'h165/* 357*/:9'h163/* 355*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[9'h168/* 360*/:9'h166/* 358*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[9'h16b/* 363*/:9'h169/* 361*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[8'h91/* 145*/:8'h90/* 144*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[9'h16e/* 366*/:9'h16c/* 364*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[8'h95/* 149*/:8'h92/* 146*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[9'h179/* 377*/:9'h16f/* 367*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[8'h97/* 151*/:8'h96/* 150*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[9'h17c/* 380*/:9'h17a/* 378*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[8'h99/* 153*/:8'h98/* 152*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[9'h17f/* 383*/:9'h17d/* 381*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[9'h182/* 386*/:9'h180/* 384*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[8'h9d/* 157*/:8'h9c/* 156*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[9'h185/* 389*/:9'h183/* 387*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[8'ha1/* 161*/:8'h9e/* 158*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[9'h190/* 400*/:9'h186/* 390*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[9'h193/* 403*/:9'h191/* 401*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[9'h196/* 406*/:9'h194/* 404*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[9'h199/* 409*/:9'h197/* 407*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[9'h19c/* 412*/:9'h19a/* 410*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[8'had/* 173*/:8'haa/* 170*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[9'h1a7/* 423*/:9'h19d/* 413*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[9'h1aa/* 426*/:9'h1a8/* 424*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[9'h1ad/* 429*/:9'h1ab/* 427*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[9'h1b0/* 432*/:9'h1ae/* 430*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[9'h1b3/* 435*/:9'h1b1/* 433*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[8'hb9/* 185*/:8'hb6/* 182*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[9'h1be/* 446*/:9'h1b4/* 436*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[8'hbb/* 187*/:8'hba/* 186*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[9'h1c1/* 449*/:9'h1bf/* 447*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[8'hbd/* 189*/:8'hbc/* 188*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[9'h1c4/* 452*/:9'h1c2/* 450*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[9'h1c7/* 455*/:9'h1c5/* 453*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[8'hc4/* 196*/:8'hc1/* 193*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h1d4/* 468*/:9'h1ca/* 458*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[8'hc5/* 197*/:8'hc5/* 197*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h1d6/* 470*/:9'h1d5/* 469*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[8'hc6/* 198*/:8'hc6/* 198*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h1d8/* 472*/:9'h1d7/* 471*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h1da/* 474*/:9'h1d9/* 473*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'hcc/* 204*/:8'hc9/* 201*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h1e7/* 487*/:9'h1dd/* 477*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'hcd/* 205*/:8'hcd/* 205*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h1e9/* 489*/:9'h1e8/* 488*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'hce/* 206*/:8'hce/* 206*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h1eb/* 491*/:9'h1ea/* 490*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'hcf/* 207*/:8'hcf/* 207*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h1ed/* 493*/:9'h1ec/* 492*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'hd4/* 212*/:8'hd1/* 209*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h1fa/* 506*/:9'h1f0/* 496*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'hd5/* 213*/:8'hd5/* 213*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h1fc/* 508*/:9'h1fb/* 507*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h1fe/* 510*/:9'h1fd/* 509*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[10'h200/* 512*/:9'h1ff/* 511*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[10'h202/* 514*/:10'h201/* 513*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'hdc/* 220*/:8'hd9/* 217*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[10'h20c/* 524*/:10'h203/* 515*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'hdd/* 221*/:8'hdd/* 221*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[10'h20e/* 526*/:10'h20d/* 525*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'hde/* 222*/:8'hde/* 222*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[10'h210/* 528*/:10'h20f/* 527*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[10'h212/* 530*/:10'h211/* 529*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[10'h214/* 532*/:10'h213/* 531*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'he4/* 228*/:8'he1/* 225*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[10'h21e/* 542*/:10'h215/* 533*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'he5/* 229*/:8'he5/* 229*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[10'h220/* 544*/:10'h21f/* 543*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'he6/* 230*/:8'he6/* 230*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[10'h222/* 546*/:10'h221/* 545*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'he7/* 231*/:8'he7/* 231*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[10'h224/* 548*/:10'h223/* 547*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[10'h226/* 550*/:10'h225/* 549*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hec/* 236*/:8'he9/* 233*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[10'h230/* 560*/:10'h227/* 551*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hed/* 237*/:8'hed/* 237*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[10'h232/* 562*/:10'h231/* 561*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hee/* 238*/:8'hee/* 238*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[10'h234/* 564*/:10'h233/* 563*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[10'h236/* 566*/:10'h235/* 565*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[10'h238/* 568*/:10'h237/* 567*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hf4/* 244*/:8'hf1/* 241*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[10'h242/* 578*/:10'h239/* 569*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hf5/* 245*/:8'hf5/* 245*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[10'h244/* 580*/:10'h243/* 579*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hf6/* 246*/:8'hf6/* 246*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[10'h246/* 582*/:10'h245/* 581*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h248/* 584*/:10'h247/* 583*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h24a/* 586*/:10'h249/* 585*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'hfc/* 252*/:8'hf9/* 249*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h254/* 596*/:10'h24b/* 587*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'hfd/* 253*/:8'hfd/* 253*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h256/* 598*/:10'h255/* 597*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hfe/* 254*/:8'hfe/* 254*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h258/* 600*/:10'h257/* 599*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hff/* 255*/:8'hff/* 255*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h25a/* 602*/:10'h259/* 601*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h25c/* 604*/:10'h25b/* 603*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[9'h104/* 260*/:9'h101/* 257*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h266/* 614*/:10'h25d/* 605*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[9'h105/* 261*/:9'h105/* 261*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h268/* 616*/:10'h267/* 615*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h106/* 262*/:9'h106/* 262*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h26a/* 618*/:10'h269/* 617*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h26b/* 619*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_21(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_10 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_11(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[10:0] T214;
  wire[10:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[10:0] T222;
  wire[10:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[10:0] T230;
  wire[10:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[10:0] T238;
  wire[10:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[10:0] T246;
  wire[10:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] T253;
  wire[10:0] T254;
  wire[10:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[10:0] T262;
  wire[10:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[9:0] T286;
  wire[9:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[9:0] T294;
  wire[9:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[9:0] T302;
  wire[9:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[9:0] T310;
  wire[9:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[9:0] T318;
  wire[9:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[9:0] T326;
  wire[9:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[3:0] T331;
  wire[3:0] T332;
  wire[3:0] T333;
  wire[10:0] T334;
  wire[10:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[10:0] T342;
  wire[10:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[10:0] T350;
  wire[10:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[10:0] T358;
  wire[10:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[10:0] T366;
  wire[10:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[3:0] T373;
  wire[10:0] T374;
  wire[10:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[10:0] T382;
  wire[10:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[10:0] T390;
  wire[10:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[10:0] T398;
  wire[10:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[9:0] T406;
  wire[9:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[9:0] T414;
  wire[9:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[9:0] T422;
  wire[9:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[9:0] T430;
  wire[9:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[9:0] T438;
  wire[9:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[9:0] T446;
  wire[9:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[1:0] T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[3:0] T467;
  wire[3:0] T468;
  wire[3:0] T469;
  wire[10:0] T470;
  wire[10:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[1:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[2:0] T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[1:0] T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire[2:0] T486;
  wire[2:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire[1:0] T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire[2:0] T502;
  wire[2:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[3:0] T507;
  wire[3:0] T508;
  wire[3:0] T509;
  wire[10:0] T510;
  wire[10:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire[1:0] T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire[2:0] T518;
  wire[2:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire[1:0] T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[2:0] T526;
  wire[2:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire[1:0] T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire[2:0] T534;
  wire[2:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire[1:0] T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire[2:0] T542;
  wire[2:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire[3:0] T547;
  wire[3:0] T548;
  wire[3:0] T549;
  wire[10:0] T550;
  wire[10:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire[1:0] T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire[2:0] T558;
  wire[2:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[1:0] T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire[2:0] T566;
  wire[2:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire[2:0] T574;
  wire[2:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[2:0] T582;
  wire[2:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[3:0] T587;
  wire[3:0] T588;
  wire[3:0] T589;
  wire[10:0] T590;
  wire[10:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire[2:0] T598;
  wire[2:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[1:0] T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire[2:0] T606;
  wire[2:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[1:0] T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire[2:0] T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[3:0] T627;
  wire[3:0] T628;
  wire[3:0] T629;
  wire[10:0] T630;
  wire[10:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[1:0] T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire[2:0] T638;
  wire[2:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[1:0] T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire[2:0] T646;
  wire[2:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire[1:0] T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire[2:0] T654;
  wire[2:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[1:0] T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire[2:0] T662;
  wire[2:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[3:0] T667;
  wire[3:0] T668;
  wire[3:0] T669;
  wire[10:0] T670;
  wire[10:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire[1:0] T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire[2:0] T678;
  wire[2:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[1:0] T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire[2:0] T686;
  wire[2:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire[3:0] T707;
  wire[3:0] T708;
  wire[3:0] T709;
  wire[10:0] T710;
  wire[10:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire T716;
  wire T717;
  wire[1:0] T718;
  wire[1:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire[3:0] T747;
  wire[3:0] T748;
  wire[3:0] T749;
  wire[10:0] T750;
  wire[10:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire[3:0] T787;
  wire[3:0] T788;
  wire[3:0] T789;
  wire[10:0] T790;
  wire[10:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[1:0] T814;
  wire[1:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire[1:0] T822;
  wire[1:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[9:0] T830;
  wire[9:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire T836;
  wire T837;
  wire[1:0] T838;
  wire[1:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire[1:0] T846;
  wire[1:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire[1:0] T854;
  wire[1:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire[1:0] T862;
  wire[1:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[3:0] T867;
  wire[3:0] T868;
  wire[3:0] T869;
  wire[9:0] T870;
  wire[9:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire[1:0] T878;
  wire[1:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire[1:0] T886;
  wire[1:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire[1:0] T894;
  wire[1:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[9:0] T910;
  wire[9:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire[1:0] T926;
  wire[1:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire[1:0] T942;
  wire[1:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire[3:0] T947;
  wire[3:0] T948;
  wire[3:0] T949;
  wire[9:0] T950;
  wire[9:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire[1:0] T958;
  wire[1:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire[1:0] T966;
  wire[1:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire[1:0] T974;
  wire[1:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire[1:0] T982;
  wire[1:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[9:0] T990;
  wire[9:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire[1:0] T998;
  wire[1:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire[1:0] T1006;
  wire[1:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire[1:0] T1022;
  wire[1:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire[3:0] T1027;
  wire[3:0] T1028;
  wire[3:0] T1029;
  wire[9:0] T1030;
  wire[9:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire[1:0] T1038;
  wire[1:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire[1:0] T1046;
  wire[1:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[7'h6c/* 108*/:7'h63/* 99*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[7'h76/* 118*/:7'h6d/* 109*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[8'h80/* 128*/:7'h77/* 119*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[8'h8a/* 138*/:8'h81/* 129*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[8'h94/* 148*/:8'h8b/* 139*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[8'h9e/* 158*/:8'h95/* 149*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[8'ha9/* 169*/:8'h9f/* 159*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[8'hb4/* 180*/:8'haa/* 170*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[8'hbf/* 191*/:8'hb5/* 181*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[8'hd5/* 213*/:8'hcb/* 203*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[8'he0/* 224*/:8'hd6/* 214*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[8'heb/* 235*/:8'he1/* 225*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[8'hf6/* 246*/:8'hec/* 236*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[9'h101/* 257*/:8'hf7/* 247*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[9'h10b/* 267*/:9'h102/* 258*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[9'h115/* 277*/:9'h10c/* 268*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[9'h11f/* 287*/:9'h116/* 278*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[9'h129/* 297*/:9'h120/* 288*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[9'h133/* 307*/:9'h12a/* 298*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[9'h13d/* 317*/:9'h134/* 308*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[9'h140/* 320*/:9'h13e/* 318*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[9'h143/* 323*/:9'h141/* 321*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[9'h14e/* 334*/:9'h144/* 324*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[8'h81/* 129*/:8'h80/* 128*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[9'h151/* 337*/:9'h14f/* 335*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[9'h154/* 340*/:9'h152/* 338*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[8'h85/* 133*/:8'h84/* 132*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[9'h157/* 343*/:9'h155/* 341*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[8'h87/* 135*/:8'h86/* 134*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[9'h15a/* 346*/:9'h158/* 344*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[9'h165/* 357*/:9'h15b/* 347*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[9'h168/* 360*/:9'h166/* 358*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[9'h16b/* 363*/:9'h169/* 361*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[8'h91/* 145*/:8'h90/* 144*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[9'h16e/* 366*/:9'h16c/* 364*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[8'h93/* 147*/:8'h92/* 146*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[9'h171/* 369*/:9'h16f/* 367*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[9'h17c/* 380*/:9'h172/* 370*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[8'h99/* 153*/:8'h98/* 152*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[9'h17f/* 383*/:9'h17d/* 381*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[9'h182/* 386*/:9'h180/* 384*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[8'h9d/* 157*/:8'h9c/* 156*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[9'h185/* 389*/:9'h183/* 387*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[8'h9f/* 159*/:8'h9e/* 158*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[9'h188/* 392*/:9'h186/* 390*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[9'h193/* 403*/:9'h189/* 393*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[9'h196/* 406*/:9'h194/* 404*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[9'h199/* 409*/:9'h197/* 407*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[9'h19c/* 412*/:9'h19a/* 410*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[9'h19f/* 415*/:9'h19d/* 413*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[9'h1aa/* 426*/:9'h1a0/* 416*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[9'h1ad/* 429*/:9'h1ab/* 427*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[9'h1b0/* 432*/:9'h1ae/* 430*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[9'h1b3/* 435*/:9'h1b1/* 433*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[9'h1b6/* 438*/:9'h1b4/* 436*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[8'hbb/* 187*/:8'hb8/* 184*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[9'h1c1/* 449*/:9'h1b7/* 439*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[8'hbd/* 189*/:8'hbc/* 188*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[9'h1c4/* 452*/:9'h1c2/* 450*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[9'h1c7/* 455*/:9'h1c5/* 453*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[8'hc5/* 197*/:8'hc2/* 194*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h1d6/* 470*/:9'h1cc/* 460*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[8'hc6/* 198*/:8'hc6/* 198*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h1d8/* 472*/:9'h1d7/* 471*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h1da/* 474*/:9'h1d9/* 473*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'hc9/* 201*/:8'hc9/* 201*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h1de/* 478*/:9'h1dd/* 477*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'hcd/* 205*/:8'hca/* 202*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h1e9/* 489*/:9'h1df/* 479*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'hce/* 206*/:8'hce/* 206*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h1eb/* 491*/:9'h1ea/* 490*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'hcf/* 207*/:8'hcf/* 207*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h1ed/* 493*/:9'h1ec/* 492*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'hd5/* 213*/:8'hd2/* 210*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h1fc/* 508*/:9'h1f2/* 498*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h1fe/* 510*/:9'h1fd/* 509*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[10'h200/* 512*/:9'h1ff/* 511*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[10'h202/* 514*/:10'h201/* 513*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[10'h204/* 516*/:10'h203/* 515*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'hdd/* 221*/:8'hda/* 218*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[10'h20e/* 526*/:10'h205/* 517*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'hde/* 222*/:8'hde/* 222*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[10'h210/* 528*/:10'h20f/* 527*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[10'h212/* 530*/:10'h211/* 529*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[10'h214/* 532*/:10'h213/* 531*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[10'h216/* 534*/:10'h215/* 533*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'he5/* 229*/:8'he2/* 226*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[10'h220/* 544*/:10'h217/* 535*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'he6/* 230*/:8'he6/* 230*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[10'h222/* 546*/:10'h221/* 545*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'he7/* 231*/:8'he7/* 231*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[10'h224/* 548*/:10'h223/* 547*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[10'h226/* 550*/:10'h225/* 549*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[10'h228/* 552*/:10'h227/* 551*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hed/* 237*/:8'hea/* 234*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[10'h232/* 562*/:10'h229/* 553*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hee/* 238*/:8'hee/* 238*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[10'h234/* 564*/:10'h233/* 563*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[10'h236/* 566*/:10'h235/* 565*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[10'h238/* 568*/:10'h237/* 567*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[10'h23a/* 570*/:10'h239/* 569*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hf5/* 245*/:8'hf2/* 242*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[10'h244/* 580*/:10'h23b/* 571*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hf6/* 246*/:8'hf6/* 246*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[10'h246/* 582*/:10'h245/* 581*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h248/* 584*/:10'h247/* 583*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h24a/* 586*/:10'h249/* 585*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h24c/* 588*/:10'h24b/* 587*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'hfd/* 253*/:8'hfa/* 250*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h256/* 598*/:10'h24d/* 589*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hfe/* 254*/:8'hfe/* 254*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h258/* 600*/:10'h257/* 599*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hff/* 255*/:8'hff/* 255*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h25a/* 602*/:10'h259/* 601*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h25c/* 604*/:10'h25b/* 603*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h25e/* 606*/:10'h25d/* 605*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[9'h105/* 261*/:9'h102/* 258*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h268/* 616*/:10'h25f/* 607*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h106/* 262*/:9'h106/* 262*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h26a/* 618*/:10'h269/* 617*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h26b/* 619*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_22(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_11 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_12(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [620:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[10:0] T214;
  wire[10:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[10:0] T222;
  wire[10:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[10:0] T230;
  wire[10:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[10:0] T238;
  wire[10:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[10:0] T246;
  wire[10:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] T253;
  wire[10:0] T254;
  wire[10:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[10:0] T262;
  wire[10:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[10:0] T270;
  wire[10:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[10:0] T278;
  wire[10:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[9:0] T286;
  wire[9:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[9:0] T294;
  wire[9:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[9:0] T302;
  wire[9:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[9:0] T310;
  wire[9:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[9:0] T318;
  wire[9:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[9:0] T326;
  wire[9:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[3:0] T331;
  wire[3:0] T332;
  wire[3:0] T333;
  wire[10:0] T334;
  wire[10:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[10:0] T342;
  wire[10:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[10:0] T350;
  wire[10:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[10:0] T358;
  wire[10:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[10:0] T366;
  wire[10:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[3:0] T373;
  wire[10:0] T374;
  wire[10:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[10:0] T382;
  wire[10:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[10:0] T390;
  wire[10:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[10:0] T398;
  wire[10:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[9:0] T406;
  wire[9:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[9:0] T414;
  wire[9:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[9:0] T422;
  wire[9:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[9:0] T430;
  wire[9:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[9:0] T438;
  wire[9:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[9:0] T446;
  wire[9:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[1:0] T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[1:0] T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire[2:0] T470;
  wire[2:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[3:0] T475;
  wire[3:0] T476;
  wire[3:0] T477;
  wire[10:0] T478;
  wire[10:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[1:0] T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire[2:0] T486;
  wire[2:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire[1:0] T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire[2:0] T502;
  wire[2:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire[1:0] T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire[2:0] T510;
  wire[2:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire[3:0] T515;
  wire[3:0] T516;
  wire[3:0] T517;
  wire[10:0] T518;
  wire[10:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire[1:0] T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[2:0] T526;
  wire[2:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire[1:0] T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire[2:0] T534;
  wire[2:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire[1:0] T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire[2:0] T542;
  wire[2:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire[1:0] T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire[2:0] T550;
  wire[2:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire[3:0] T555;
  wire[3:0] T556;
  wire[3:0] T557;
  wire[10:0] T558;
  wire[10:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire[1:0] T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire[2:0] T566;
  wire[2:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire[2:0] T574;
  wire[2:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[2:0] T582;
  wire[2:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[2:0] T590;
  wire[2:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[3:0] T595;
  wire[3:0] T596;
  wire[3:0] T597;
  wire[10:0] T598;
  wire[10:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[1:0] T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire[2:0] T606;
  wire[2:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire[1:0] T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire[2:0] T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire[1:0] T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire[2:0] T630;
  wire[2:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire[3:0] T635;
  wire[3:0] T636;
  wire[3:0] T637;
  wire[10:0] T638;
  wire[10:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire[1:0] T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire[2:0] T646;
  wire[2:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire[1:0] T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire[2:0] T654;
  wire[2:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire[1:0] T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire[2:0] T662;
  wire[2:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire[1:0] T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire[2:0] T670;
  wire[2:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire[3:0] T675;
  wire[3:0] T676;
  wire[3:0] T677;
  wire[10:0] T678;
  wire[10:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire[1:0] T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire[2:0] T686;
  wire[2:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire T692;
  wire T693;
  wire[1:0] T694;
  wire[1:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire T700;
  wire T701;
  wire[1:0] T702;
  wire[1:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire[1:0] T710;
  wire[1:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire[3:0] T715;
  wire[3:0] T716;
  wire[3:0] T717;
  wire[10:0] T718;
  wire[10:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire T724;
  wire T725;
  wire[1:0] T726;
  wire[1:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire[1:0] T734;
  wire[1:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire[3:0] T755;
  wire[3:0] T756;
  wire[3:0] T757;
  wire[10:0] T758;
  wire[10:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire[3:0] T795;
  wire[3:0] T796;
  wire[3:0] T797;
  wire[10:0] T798;
  wire[10:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire[1:0] T814;
  wire[1:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire T820;
  wire T821;
  wire[1:0] T822;
  wire[1:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire T828;
  wire T829;
  wire[1:0] T830;
  wire[1:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[3:0] T835;
  wire[3:0] T836;
  wire[3:0] T837;
  wire[9:0] T838;
  wire[9:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire T844;
  wire T845;
  wire[1:0] T846;
  wire[1:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire[1:0] T854;
  wire[1:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire T860;
  wire T861;
  wire[1:0] T862;
  wire[1:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire[1:0] T870;
  wire[1:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[9:0] T878;
  wire[9:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire[1:0] T886;
  wire[1:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire[1:0] T894;
  wire[1:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire[1:0] T902;
  wire[1:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire[1:0] T910;
  wire[1:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire[3:0] T915;
  wire[3:0] T916;
  wire[3:0] T917;
  wire[9:0] T918;
  wire[9:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire T924;
  wire T925;
  wire[1:0] T926;
  wire[1:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire[1:0] T942;
  wire[1:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire[1:0] T950;
  wire[1:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[9:0] T958;
  wire[9:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire[1:0] T966;
  wire[1:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire T972;
  wire T973;
  wire[1:0] T974;
  wire[1:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire[1:0] T982;
  wire[1:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire T988;
  wire T989;
  wire[1:0] T990;
  wire[1:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire[3:0] T995;
  wire[3:0] T996;
  wire[3:0] T997;
  wire[9:0] T998;
  wire[9:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire T1004;
  wire T1005;
  wire[1:0] T1006;
  wire[1:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire[1:0] T1022;
  wire[1:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire[1:0] T1046;
  wire[1:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[7'h6c/* 108*/:7'h63/* 99*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[7'h76/* 118*/:7'h6d/* 109*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[8'h80/* 128*/:7'h77/* 119*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[8'h8a/* 138*/:8'h81/* 129*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[8'h94/* 148*/:8'h8b/* 139*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[8'h9e/* 158*/:8'h95/* 149*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[8'ha9/* 169*/:8'h9f/* 159*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[8'hb4/* 180*/:8'haa/* 170*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[8'hbf/* 191*/:8'hb5/* 181*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[8'hd5/* 213*/:8'hcb/* 203*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[8'he0/* 224*/:8'hd6/* 214*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[8'heb/* 235*/:8'he1/* 225*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[8'hf6/* 246*/:8'hec/* 236*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[9'h101/* 257*/:8'hf7/* 247*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[9'h10b/* 267*/:9'h102/* 258*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[9'h115/* 277*/:9'h10c/* 268*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[9'h11f/* 287*/:9'h116/* 278*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[9'h129/* 297*/:9'h120/* 288*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[9'h133/* 307*/:9'h12a/* 298*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[9'h13d/* 317*/:9'h134/* 308*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[9'h140/* 320*/:9'h13e/* 318*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[9'h143/* 323*/:9'h141/* 321*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[9'h146/* 326*/:9'h144/* 324*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[8'h81/* 129*/:7'h7e/* 126*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[9'h151/* 337*/:9'h147/* 327*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[9'h154/* 340*/:9'h152/* 338*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[8'h85/* 133*/:8'h84/* 132*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[9'h157/* 343*/:9'h155/* 341*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[8'h87/* 135*/:8'h86/* 134*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[9'h15a/* 346*/:9'h158/* 344*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[8'h89/* 137*/:8'h88/* 136*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[9'h15d/* 349*/:9'h15b/* 347*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[9'h168/* 360*/:9'h15e/* 350*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[9'h16b/* 363*/:9'h169/* 361*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[8'h91/* 145*/:8'h90/* 144*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[9'h16e/* 366*/:9'h16c/* 364*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[8'h93/* 147*/:8'h92/* 146*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[9'h171/* 369*/:9'h16f/* 367*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[8'h95/* 149*/:8'h94/* 148*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[9'h174/* 372*/:9'h172/* 370*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[9'h17f/* 383*/:9'h175/* 373*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[8'h9b/* 155*/:8'h9a/* 154*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[9'h182/* 386*/:9'h180/* 384*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[8'h9d/* 157*/:8'h9c/* 156*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[9'h185/* 389*/:9'h183/* 387*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[8'h9f/* 159*/:8'h9e/* 158*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[9'h188/* 392*/:9'h186/* 390*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[9'h18b/* 395*/:9'h189/* 393*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[8'ha5/* 165*/:8'ha2/* 162*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[9'h196/* 406*/:9'h18c/* 396*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[9'h199/* 409*/:9'h197/* 407*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[9'h19c/* 412*/:9'h19a/* 410*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[9'h19f/* 415*/:9'h19d/* 413*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[9'h1a2/* 418*/:9'h1a0/* 416*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[8'hb1/* 177*/:8'hae/* 174*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[9'h1ad/* 429*/:9'h1a3/* 419*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[9'h1b0/* 432*/:9'h1ae/* 430*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[9'h1b3/* 435*/:9'h1b1/* 433*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[9'h1b6/* 438*/:9'h1b4/* 436*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[9'h1b9/* 441*/:9'h1b7/* 439*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[8'hbd/* 189*/:8'hba/* 186*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[9'h1c4/* 452*/:9'h1ba/* 442*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[9'h1c7/* 455*/:9'h1c5/* 453*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h1cd/* 461*/:9'h1cc/* 460*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h1da/* 474*/:9'h1d9/* 473*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h1dc/* 476*/:9'h1db/* 475*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'hc9/* 201*/:8'hc9/* 201*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h1de/* 478*/:9'h1dd/* 477*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'hca/* 202*/:8'hca/* 202*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h1e0/* 480*/:9'h1df/* 479*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'hce/* 206*/:8'hcb/* 203*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h1eb/* 491*/:9'h1e1/* 481*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'hcf/* 207*/:8'hcf/* 207*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h1ed/* 493*/:9'h1ec/* 492*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h1f3/* 499*/:9'h1f2/* 498*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'hd6/* 214*/:8'hd3/* 211*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h1fe/* 510*/:9'h1f4/* 500*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[10'h200/* 512*/:9'h1ff/* 511*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[10'h202/* 514*/:10'h201/* 513*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[10'h204/* 516*/:10'h203/* 515*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[10'h206/* 518*/:10'h205/* 517*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'hde/* 222*/:8'hdb/* 219*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[10'h210/* 528*/:10'h207/* 519*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[10'h212/* 530*/:10'h211/* 529*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[10'h214/* 532*/:10'h213/* 531*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[10'h216/* 534*/:10'h215/* 533*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'he2/* 226*/:8'he2/* 226*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[10'h218/* 536*/:10'h217/* 535*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'he6/* 230*/:8'he3/* 227*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[10'h222/* 546*/:10'h219/* 537*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'he7/* 231*/:8'he7/* 231*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[10'h224/* 548*/:10'h223/* 547*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[10'h226/* 550*/:10'h225/* 549*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[10'h228/* 552*/:10'h227/* 551*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[10'h22a/* 554*/:10'h229/* 553*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hee/* 238*/:8'heb/* 235*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[10'h234/* 564*/:10'h22b/* 555*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[10'h236/* 566*/:10'h235/* 565*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[10'h238/* 568*/:10'h237/* 567*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[10'h23a/* 570*/:10'h239/* 569*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[10'h23c/* 572*/:10'h23b/* 571*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hf6/* 246*/:8'hf3/* 243*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[10'h246/* 582*/:10'h23d/* 573*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h248/* 584*/:10'h247/* 583*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h24a/* 586*/:10'h249/* 585*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h24c/* 588*/:10'h24b/* 587*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'hfa/* 250*/:8'hfa/* 250*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h24e/* 590*/:10'h24d/* 589*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hfe/* 254*/:8'hfb/* 251*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h258/* 600*/:10'h24f/* 591*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hff/* 255*/:8'hff/* 255*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h25a/* 602*/:10'h259/* 601*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h25c/* 604*/:10'h25b/* 603*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h25e/* 606*/:10'h25d/* 605*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h260/* 608*/:10'h25f/* 607*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h106/* 262*/:9'h103/* 259*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h26a/* 618*/:10'h261/* 609*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h26c/* 620*/:10'h26b/* 619*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_23(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_12 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_24(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_9 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_25(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_10 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_26(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_11 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_27(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [620:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_12 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_13(
    input [275:0] io_ipin_in,
    input [91:0] io_ipin_config,
    input [572:0] io_chanxy_in,
    input [263:0] io_chanxy_config,
    output[22:0] io_ipin_out,
    output[104:0] io_chanxy_out);

  wire[104:0] T0;
  wire[104:0] T1;
  wire[103:0] T2;
  wire[103:0] T3;
  wire[102:0] T4;
  wire[102:0] T5;
  wire[101:0] T6;
  wire[101:0] T7;
  wire[100:0] T8;
  wire[100:0] T9;
  wire[99:0] T10;
  wire[99:0] T11;
  wire[98:0] T12;
  wire[98:0] T13;
  wire[97:0] T14;
  wire[97:0] T15;
  wire[96:0] T16;
  wire[96:0] T17;
  wire[95:0] T18;
  wire[95:0] T19;
  wire[94:0] T20;
  wire[94:0] T21;
  wire[93:0] T22;
  wire[93:0] T23;
  wire[92:0] T24;
  wire[92:0] T25;
  wire[91:0] T26;
  wire[91:0] T27;
  wire[90:0] T28;
  wire[90:0] T29;
  wire[89:0] T30;
  wire[89:0] T31;
  wire[88:0] T32;
  wire[88:0] T33;
  wire[87:0] T34;
  wire[87:0] T35;
  wire[86:0] T36;
  wire[86:0] T37;
  wire[85:0] T38;
  wire[85:0] T39;
  wire[84:0] T40;
  wire[84:0] T41;
  wire[83:0] T42;
  wire[83:0] T43;
  wire[82:0] T44;
  wire[82:0] T45;
  wire[81:0] T46;
  wire[81:0] T47;
  wire[80:0] T48;
  wire[80:0] T49;
  wire[79:0] T50;
  wire[79:0] T51;
  wire[78:0] T52;
  wire[78:0] T53;
  wire[77:0] T54;
  wire[77:0] T55;
  wire[76:0] T56;
  wire[76:0] T57;
  wire[75:0] T58;
  wire[75:0] T59;
  wire[74:0] T60;
  wire[74:0] T61;
  wire[73:0] T62;
  wire[73:0] T63;
  wire[72:0] T64;
  wire[72:0] T65;
  wire[71:0] T66;
  wire[71:0] T67;
  wire[70:0] T68;
  wire[70:0] T69;
  wire[69:0] T70;
  wire[69:0] T71;
  wire[68:0] T72;
  wire[68:0] T73;
  wire[67:0] T74;
  wire[67:0] T75;
  wire[66:0] T76;
  wire[66:0] T77;
  wire[65:0] T78;
  wire[65:0] T79;
  wire[64:0] T80;
  wire[64:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[62:0] T84;
  wire[62:0] T85;
  wire[61:0] T86;
  wire[61:0] T87;
  wire[60:0] T88;
  wire[60:0] T89;
  wire[59:0] T90;
  wire[59:0] T91;
  wire[58:0] T92;
  wire[58:0] T93;
  wire[57:0] T94;
  wire[57:0] T95;
  wire[56:0] T96;
  wire[56:0] T97;
  wire[55:0] T98;
  wire[55:0] T99;
  wire[54:0] T100;
  wire[54:0] T101;
  wire[53:0] T102;
  wire[53:0] T103;
  wire[52:0] T104;
  wire[52:0] T105;
  wire[51:0] T106;
  wire[51:0] T107;
  wire[50:0] T108;
  wire[50:0] T109;
  wire[49:0] T110;
  wire[49:0] T111;
  wire[48:0] T112;
  wire[48:0] T113;
  wire[47:0] T114;
  wire[47:0] T115;
  wire[46:0] T116;
  wire[46:0] T117;
  wire[45:0] T118;
  wire[45:0] T119;
  wire[44:0] T120;
  wire[44:0] T121;
  wire[43:0] T122;
  wire[43:0] T123;
  wire[42:0] T124;
  wire[42:0] T125;
  wire[41:0] T126;
  wire[41:0] T127;
  wire[40:0] T128;
  wire[40:0] T129;
  wire[39:0] T130;
  wire[39:0] T131;
  wire[38:0] T132;
  wire[38:0] T133;
  wire[37:0] T134;
  wire[37:0] T135;
  wire[36:0] T136;
  wire[36:0] T137;
  wire[35:0] T138;
  wire[35:0] T139;
  wire[34:0] T140;
  wire[34:0] T141;
  wire[33:0] T142;
  wire[33:0] T143;
  wire[32:0] T144;
  wire[32:0] T145;
  wire[31:0] T146;
  wire[31:0] T147;
  wire[30:0] T148;
  wire[30:0] T149;
  wire[29:0] T150;
  wire[29:0] T151;
  wire[28:0] T152;
  wire[28:0] T153;
  wire[27:0] T154;
  wire[27:0] T155;
  wire[26:0] T156;
  wire[26:0] T157;
  wire[25:0] T158;
  wire[25:0] T159;
  wire[24:0] T160;
  wire[24:0] T161;
  wire[23:0] T162;
  wire[23:0] T163;
  wire[22:0] T164;
  wire[22:0] T165;
  wire[21:0] T166;
  wire[21:0] T167;
  wire[20:0] T168;
  wire[20:0] T169;
  wire[19:0] T170;
  wire[19:0] T171;
  wire[18:0] T172;
  wire[18:0] T173;
  wire[17:0] T174;
  wire[17:0] T175;
  wire[16:0] T176;
  wire[16:0] T177;
  wire[15:0] T178;
  wire[15:0] T179;
  wire[14:0] T180;
  wire[14:0] T181;
  wire[13:0] T182;
  wire[13:0] T183;
  wire[12:0] T184;
  wire[12:0] T185;
  wire[11:0] T186;
  wire[11:0] T187;
  wire[10:0] T188;
  wire[10:0] T189;
  wire[9:0] T190;
  wire[9:0] T191;
  wire[8:0] T192;
  wire[8:0] T193;
  wire[7:0] T194;
  wire[7:0] T195;
  wire[6:0] T196;
  wire[6:0] T197;
  wire[5:0] T198;
  wire[5:0] T199;
  wire[4:0] T200;
  wire[4:0] T201;
  wire[3:0] T202;
  wire[3:0] T203;
  wire[2:0] T204;
  wire[2:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire T208;
  wire T209;
  wire T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[8:0] T214;
  wire[8:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire[3:0] T219;
  wire[3:0] T220;
  wire[3:0] T221;
  wire[8:0] T222;
  wire[8:0] T223;
  wire T224;
  wire T225;
  wire T226;
  wire[3:0] T227;
  wire[3:0] T228;
  wire[3:0] T229;
  wire[8:0] T230;
  wire[8:0] T231;
  wire T232;
  wire T233;
  wire T234;
  wire[3:0] T235;
  wire[3:0] T236;
  wire[3:0] T237;
  wire[8:0] T238;
  wire[8:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire[3:0] T243;
  wire[3:0] T244;
  wire[3:0] T245;
  wire[8:0] T246;
  wire[8:0] T247;
  wire T248;
  wire T249;
  wire T250;
  wire[3:0] T251;
  wire[3:0] T252;
  wire[3:0] T253;
  wire[8:0] T254;
  wire[8:0] T255;
  wire T256;
  wire T257;
  wire T258;
  wire[3:0] T259;
  wire[3:0] T260;
  wire[3:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire[3:0] T267;
  wire[3:0] T268;
  wire[3:0] T269;
  wire[8:0] T270;
  wire[8:0] T271;
  wire T272;
  wire T273;
  wire T274;
  wire[3:0] T275;
  wire[3:0] T276;
  wire[3:0] T277;
  wire[8:0] T278;
  wire[8:0] T279;
  wire T280;
  wire T281;
  wire T282;
  wire[3:0] T283;
  wire[3:0] T284;
  wire[3:0] T285;
  wire[8:0] T286;
  wire[8:0] T287;
  wire T288;
  wire T289;
  wire T290;
  wire[3:0] T291;
  wire[3:0] T292;
  wire[3:0] T293;
  wire[8:0] T294;
  wire[8:0] T295;
  wire T296;
  wire T297;
  wire T298;
  wire[3:0] T299;
  wire[3:0] T300;
  wire[3:0] T301;
  wire[8:0] T302;
  wire[8:0] T303;
  wire T304;
  wire T305;
  wire T306;
  wire[3:0] T307;
  wire[3:0] T308;
  wire[3:0] T309;
  wire[8:0] T310;
  wire[8:0] T311;
  wire T312;
  wire T313;
  wire T314;
  wire[3:0] T315;
  wire[3:0] T316;
  wire[3:0] T317;
  wire[8:0] T318;
  wire[8:0] T319;
  wire T320;
  wire T321;
  wire T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire[3:0] T325;
  wire[8:0] T326;
  wire[8:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire[3:0] T331;
  wire[3:0] T332;
  wire[3:0] T333;
  wire[8:0] T334;
  wire[8:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire[3:0] T339;
  wire[3:0] T340;
  wire[3:0] T341;
  wire[8:0] T342;
  wire[8:0] T343;
  wire T344;
  wire T345;
  wire T346;
  wire[3:0] T347;
  wire[3:0] T348;
  wire[3:0] T349;
  wire[8:0] T350;
  wire[8:0] T351;
  wire T352;
  wire T353;
  wire T354;
  wire[3:0] T355;
  wire[3:0] T356;
  wire[3:0] T357;
  wire[8:0] T358;
  wire[8:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire[3:0] T363;
  wire[3:0] T364;
  wire[3:0] T365;
  wire[8:0] T366;
  wire[8:0] T367;
  wire T368;
  wire T369;
  wire T370;
  wire[3:0] T371;
  wire[3:0] T372;
  wire[3:0] T373;
  wire[8:0] T374;
  wire[8:0] T375;
  wire T376;
  wire T377;
  wire T378;
  wire[3:0] T379;
  wire[3:0] T380;
  wire[3:0] T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire T384;
  wire T385;
  wire T386;
  wire[3:0] T387;
  wire[3:0] T388;
  wire[3:0] T389;
  wire[8:0] T390;
  wire[8:0] T391;
  wire T392;
  wire T393;
  wire T394;
  wire[3:0] T395;
  wire[3:0] T396;
  wire[3:0] T397;
  wire[8:0] T398;
  wire[8:0] T399;
  wire T400;
  wire T401;
  wire T402;
  wire[3:0] T403;
  wire[3:0] T404;
  wire[3:0] T405;
  wire[8:0] T406;
  wire[8:0] T407;
  wire T408;
  wire T409;
  wire T410;
  wire[3:0] T411;
  wire[3:0] T412;
  wire[3:0] T413;
  wire[8:0] T414;
  wire[8:0] T415;
  wire T416;
  wire T417;
  wire T418;
  wire[3:0] T419;
  wire[3:0] T420;
  wire[3:0] T421;
  wire[8:0] T422;
  wire[8:0] T423;
  wire T424;
  wire T425;
  wire T426;
  wire[3:0] T427;
  wire[3:0] T428;
  wire[3:0] T429;
  wire[8:0] T430;
  wire[8:0] T431;
  wire T432;
  wire T433;
  wire T434;
  wire[3:0] T435;
  wire[3:0] T436;
  wire[3:0] T437;
  wire[8:0] T438;
  wire[8:0] T439;
  wire T440;
  wire T441;
  wire T442;
  wire[3:0] T443;
  wire[3:0] T444;
  wire[3:0] T445;
  wire[8:0] T446;
  wire[8:0] T447;
  wire T448;
  wire T449;
  wire T450;
  wire[1:0] T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire[2:0] T454;
  wire[2:0] T455;
  wire T456;
  wire T457;
  wire T458;
  wire[1:0] T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire[2:0] T462;
  wire[2:0] T463;
  wire T464;
  wire T465;
  wire T466;
  wire[1:0] T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire[2:0] T470;
  wire[2:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire[1:0] T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire[2:0] T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire[1:0] T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire[2:0] T486;
  wire[2:0] T487;
  wire T488;
  wire T489;
  wire T490;
  wire[1:0] T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire[2:0] T494;
  wire[2:0] T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire T500;
  wire T501;
  wire[1:0] T502;
  wire[1:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire[1:0] T510;
  wire[1:0] T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire[1:0] T518;
  wire[1:0] T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire[1:0] T526;
  wire[1:0] T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire[1:0] T534;
  wire[1:0] T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire[1:0] T542;
  wire[1:0] T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire[1:0] T550;
  wire[1:0] T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire[1:0] T558;
  wire[1:0] T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire[1:0] T566;
  wire[1:0] T567;
  wire T568;
  wire T569;
  wire T570;
  wire[1:0] T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire[2:0] T574;
  wire[2:0] T575;
  wire T576;
  wire T577;
  wire T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire[2:0] T582;
  wire[2:0] T583;
  wire T584;
  wire T585;
  wire T586;
  wire[1:0] T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire[2:0] T590;
  wire[2:0] T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire[2:0] T598;
  wire[2:0] T599;
  wire T600;
  wire T601;
  wire T602;
  wire[1:0] T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire[2:0] T606;
  wire[2:0] T607;
  wire T608;
  wire T609;
  wire T610;
  wire[1:0] T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire[2:0] T614;
  wire[2:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire[1:0] T622;
  wire[1:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire[1:0] T630;
  wire[1:0] T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire[1:0] T638;
  wire[1:0] T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire[1:0] T646;
  wire[1:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire[1:0] T654;
  wire[1:0] T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire[1:0] T662;
  wire[1:0] T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire[1:0] T670;
  wire[1:0] T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire[1:0] T678;
  wire[1:0] T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire[1:0] T686;
  wire[1:0] T687;
  wire T688;
  wire T689;
  wire T690;
  wire[1:0] T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire[2:0] T694;
  wire[2:0] T695;
  wire T696;
  wire T697;
  wire T698;
  wire[1:0] T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire[2:0] T702;
  wire[2:0] T703;
  wire T704;
  wire T705;
  wire T706;
  wire[1:0] T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire[2:0] T710;
  wire[2:0] T711;
  wire T712;
  wire T713;
  wire T714;
  wire[1:0] T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire[2:0] T718;
  wire[2:0] T719;
  wire T720;
  wire T721;
  wire T722;
  wire[1:0] T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire[2:0] T726;
  wire[2:0] T727;
  wire T728;
  wire T729;
  wire T730;
  wire[1:0] T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire[2:0] T734;
  wire[2:0] T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire T740;
  wire T741;
  wire[1:0] T742;
  wire[1:0] T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire[1:0] T750;
  wire[1:0] T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire[1:0] T758;
  wire[1:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire[1:0] T766;
  wire[1:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire[1:0] T774;
  wire[1:0] T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire[1:0] T782;
  wire[1:0] T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire[1:0] T790;
  wire[1:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire[1:0] T798;
  wire[1:0] T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire[1:0] T806;
  wire[1:0] T807;
  wire T808;
  wire T809;
  wire T810;
  wire[3:0] T811;
  wire[3:0] T812;
  wire[3:0] T813;
  wire[10:0] T814;
  wire[10:0] T815;
  wire T816;
  wire T817;
  wire T818;
  wire[1:0] T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire[2:0] T822;
  wire[2:0] T823;
  wire T824;
  wire T825;
  wire T826;
  wire[3:0] T827;
  wire[3:0] T828;
  wire[3:0] T829;
  wire[10:0] T830;
  wire[10:0] T831;
  wire T832;
  wire T833;
  wire T834;
  wire[1:0] T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire[2:0] T838;
  wire[2:0] T839;
  wire T840;
  wire T841;
  wire T842;
  wire[3:0] T843;
  wire[3:0] T844;
  wire[3:0] T845;
  wire[10:0] T846;
  wire[10:0] T847;
  wire T848;
  wire T849;
  wire T850;
  wire[1:0] T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire[2:0] T854;
  wire[2:0] T855;
  wire T856;
  wire T857;
  wire T858;
  wire[3:0] T859;
  wire[3:0] T860;
  wire[3:0] T861;
  wire[10:0] T862;
  wire[10:0] T863;
  wire T864;
  wire T865;
  wire T866;
  wire[1:0] T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire[2:0] T870;
  wire[2:0] T871;
  wire T872;
  wire T873;
  wire T874;
  wire[3:0] T875;
  wire[3:0] T876;
  wire[3:0] T877;
  wire[10:0] T878;
  wire[10:0] T879;
  wire T880;
  wire T881;
  wire T882;
  wire[1:0] T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire[2:0] T886;
  wire[2:0] T887;
  wire T888;
  wire T889;
  wire T890;
  wire[3:0] T891;
  wire[3:0] T892;
  wire[3:0] T893;
  wire[10:0] T894;
  wire[10:0] T895;
  wire T896;
  wire T897;
  wire T898;
  wire[1:0] T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire[2:0] T902;
  wire[2:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire[3:0] T907;
  wire[3:0] T908;
  wire[3:0] T909;
  wire[10:0] T910;
  wire[10:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire[1:0] T918;
  wire[1:0] T919;
  wire T920;
  wire T921;
  wire T922;
  wire[3:0] T923;
  wire[3:0] T924;
  wire[3:0] T925;
  wire[10:0] T926;
  wire[10:0] T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire T932;
  wire T933;
  wire[1:0] T934;
  wire[1:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire[3:0] T939;
  wire[3:0] T940;
  wire[3:0] T941;
  wire[10:0] T942;
  wire[10:0] T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire[1:0] T950;
  wire[1:0] T951;
  wire T952;
  wire T953;
  wire T954;
  wire[3:0] T955;
  wire[3:0] T956;
  wire[3:0] T957;
  wire[9:0] T958;
  wire[9:0] T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire T964;
  wire T965;
  wire[1:0] T966;
  wire[1:0] T967;
  wire T968;
  wire T969;
  wire T970;
  wire[3:0] T971;
  wire[3:0] T972;
  wire[3:0] T973;
  wire[9:0] T974;
  wire[9:0] T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire T980;
  wire T981;
  wire[1:0] T982;
  wire[1:0] T983;
  wire T984;
  wire T985;
  wire T986;
  wire[3:0] T987;
  wire[3:0] T988;
  wire[3:0] T989;
  wire[9:0] T990;
  wire[9:0] T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire[1:0] T998;
  wire[1:0] T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire[3:0] T1003;
  wire[3:0] T1004;
  wire[3:0] T1005;
  wire[9:0] T1006;
  wire[9:0] T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire T1012;
  wire T1013;
  wire[1:0] T1014;
  wire[1:0] T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire[3:0] T1019;
  wire[3:0] T1020;
  wire[3:0] T1021;
  wire[9:0] T1022;
  wire[9:0] T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire[1:0] T1030;
  wire[1:0] T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire[3:0] T1035;
  wire[3:0] T1036;
  wire[3:0] T1037;
  wire[9:0] T1038;
  wire[9:0] T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire T1044;
  wire T1045;
  wire[1:0] T1046;
  wire[1:0] T1047;
  wire[22:0] T1048;
  wire[22:0] T1049;
  wire[21:0] T1050;
  wire[21:0] T1051;
  wire[20:0] T1052;
  wire[20:0] T1053;
  wire[19:0] T1054;
  wire[19:0] T1055;
  wire[18:0] T1056;
  wire[18:0] T1057;
  wire[17:0] T1058;
  wire[17:0] T1059;
  wire[16:0] T1060;
  wire[16:0] T1061;
  wire[15:0] T1062;
  wire[15:0] T1063;
  wire[14:0] T1064;
  wire[14:0] T1065;
  wire[13:0] T1066;
  wire[13:0] T1067;
  wire[12:0] T1068;
  wire[12:0] T1069;
  wire[11:0] T1070;
  wire[11:0] T1071;
  wire[10:0] T1072;
  wire[10:0] T1073;
  wire[9:0] T1074;
  wire[9:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire[7:0] T1078;
  wire[7:0] T1079;
  wire[6:0] T1080;
  wire[6:0] T1081;
  wire[5:0] T1082;
  wire[5:0] T1083;
  wire[4:0] T1084;
  wire[4:0] T1085;
  wire[3:0] T1086;
  wire[3:0] T1087;
  wire[2:0] T1088;
  wire[2:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire[3:0] T1095;
  wire[3:0] T1096;
  wire[3:0] T1097;
  wire[11:0] T1098;
  wire[11:0] T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire[3:0] T1103;
  wire[3:0] T1104;
  wire[3:0] T1105;
  wire[11:0] T1106;
  wire[11:0] T1107;
  wire T1108;
  wire T1109;
  wire T1110;
  wire[3:0] T1111;
  wire[3:0] T1112;
  wire[3:0] T1113;
  wire[11:0] T1114;
  wire[11:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire[3:0] T1119;
  wire[3:0] T1120;
  wire[3:0] T1121;
  wire[11:0] T1122;
  wire[11:0] T1123;
  wire T1124;
  wire T1125;
  wire T1126;
  wire[3:0] T1127;
  wire[3:0] T1128;
  wire[3:0] T1129;
  wire[11:0] T1130;
  wire[11:0] T1131;
  wire T1132;
  wire T1133;
  wire T1134;
  wire[3:0] T1135;
  wire[3:0] T1136;
  wire[3:0] T1137;
  wire[11:0] T1138;
  wire[11:0] T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire[3:0] T1143;
  wire[3:0] T1144;
  wire[3:0] T1145;
  wire[11:0] T1146;
  wire[11:0] T1147;
  wire T1148;
  wire T1149;
  wire T1150;
  wire[3:0] T1151;
  wire[3:0] T1152;
  wire[3:0] T1153;
  wire[11:0] T1154;
  wire[11:0] T1155;
  wire T1156;
  wire T1157;
  wire T1158;
  wire[3:0] T1159;
  wire[3:0] T1160;
  wire[3:0] T1161;
  wire[11:0] T1162;
  wire[11:0] T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire[3:0] T1167;
  wire[3:0] T1168;
  wire[3:0] T1169;
  wire[11:0] T1170;
  wire[11:0] T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire[3:0] T1175;
  wire[3:0] T1176;
  wire[3:0] T1177;
  wire[11:0] T1178;
  wire[11:0] T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire[3:0] T1183;
  wire[3:0] T1184;
  wire[3:0] T1185;
  wire[11:0] T1186;
  wire[11:0] T1187;
  wire T1188;
  wire T1189;
  wire T1190;
  wire[3:0] T1191;
  wire[3:0] T1192;
  wire[3:0] T1193;
  wire[11:0] T1194;
  wire[11:0] T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[3:0] T1199;
  wire[3:0] T1200;
  wire[3:0] T1201;
  wire[11:0] T1202;
  wire[11:0] T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire[3:0] T1207;
  wire[3:0] T1208;
  wire[3:0] T1209;
  wire[11:0] T1210;
  wire[11:0] T1211;
  wire T1212;
  wire T1213;
  wire T1214;
  wire[3:0] T1215;
  wire[3:0] T1216;
  wire[3:0] T1217;
  wire[11:0] T1218;
  wire[11:0] T1219;
  wire T1220;
  wire T1221;
  wire T1222;
  wire[3:0] T1223;
  wire[3:0] T1224;
  wire[3:0] T1225;
  wire[11:0] T1226;
  wire[11:0] T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire[3:0] T1231;
  wire[3:0] T1232;
  wire[3:0] T1233;
  wire[11:0] T1234;
  wire[11:0] T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire[3:0] T1239;
  wire[3:0] T1240;
  wire[3:0] T1241;
  wire[11:0] T1242;
  wire[11:0] T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire[3:0] T1247;
  wire[3:0] T1248;
  wire[3:0] T1249;
  wire[11:0] T1250;
  wire[11:0] T1251;
  wire T1252;
  wire T1253;
  wire T1254;
  wire[3:0] T1255;
  wire[3:0] T1256;
  wire[3:0] T1257;
  wire[11:0] T1258;
  wire[11:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire[3:0] T1263;
  wire[3:0] T1264;
  wire[3:0] T1265;
  wire[11:0] T1266;
  wire[11:0] T1267;
  wire T1268;
  wire T1269;
  wire T1270;
  wire[3:0] T1271;
  wire[3:0] T1272;
  wire[3:0] T1273;
  wire[11:0] T1274;
  wire[11:0] T1275;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1040, T2};
  assign T2 = T3;
  assign T3 = {T1032, T4};
  assign T4 = T5;
  assign T5 = {T1024, T6};
  assign T6 = T7;
  assign T7 = {T1016, T8};
  assign T8 = T9;
  assign T9 = {T1008, T10};
  assign T10 = T11;
  assign T11 = {T1000, T12};
  assign T12 = T13;
  assign T13 = {T992, T14};
  assign T14 = T15;
  assign T15 = {T984, T16};
  assign T16 = T17;
  assign T17 = {T976, T18};
  assign T18 = T19;
  assign T19 = {T968, T20};
  assign T20 = T21;
  assign T21 = {T960, T22};
  assign T22 = T23;
  assign T23 = {T952, T24};
  assign T24 = T25;
  assign T25 = {T944, T26};
  assign T26 = T27;
  assign T27 = {T936, T28};
  assign T28 = T29;
  assign T29 = {T928, T30};
  assign T30 = T31;
  assign T31 = {T920, T32};
  assign T32 = T33;
  assign T33 = {T912, T34};
  assign T34 = T35;
  assign T35 = {T904, T36};
  assign T36 = T37;
  assign T37 = {T896, T38};
  assign T38 = T39;
  assign T39 = {T888, T40};
  assign T40 = T41;
  assign T41 = {T880, T42};
  assign T42 = T43;
  assign T43 = {T872, T44};
  assign T44 = T45;
  assign T45 = {T864, T46};
  assign T46 = T47;
  assign T47 = {T856, T48};
  assign T48 = T49;
  assign T49 = {T848, T50};
  assign T50 = T51;
  assign T51 = {T840, T52};
  assign T52 = T53;
  assign T53 = {T832, T54};
  assign T54 = T55;
  assign T55 = {T824, T56};
  assign T56 = T57;
  assign T57 = {T816, T58};
  assign T58 = T59;
  assign T59 = {T808, T60};
  assign T60 = T61;
  assign T61 = {T800, T62};
  assign T62 = T63;
  assign T63 = {T792, T64};
  assign T64 = T65;
  assign T65 = {T784, T66};
  assign T66 = T67;
  assign T67 = {T776, T68};
  assign T68 = T69;
  assign T69 = {T768, T70};
  assign T70 = T71;
  assign T71 = {T760, T72};
  assign T72 = T73;
  assign T73 = {T752, T74};
  assign T74 = T75;
  assign T75 = {T744, T76};
  assign T76 = T77;
  assign T77 = {T736, T78};
  assign T78 = T79;
  assign T79 = {T728, T80};
  assign T80 = T81;
  assign T81 = {T720, T82};
  assign T82 = T83;
  assign T83 = {T712, T84};
  assign T84 = T85;
  assign T85 = {T704, T86};
  assign T86 = T87;
  assign T87 = {T696, T88};
  assign T88 = T89;
  assign T89 = {T688, T90};
  assign T90 = T91;
  assign T91 = {T680, T92};
  assign T92 = T93;
  assign T93 = {T672, T94};
  assign T94 = T95;
  assign T95 = {T664, T96};
  assign T96 = T97;
  assign T97 = {T656, T98};
  assign T98 = T99;
  assign T99 = {T648, T100};
  assign T100 = T101;
  assign T101 = {T640, T102};
  assign T102 = T103;
  assign T103 = {T632, T104};
  assign T104 = T105;
  assign T105 = {T624, T106};
  assign T106 = T107;
  assign T107 = {T616, T108};
  assign T108 = T109;
  assign T109 = {T608, T110};
  assign T110 = T111;
  assign T111 = {T600, T112};
  assign T112 = T113;
  assign T113 = {T592, T114};
  assign T114 = T115;
  assign T115 = {T584, T116};
  assign T116 = T117;
  assign T117 = {T576, T118};
  assign T118 = T119;
  assign T119 = {T568, T120};
  assign T120 = T121;
  assign T121 = {T560, T122};
  assign T122 = T123;
  assign T123 = {T552, T124};
  assign T124 = T125;
  assign T125 = {T544, T126};
  assign T126 = T127;
  assign T127 = {T536, T128};
  assign T128 = T129;
  assign T129 = {T528, T130};
  assign T130 = T131;
  assign T131 = {T520, T132};
  assign T132 = T133;
  assign T133 = {T512, T134};
  assign T134 = T135;
  assign T135 = {T504, T136};
  assign T136 = T137;
  assign T137 = {T496, T138};
  assign T138 = T139;
  assign T139 = {T488, T140};
  assign T140 = T141;
  assign T141 = {T480, T142};
  assign T142 = T143;
  assign T143 = {T472, T144};
  assign T144 = T145;
  assign T145 = {T464, T146};
  assign T146 = T147;
  assign T147 = {T456, T148};
  assign T148 = T149;
  assign T149 = {T448, T150};
  assign T150 = T151;
  assign T151 = {T440, T152};
  assign T152 = T153;
  assign T153 = {T432, T154};
  assign T154 = T155;
  assign T155 = {T424, T156};
  assign T156 = T157;
  assign T157 = {T416, T158};
  assign T158 = T159;
  assign T159 = {T408, T160};
  assign T160 = T161;
  assign T161 = {T400, T162};
  assign T162 = T163;
  assign T163 = {T392, T164};
  assign T164 = T165;
  assign T165 = {T384, T166};
  assign T166 = T167;
  assign T167 = {T376, T168};
  assign T168 = T169;
  assign T169 = {T368, T170};
  assign T170 = T171;
  assign T171 = {T360, T172};
  assign T172 = T173;
  assign T173 = {T352, T174};
  assign T174 = T175;
  assign T175 = {T344, T176};
  assign T176 = T177;
  assign T177 = {T336, T178};
  assign T178 = T179;
  assign T179 = {T328, T180};
  assign T180 = T181;
  assign T181 = {T320, T182};
  assign T182 = T183;
  assign T183 = {T312, T184};
  assign T184 = T185;
  assign T185 = {T304, T186};
  assign T186 = T187;
  assign T187 = {T296, T188};
  assign T188 = T189;
  assign T189 = {T288, T190};
  assign T190 = T191;
  assign T191 = {T280, T192};
  assign T192 = T193;
  assign T193 = {T272, T194};
  assign T194 = T195;
  assign T195 = {T264, T196};
  assign T196 = T197;
  assign T197 = {T256, T198};
  assign T198 = T199;
  assign T199 = {T248, T200};
  assign T200 = T201;
  assign T201 = {T240, T202};
  assign T202 = T203;
  assign T203 = {T232, T204};
  assign T204 = T205;
  assign T205 = {T224, T206};
  assign T206 = T207;
  assign T207 = {T216, T208};
  assign T208 = T209;
  assign T209 = T210;
  assign T210 = T214[T211];
  assign T211 = T212;
  assign T212 = T213;
  assign T213 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T214 = T215;
  assign T215 = io_chanxy_in[4'h8/* 8*/:1'h0/* 0*/];
  assign T216 = T217;
  assign T217 = T218;
  assign T218 = T222[T219];
  assign T219 = T220;
  assign T220 = T221;
  assign T221 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T222 = T223;
  assign T223 = io_chanxy_in[5'h11/* 17*/:4'h9/* 9*/];
  assign T224 = T225;
  assign T225 = T226;
  assign T226 = T230[T227];
  assign T227 = T228;
  assign T228 = T229;
  assign T229 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T230 = T231;
  assign T231 = io_chanxy_in[5'h1a/* 26*/:5'h12/* 18*/];
  assign T232 = T233;
  assign T233 = T234;
  assign T234 = T238[T235];
  assign T235 = T236;
  assign T236 = T237;
  assign T237 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T238 = T239;
  assign T239 = io_chanxy_in[6'h23/* 35*/:5'h1b/* 27*/];
  assign T240 = T241;
  assign T241 = T242;
  assign T242 = T246[T243];
  assign T243 = T244;
  assign T244 = T245;
  assign T245 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T246 = T247;
  assign T247 = io_chanxy_in[6'h2c/* 44*/:6'h24/* 36*/];
  assign T248 = T249;
  assign T249 = T250;
  assign T250 = T254[T251];
  assign T251 = T252;
  assign T252 = T253;
  assign T253 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T254 = T255;
  assign T255 = io_chanxy_in[6'h35/* 53*/:6'h2d/* 45*/];
  assign T256 = T257;
  assign T257 = T258;
  assign T258 = T262[T259];
  assign T259 = T260;
  assign T260 = T261;
  assign T261 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T262 = T263;
  assign T263 = io_chanxy_in[6'h3e/* 62*/:6'h36/* 54*/];
  assign T264 = T265;
  assign T265 = T266;
  assign T266 = T270[T267];
  assign T267 = T268;
  assign T268 = T269;
  assign T269 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T270 = T271;
  assign T271 = io_chanxy_in[7'h47/* 71*/:6'h3f/* 63*/];
  assign T272 = T273;
  assign T273 = T274;
  assign T274 = T278[T275];
  assign T275 = T276;
  assign T276 = T277;
  assign T277 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T278 = T279;
  assign T279 = io_chanxy_in[7'h50/* 80*/:7'h48/* 72*/];
  assign T280 = T281;
  assign T281 = T282;
  assign T282 = T286[T283];
  assign T283 = T284;
  assign T284 = T285;
  assign T285 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T286 = T287;
  assign T287 = io_chanxy_in[7'h59/* 89*/:7'h51/* 81*/];
  assign T288 = T289;
  assign T289 = T290;
  assign T290 = T294[T291];
  assign T291 = T292;
  assign T292 = T293;
  assign T293 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T294 = T295;
  assign T295 = io_chanxy_in[7'h62/* 98*/:7'h5a/* 90*/];
  assign T296 = T297;
  assign T297 = T298;
  assign T298 = T302[T299];
  assign T299 = T300;
  assign T300 = T301;
  assign T301 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T302 = T303;
  assign T303 = io_chanxy_in[7'h6b/* 107*/:7'h63/* 99*/];
  assign T304 = T305;
  assign T305 = T306;
  assign T306 = T310[T307];
  assign T307 = T308;
  assign T308 = T309;
  assign T309 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T310 = T311;
  assign T311 = io_chanxy_in[7'h74/* 116*/:7'h6c/* 108*/];
  assign T312 = T313;
  assign T313 = T314;
  assign T314 = T318[T315];
  assign T315 = T316;
  assign T316 = T317;
  assign T317 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T318 = T319;
  assign T319 = io_chanxy_in[7'h7d/* 125*/:7'h75/* 117*/];
  assign T320 = T321;
  assign T321 = T322;
  assign T322 = T326[T323];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T326 = T327;
  assign T327 = io_chanxy_in[8'h86/* 134*/:7'h7e/* 126*/];
  assign T328 = T329;
  assign T329 = T330;
  assign T330 = T334[T331];
  assign T331 = T332;
  assign T332 = T333;
  assign T333 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T334 = T335;
  assign T335 = io_chanxy_in[8'h8f/* 143*/:8'h87/* 135*/];
  assign T336 = T337;
  assign T337 = T338;
  assign T338 = T342[T339];
  assign T339 = T340;
  assign T340 = T341;
  assign T341 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T342 = T343;
  assign T343 = io_chanxy_in[8'h98/* 152*/:8'h90/* 144*/];
  assign T344 = T345;
  assign T345 = T346;
  assign T346 = T350[T347];
  assign T347 = T348;
  assign T348 = T349;
  assign T349 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T350 = T351;
  assign T351 = io_chanxy_in[8'ha1/* 161*/:8'h99/* 153*/];
  assign T352 = T353;
  assign T353 = T354;
  assign T354 = T358[T355];
  assign T355 = T356;
  assign T356 = T357;
  assign T357 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T358 = T359;
  assign T359 = io_chanxy_in[8'haa/* 170*/:8'ha2/* 162*/];
  assign T360 = T361;
  assign T361 = T362;
  assign T362 = T366[T363];
  assign T363 = T364;
  assign T364 = T365;
  assign T365 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T366 = T367;
  assign T367 = io_chanxy_in[8'hb3/* 179*/:8'hab/* 171*/];
  assign T368 = T369;
  assign T369 = T370;
  assign T370 = T374[T371];
  assign T371 = T372;
  assign T372 = T373;
  assign T373 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T374 = T375;
  assign T375 = io_chanxy_in[8'hbc/* 188*/:8'hb4/* 180*/];
  assign T376 = T377;
  assign T377 = T378;
  assign T378 = T382[T379];
  assign T379 = T380;
  assign T380 = T381;
  assign T381 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T382 = T383;
  assign T383 = io_chanxy_in[8'hc5/* 197*/:8'hbd/* 189*/];
  assign T384 = T385;
  assign T385 = T386;
  assign T386 = T390[T387];
  assign T387 = T388;
  assign T388 = T389;
  assign T389 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T390 = T391;
  assign T391 = io_chanxy_in[8'hce/* 206*/:8'hc6/* 198*/];
  assign T392 = T393;
  assign T393 = T394;
  assign T394 = T398[T395];
  assign T395 = T396;
  assign T396 = T397;
  assign T397 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T398 = T399;
  assign T399 = io_chanxy_in[8'hd7/* 215*/:8'hcf/* 207*/];
  assign T400 = T401;
  assign T401 = T402;
  assign T402 = T406[T403];
  assign T403 = T404;
  assign T404 = T405;
  assign T405 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T406 = T407;
  assign T407 = io_chanxy_in[8'he0/* 224*/:8'hd8/* 216*/];
  assign T408 = T409;
  assign T409 = T410;
  assign T410 = T414[T411];
  assign T411 = T412;
  assign T412 = T413;
  assign T413 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T414 = T415;
  assign T415 = io_chanxy_in[8'he9/* 233*/:8'he1/* 225*/];
  assign T416 = T417;
  assign T417 = T418;
  assign T418 = T422[T419];
  assign T419 = T420;
  assign T420 = T421;
  assign T421 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T422 = T423;
  assign T423 = io_chanxy_in[8'hf2/* 242*/:8'hea/* 234*/];
  assign T424 = T425;
  assign T425 = T426;
  assign T426 = T430[T427];
  assign T427 = T428;
  assign T428 = T429;
  assign T429 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T430 = T431;
  assign T431 = io_chanxy_in[8'hfb/* 251*/:8'hf3/* 243*/];
  assign T432 = T433;
  assign T433 = T434;
  assign T434 = T438[T435];
  assign T435 = T436;
  assign T436 = T437;
  assign T437 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T438 = T439;
  assign T439 = io_chanxy_in[9'h104/* 260*/:8'hfc/* 252*/];
  assign T440 = T441;
  assign T441 = T442;
  assign T442 = T446[T443];
  assign T443 = T444;
  assign T444 = T445;
  assign T445 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T446 = T447;
  assign T447 = io_chanxy_in[9'h10d/* 269*/:9'h105/* 261*/];
  assign T448 = T449;
  assign T449 = T450;
  assign T450 = T454[T451];
  assign T451 = T452;
  assign T452 = T453;
  assign T453 = io_chanxy_config[7'h79/* 121*/:7'h78/* 120*/];
  assign T454 = T455;
  assign T455 = io_chanxy_in[9'h110/* 272*/:9'h10e/* 270*/];
  assign T456 = T457;
  assign T457 = T458;
  assign T458 = T462[T459];
  assign T459 = T460;
  assign T460 = T461;
  assign T461 = io_chanxy_config[7'h7b/* 123*/:7'h7a/* 122*/];
  assign T462 = T463;
  assign T463 = io_chanxy_in[9'h113/* 275*/:9'h111/* 273*/];
  assign T464 = T465;
  assign T465 = T466;
  assign T466 = T470[T467];
  assign T467 = T468;
  assign T468 = T469;
  assign T469 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T470 = T471;
  assign T471 = io_chanxy_in[9'h116/* 278*/:9'h114/* 276*/];
  assign T472 = T473;
  assign T473 = T474;
  assign T474 = T478[T475];
  assign T475 = T476;
  assign T476 = T477;
  assign T477 = io_chanxy_config[7'h7f/* 127*/:7'h7e/* 126*/];
  assign T478 = T479;
  assign T479 = io_chanxy_in[9'h119/* 281*/:9'h117/* 279*/];
  assign T480 = T481;
  assign T481 = T482;
  assign T482 = T486[T483];
  assign T483 = T484;
  assign T484 = T485;
  assign T485 = io_chanxy_config[8'h81/* 129*/:8'h80/* 128*/];
  assign T486 = T487;
  assign T487 = io_chanxy_in[9'h11c/* 284*/:9'h11a/* 282*/];
  assign T488 = T489;
  assign T489 = T490;
  assign T490 = T494[T491];
  assign T491 = T492;
  assign T492 = T493;
  assign T493 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T494 = T495;
  assign T495 = io_chanxy_in[9'h11f/* 287*/:9'h11d/* 285*/];
  assign T496 = T497;
  assign T497 = T498;
  assign T498 = T502[T499];
  assign T499 = T500;
  assign T500 = T501;
  assign T501 = io_chanxy_config[8'h84/* 132*/:8'h84/* 132*/];
  assign T502 = T503;
  assign T503 = io_chanxy_in[9'h121/* 289*/:9'h120/* 288*/];
  assign T504 = T505;
  assign T505 = T506;
  assign T506 = T510[T507];
  assign T507 = T508;
  assign T508 = T509;
  assign T509 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T510 = T511;
  assign T511 = io_chanxy_in[9'h123/* 291*/:9'h122/* 290*/];
  assign T512 = T513;
  assign T513 = T514;
  assign T514 = T518[T515];
  assign T515 = T516;
  assign T516 = T517;
  assign T517 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T518 = T519;
  assign T519 = io_chanxy_in[9'h125/* 293*/:9'h124/* 292*/];
  assign T520 = T521;
  assign T521 = T522;
  assign T522 = T526[T523];
  assign T523 = T524;
  assign T524 = T525;
  assign T525 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T526 = T527;
  assign T527 = io_chanxy_in[9'h127/* 295*/:9'h126/* 294*/];
  assign T528 = T529;
  assign T529 = T530;
  assign T530 = T534[T531];
  assign T531 = T532;
  assign T532 = T533;
  assign T533 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T534 = T535;
  assign T535 = io_chanxy_in[9'h129/* 297*/:9'h128/* 296*/];
  assign T536 = T537;
  assign T537 = T538;
  assign T538 = T542[T539];
  assign T539 = T540;
  assign T540 = T541;
  assign T541 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T542 = T543;
  assign T543 = io_chanxy_in[9'h12b/* 299*/:9'h12a/* 298*/];
  assign T544 = T545;
  assign T545 = T546;
  assign T546 = T550[T547];
  assign T547 = T548;
  assign T548 = T549;
  assign T549 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T550 = T551;
  assign T551 = io_chanxy_in[9'h12d/* 301*/:9'h12c/* 300*/];
  assign T552 = T553;
  assign T553 = T554;
  assign T554 = T558[T555];
  assign T555 = T556;
  assign T556 = T557;
  assign T557 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T558 = T559;
  assign T559 = io_chanxy_in[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T560 = T561;
  assign T561 = T562;
  assign T562 = T566[T563];
  assign T563 = T564;
  assign T564 = T565;
  assign T565 = io_chanxy_config[8'h8c/* 140*/:8'h8c/* 140*/];
  assign T566 = T567;
  assign T567 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T568 = T569;
  assign T569 = T570;
  assign T570 = T574[T571];
  assign T571 = T572;
  assign T572 = T573;
  assign T573 = io_chanxy_config[8'h8e/* 142*/:8'h8d/* 141*/];
  assign T574 = T575;
  assign T575 = io_chanxy_in[9'h134/* 308*/:9'h132/* 306*/];
  assign T576 = T577;
  assign T577 = T578;
  assign T578 = T582[T579];
  assign T579 = T580;
  assign T580 = T581;
  assign T581 = io_chanxy_config[8'h90/* 144*/:8'h8f/* 143*/];
  assign T582 = T583;
  assign T583 = io_chanxy_in[9'h137/* 311*/:9'h135/* 309*/];
  assign T584 = T585;
  assign T585 = T586;
  assign T586 = T590[T587];
  assign T587 = T588;
  assign T588 = T589;
  assign T589 = io_chanxy_config[8'h92/* 146*/:8'h91/* 145*/];
  assign T590 = T591;
  assign T591 = io_chanxy_in[9'h13a/* 314*/:9'h138/* 312*/];
  assign T592 = T593;
  assign T593 = T594;
  assign T594 = T598[T595];
  assign T595 = T596;
  assign T596 = T597;
  assign T597 = io_chanxy_config[8'h94/* 148*/:8'h93/* 147*/];
  assign T598 = T599;
  assign T599 = io_chanxy_in[9'h13d/* 317*/:9'h13b/* 315*/];
  assign T600 = T601;
  assign T601 = T602;
  assign T602 = T606[T603];
  assign T603 = T604;
  assign T604 = T605;
  assign T605 = io_chanxy_config[8'h96/* 150*/:8'h95/* 149*/];
  assign T606 = T607;
  assign T607 = io_chanxy_in[9'h140/* 320*/:9'h13e/* 318*/];
  assign T608 = T609;
  assign T609 = T610;
  assign T610 = T614[T611];
  assign T611 = T612;
  assign T612 = T613;
  assign T613 = io_chanxy_config[8'h98/* 152*/:8'h97/* 151*/];
  assign T614 = T615;
  assign T615 = io_chanxy_in[9'h143/* 323*/:9'h141/* 321*/];
  assign T616 = T617;
  assign T617 = T618;
  assign T618 = T622[T619];
  assign T619 = T620;
  assign T620 = T621;
  assign T621 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T622 = T623;
  assign T623 = io_chanxy_in[9'h145/* 325*/:9'h144/* 324*/];
  assign T624 = T625;
  assign T625 = T626;
  assign T626 = T630[T627];
  assign T627 = T628;
  assign T628 = T629;
  assign T629 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T630 = T631;
  assign T631 = io_chanxy_in[9'h147/* 327*/:9'h146/* 326*/];
  assign T632 = T633;
  assign T633 = T634;
  assign T634 = T638[T635];
  assign T635 = T636;
  assign T636 = T637;
  assign T637 = io_chanxy_config[8'h9b/* 155*/:8'h9b/* 155*/];
  assign T638 = T639;
  assign T639 = io_chanxy_in[9'h149/* 329*/:9'h148/* 328*/];
  assign T640 = T641;
  assign T641 = T642;
  assign T642 = T646[T643];
  assign T643 = T644;
  assign T644 = T645;
  assign T645 = io_chanxy_config[8'h9c/* 156*/:8'h9c/* 156*/];
  assign T646 = T647;
  assign T647 = io_chanxy_in[9'h14b/* 331*/:9'h14a/* 330*/];
  assign T648 = T649;
  assign T649 = T650;
  assign T650 = T654[T651];
  assign T651 = T652;
  assign T652 = T653;
  assign T653 = io_chanxy_config[8'h9d/* 157*/:8'h9d/* 157*/];
  assign T654 = T655;
  assign T655 = io_chanxy_in[9'h14d/* 333*/:9'h14c/* 332*/];
  assign T656 = T657;
  assign T657 = T658;
  assign T658 = T662[T659];
  assign T659 = T660;
  assign T660 = T661;
  assign T661 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T662 = T663;
  assign T663 = io_chanxy_in[9'h14f/* 335*/:9'h14e/* 334*/];
  assign T664 = T665;
  assign T665 = T666;
  assign T666 = T670[T667];
  assign T667 = T668;
  assign T668 = T669;
  assign T669 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T670 = T671;
  assign T671 = io_chanxy_in[9'h151/* 337*/:9'h150/* 336*/];
  assign T672 = T673;
  assign T673 = T674;
  assign T674 = T678[T675];
  assign T675 = T676;
  assign T676 = T677;
  assign T677 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T678 = T679;
  assign T679 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign T680 = T681;
  assign T681 = T682;
  assign T682 = T686[T683];
  assign T683 = T684;
  assign T684 = T685;
  assign T685 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T686 = T687;
  assign T687 = io_chanxy_in[9'h155/* 341*/:9'h154/* 340*/];
  assign T688 = T689;
  assign T689 = T690;
  assign T690 = T694[T691];
  assign T691 = T692;
  assign T692 = T693;
  assign T693 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T694 = T695;
  assign T695 = io_chanxy_in[9'h158/* 344*/:9'h156/* 342*/];
  assign T696 = T697;
  assign T697 = T698;
  assign T698 = T702[T699];
  assign T699 = T700;
  assign T700 = T701;
  assign T701 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T702 = T703;
  assign T703 = io_chanxy_in[9'h15b/* 347*/:9'h159/* 345*/];
  assign T704 = T705;
  assign T705 = T706;
  assign T706 = T710[T707];
  assign T707 = T708;
  assign T708 = T709;
  assign T709 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T710 = T711;
  assign T711 = io_chanxy_in[9'h15e/* 350*/:9'h15c/* 348*/];
  assign T712 = T713;
  assign T713 = T714;
  assign T714 = T718[T715];
  assign T715 = T716;
  assign T716 = T717;
  assign T717 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T718 = T719;
  assign T719 = io_chanxy_in[9'h161/* 353*/:9'h15f/* 351*/];
  assign T720 = T721;
  assign T721 = T722;
  assign T722 = T726[T723];
  assign T723 = T724;
  assign T724 = T725;
  assign T725 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T726 = T727;
  assign T727 = io_chanxy_in[9'h164/* 356*/:9'h162/* 354*/];
  assign T728 = T729;
  assign T729 = T730;
  assign T730 = T734[T731];
  assign T731 = T732;
  assign T732 = T733;
  assign T733 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T734 = T735;
  assign T735 = io_chanxy_in[9'h167/* 359*/:9'h165/* 357*/];
  assign T736 = T737;
  assign T737 = T738;
  assign T738 = T742[T739];
  assign T739 = T740;
  assign T740 = T741;
  assign T741 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T742 = T743;
  assign T743 = io_chanxy_in[9'h169/* 361*/:9'h168/* 360*/];
  assign T744 = T745;
  assign T745 = T746;
  assign T746 = T750[T747];
  assign T747 = T748;
  assign T748 = T749;
  assign T749 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T750 = T751;
  assign T751 = io_chanxy_in[9'h16b/* 363*/:9'h16a/* 362*/];
  assign T752 = T753;
  assign T753 = T754;
  assign T754 = T758[T755];
  assign T755 = T756;
  assign T756 = T757;
  assign T757 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T758 = T759;
  assign T759 = io_chanxy_in[9'h16d/* 365*/:9'h16c/* 364*/];
  assign T760 = T761;
  assign T761 = T762;
  assign T762 = T766[T763];
  assign T763 = T764;
  assign T764 = T765;
  assign T765 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T766 = T767;
  assign T767 = io_chanxy_in[9'h16f/* 367*/:9'h16e/* 366*/];
  assign T768 = T769;
  assign T769 = T770;
  assign T770 = T774[T771];
  assign T771 = T772;
  assign T772 = T773;
  assign T773 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T774 = T775;
  assign T775 = io_chanxy_in[9'h171/* 369*/:9'h170/* 368*/];
  assign T776 = T777;
  assign T777 = T778;
  assign T778 = T782[T779];
  assign T779 = T780;
  assign T780 = T781;
  assign T781 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T782 = T783;
  assign T783 = io_chanxy_in[9'h173/* 371*/:9'h172/* 370*/];
  assign T784 = T785;
  assign T785 = T786;
  assign T786 = T790[T787];
  assign T787 = T788;
  assign T788 = T789;
  assign T789 = io_chanxy_config[8'hb4/* 180*/:8'hb4/* 180*/];
  assign T790 = T791;
  assign T791 = io_chanxy_in[9'h175/* 373*/:9'h174/* 372*/];
  assign T792 = T793;
  assign T793 = T794;
  assign T794 = T798[T795];
  assign T795 = T796;
  assign T796 = T797;
  assign T797 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T798 = T799;
  assign T799 = io_chanxy_in[9'h177/* 375*/:9'h176/* 374*/];
  assign T800 = T801;
  assign T801 = T802;
  assign T802 = T806[T803];
  assign T803 = T804;
  assign T804 = T805;
  assign T805 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T806 = T807;
  assign T807 = io_chanxy_in[9'h179/* 377*/:9'h178/* 376*/];
  assign T808 = T809;
  assign T809 = T810;
  assign T810 = T814[T811];
  assign T811 = T812;
  assign T812 = T813;
  assign T813 = io_chanxy_config[8'hba/* 186*/:8'hb7/* 183*/];
  assign T814 = T815;
  assign T815 = io_chanxy_in[9'h184/* 388*/:9'h17a/* 378*/];
  assign T816 = T817;
  assign T817 = T818;
  assign T818 = T822[T819];
  assign T819 = T820;
  assign T820 = T821;
  assign T821 = io_chanxy_config[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T822 = T823;
  assign T823 = io_chanxy_in[9'h187/* 391*/:9'h185/* 389*/];
  assign T824 = T825;
  assign T825 = T826;
  assign T826 = T830[T827];
  assign T827 = T828;
  assign T828 = T829;
  assign T829 = io_chanxy_config[8'hc0/* 192*/:8'hbd/* 189*/];
  assign T830 = T831;
  assign T831 = io_chanxy_in[9'h192/* 402*/:9'h188/* 392*/];
  assign T832 = T833;
  assign T833 = T834;
  assign T834 = T838[T835];
  assign T835 = T836;
  assign T836 = T837;
  assign T837 = io_chanxy_config[8'hc2/* 194*/:8'hc1/* 193*/];
  assign T838 = T839;
  assign T839 = io_chanxy_in[9'h195/* 405*/:9'h193/* 403*/];
  assign T840 = T841;
  assign T841 = T842;
  assign T842 = T846[T843];
  assign T843 = T844;
  assign T844 = T845;
  assign T845 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T846 = T847;
  assign T847 = io_chanxy_in[9'h1a0/* 416*/:9'h196/* 406*/];
  assign T848 = T849;
  assign T849 = T850;
  assign T850 = T854[T851];
  assign T851 = T852;
  assign T852 = T853;
  assign T853 = io_chanxy_config[8'hc8/* 200*/:8'hc7/* 199*/];
  assign T854 = T855;
  assign T855 = io_chanxy_in[9'h1a3/* 419*/:9'h1a1/* 417*/];
  assign T856 = T857;
  assign T857 = T858;
  assign T858 = T862[T859];
  assign T859 = T860;
  assign T860 = T861;
  assign T861 = io_chanxy_config[8'hcc/* 204*/:8'hc9/* 201*/];
  assign T862 = T863;
  assign T863 = io_chanxy_in[9'h1ae/* 430*/:9'h1a4/* 420*/];
  assign T864 = T865;
  assign T865 = T866;
  assign T866 = T870[T867];
  assign T867 = T868;
  assign T868 = T869;
  assign T869 = io_chanxy_config[8'hce/* 206*/:8'hcd/* 205*/];
  assign T870 = T871;
  assign T871 = io_chanxy_in[9'h1b1/* 433*/:9'h1af/* 431*/];
  assign T872 = T873;
  assign T873 = T874;
  assign T874 = T878[T875];
  assign T875 = T876;
  assign T876 = T877;
  assign T877 = io_chanxy_config[8'hd2/* 210*/:8'hcf/* 207*/];
  assign T878 = T879;
  assign T879 = io_chanxy_in[9'h1bc/* 444*/:9'h1b2/* 434*/];
  assign T880 = T881;
  assign T881 = T882;
  assign T882 = T886[T883];
  assign T883 = T884;
  assign T884 = T885;
  assign T885 = io_chanxy_config[8'hd4/* 212*/:8'hd3/* 211*/];
  assign T886 = T887;
  assign T887 = io_chanxy_in[9'h1bf/* 447*/:9'h1bd/* 445*/];
  assign T888 = T889;
  assign T889 = T890;
  assign T890 = T894[T891];
  assign T891 = T892;
  assign T892 = T893;
  assign T893 = io_chanxy_config[8'hd8/* 216*/:8'hd5/* 213*/];
  assign T894 = T895;
  assign T895 = io_chanxy_in[9'h1ca/* 458*/:9'h1c0/* 448*/];
  assign T896 = T897;
  assign T897 = T898;
  assign T898 = T902[T899];
  assign T899 = T900;
  assign T900 = T901;
  assign T901 = io_chanxy_config[8'hda/* 218*/:8'hd9/* 217*/];
  assign T902 = T903;
  assign T903 = io_chanxy_in[9'h1cd/* 461*/:9'h1cb/* 459*/];
  assign T904 = T905;
  assign T905 = T906;
  assign T906 = T910[T907];
  assign T907 = T908;
  assign T908 = T909;
  assign T909 = io_chanxy_config[8'hde/* 222*/:8'hdb/* 219*/];
  assign T910 = T911;
  assign T911 = io_chanxy_in[9'h1d8/* 472*/:9'h1ce/* 462*/];
  assign T912 = T913;
  assign T913 = T914;
  assign T914 = T918[T915];
  assign T915 = T916;
  assign T916 = T917;
  assign T917 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T918 = T919;
  assign T919 = io_chanxy_in[9'h1da/* 474*/:9'h1d9/* 473*/];
  assign T920 = T921;
  assign T921 = T922;
  assign T922 = T926[T923];
  assign T923 = T924;
  assign T924 = T925;
  assign T925 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T926 = T927;
  assign T927 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T928 = T929;
  assign T929 = T930;
  assign T930 = T934[T931];
  assign T931 = T932;
  assign T932 = T933;
  assign T933 = io_chanxy_config[8'he4/* 228*/:8'he4/* 228*/];
  assign T934 = T935;
  assign T935 = io_chanxy_in[9'h1e7/* 487*/:9'h1e6/* 486*/];
  assign T936 = T937;
  assign T937 = T938;
  assign T938 = T942[T939];
  assign T939 = T940;
  assign T940 = T941;
  assign T941 = io_chanxy_config[8'he8/* 232*/:8'he5/* 229*/];
  assign T942 = T943;
  assign T943 = io_chanxy_in[9'h1f2/* 498*/:9'h1e8/* 488*/];
  assign T944 = T945;
  assign T945 = T946;
  assign T946 = T950[T947];
  assign T947 = T948;
  assign T948 = T949;
  assign T949 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T950 = T951;
  assign T951 = io_chanxy_in[9'h1f4/* 500*/:9'h1f3/* 499*/];
  assign T952 = T953;
  assign T953 = T954;
  assign T954 = T958[T955];
  assign T955 = T956;
  assign T956 = T957;
  assign T957 = io_chanxy_config[8'hed/* 237*/:8'hea/* 234*/];
  assign T958 = T959;
  assign T959 = io_chanxy_in[9'h1fe/* 510*/:9'h1f5/* 501*/];
  assign T960 = T961;
  assign T961 = T962;
  assign T962 = T966[T963];
  assign T963 = T964;
  assign T964 = T965;
  assign T965 = io_chanxy_config[8'hee/* 238*/:8'hee/* 238*/];
  assign T966 = T967;
  assign T967 = io_chanxy_in[10'h200/* 512*/:9'h1ff/* 511*/];
  assign T968 = T969;
  assign T969 = T970;
  assign T970 = T974[T971];
  assign T971 = T972;
  assign T972 = T973;
  assign T973 = io_chanxy_config[8'hf2/* 242*/:8'hef/* 239*/];
  assign T974 = T975;
  assign T975 = io_chanxy_in[10'h20a/* 522*/:10'h201/* 513*/];
  assign T976 = T977;
  assign T977 = T978;
  assign T978 = T982[T979];
  assign T979 = T980;
  assign T980 = T981;
  assign T981 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T982 = T983;
  assign T983 = io_chanxy_in[10'h20c/* 524*/:10'h20b/* 523*/];
  assign T984 = T985;
  assign T985 = T986;
  assign T986 = T990[T987];
  assign T987 = T988;
  assign T988 = T989;
  assign T989 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T990 = T991;
  assign T991 = io_chanxy_in[10'h216/* 534*/:10'h20d/* 525*/];
  assign T992 = T993;
  assign T993 = T994;
  assign T994 = T998[T995];
  assign T995 = T996;
  assign T996 = T997;
  assign T997 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T998 = T999;
  assign T999 = io_chanxy_in[10'h218/* 536*/:10'h217/* 535*/];
  assign T1000 = T1001;
  assign T1001 = T1002;
  assign T1002 = T1006[T1003];
  assign T1003 = T1004;
  assign T1004 = T1005;
  assign T1005 = io_chanxy_config[8'hfc/* 252*/:8'hf9/* 249*/];
  assign T1006 = T1007;
  assign T1007 = io_chanxy_in[10'h222/* 546*/:10'h219/* 537*/];
  assign T1008 = T1009;
  assign T1009 = T1010;
  assign T1010 = T1014[T1011];
  assign T1011 = T1012;
  assign T1012 = T1013;
  assign T1013 = io_chanxy_config[8'hfd/* 253*/:8'hfd/* 253*/];
  assign T1014 = T1015;
  assign T1015 = io_chanxy_in[10'h224/* 548*/:10'h223/* 547*/];
  assign T1016 = T1017;
  assign T1017 = T1018;
  assign T1018 = T1022[T1019];
  assign T1019 = T1020;
  assign T1020 = T1021;
  assign T1021 = io_chanxy_config[9'h101/* 257*/:8'hfe/* 254*/];
  assign T1022 = T1023;
  assign T1023 = io_chanxy_in[10'h22e/* 558*/:10'h225/* 549*/];
  assign T1024 = T1025;
  assign T1025 = T1026;
  assign T1026 = T1030[T1027];
  assign T1027 = T1028;
  assign T1028 = T1029;
  assign T1029 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1030 = T1031;
  assign T1031 = io_chanxy_in[10'h230/* 560*/:10'h22f/* 559*/];
  assign T1032 = T1033;
  assign T1033 = T1034;
  assign T1034 = T1038[T1035];
  assign T1035 = T1036;
  assign T1036 = T1037;
  assign T1037 = io_chanxy_config[9'h106/* 262*/:9'h103/* 259*/];
  assign T1038 = T1039;
  assign T1039 = io_chanxy_in[10'h23a/* 570*/:10'h231/* 561*/];
  assign T1040 = T1041;
  assign T1041 = T1042;
  assign T1042 = T1046[T1043];
  assign T1043 = T1044;
  assign T1044 = T1045;
  assign T1045 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1046 = T1047;
  assign T1047 = io_chanxy_in[10'h23c/* 572*/:10'h23b/* 571*/];
  assign io_ipin_out = T1048;
  assign T1048 = T1049;
  assign T1049 = {T1268, T1050};
  assign T1050 = T1051;
  assign T1051 = {T1260, T1052};
  assign T1052 = T1053;
  assign T1053 = {T1252, T1054};
  assign T1054 = T1055;
  assign T1055 = {T1244, T1056};
  assign T1056 = T1057;
  assign T1057 = {T1236, T1058};
  assign T1058 = T1059;
  assign T1059 = {T1228, T1060};
  assign T1060 = T1061;
  assign T1061 = {T1220, T1062};
  assign T1062 = T1063;
  assign T1063 = {T1212, T1064};
  assign T1064 = T1065;
  assign T1065 = {T1204, T1066};
  assign T1066 = T1067;
  assign T1067 = {T1196, T1068};
  assign T1068 = T1069;
  assign T1069 = {T1188, T1070};
  assign T1070 = T1071;
  assign T1071 = {T1180, T1072};
  assign T1072 = T1073;
  assign T1073 = {T1172, T1074};
  assign T1074 = T1075;
  assign T1075 = {T1164, T1076};
  assign T1076 = T1077;
  assign T1077 = {T1156, T1078};
  assign T1078 = T1079;
  assign T1079 = {T1148, T1080};
  assign T1080 = T1081;
  assign T1081 = {T1140, T1082};
  assign T1082 = T1083;
  assign T1083 = {T1132, T1084};
  assign T1084 = T1085;
  assign T1085 = {T1124, T1086};
  assign T1086 = T1087;
  assign T1087 = {T1116, T1088};
  assign T1088 = T1089;
  assign T1089 = {T1108, T1090};
  assign T1090 = T1091;
  assign T1091 = {T1100, T1092};
  assign T1092 = T1093;
  assign T1093 = T1094;
  assign T1094 = T1098[T1095];
  assign T1095 = T1096;
  assign T1096 = T1097;
  assign T1097 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1098 = T1099;
  assign T1099 = io_ipin_in[4'hb/* 11*/:1'h0/* 0*/];
  assign T1100 = T1101;
  assign T1101 = T1102;
  assign T1102 = T1106[T1103];
  assign T1103 = T1104;
  assign T1104 = T1105;
  assign T1105 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1106 = T1107;
  assign T1107 = io_ipin_in[5'h17/* 23*/:4'hc/* 12*/];
  assign T1108 = T1109;
  assign T1109 = T1110;
  assign T1110 = T1114[T1111];
  assign T1111 = T1112;
  assign T1112 = T1113;
  assign T1113 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1114 = T1115;
  assign T1115 = io_ipin_in[6'h23/* 35*/:5'h18/* 24*/];
  assign T1116 = T1117;
  assign T1117 = T1118;
  assign T1118 = T1122[T1119];
  assign T1119 = T1120;
  assign T1120 = T1121;
  assign T1121 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1122 = T1123;
  assign T1123 = io_ipin_in[6'h2f/* 47*/:6'h24/* 36*/];
  assign T1124 = T1125;
  assign T1125 = T1126;
  assign T1126 = T1130[T1127];
  assign T1127 = T1128;
  assign T1128 = T1129;
  assign T1129 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1130 = T1131;
  assign T1131 = io_ipin_in[6'h3b/* 59*/:6'h30/* 48*/];
  assign T1132 = T1133;
  assign T1133 = T1134;
  assign T1134 = T1138[T1135];
  assign T1135 = T1136;
  assign T1136 = T1137;
  assign T1137 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1138 = T1139;
  assign T1139 = io_ipin_in[7'h47/* 71*/:6'h3c/* 60*/];
  assign T1140 = T1141;
  assign T1141 = T1142;
  assign T1142 = T1146[T1143];
  assign T1143 = T1144;
  assign T1144 = T1145;
  assign T1145 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1146 = T1147;
  assign T1147 = io_ipin_in[7'h53/* 83*/:7'h48/* 72*/];
  assign T1148 = T1149;
  assign T1149 = T1150;
  assign T1150 = T1154[T1151];
  assign T1151 = T1152;
  assign T1152 = T1153;
  assign T1153 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1154 = T1155;
  assign T1155 = io_ipin_in[7'h5f/* 95*/:7'h54/* 84*/];
  assign T1156 = T1157;
  assign T1157 = T1158;
  assign T1158 = T1162[T1159];
  assign T1159 = T1160;
  assign T1160 = T1161;
  assign T1161 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1162 = T1163;
  assign T1163 = io_ipin_in[7'h6b/* 107*/:7'h60/* 96*/];
  assign T1164 = T1165;
  assign T1165 = T1166;
  assign T1166 = T1170[T1167];
  assign T1167 = T1168;
  assign T1168 = T1169;
  assign T1169 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1170 = T1171;
  assign T1171 = io_ipin_in[7'h77/* 119*/:7'h6c/* 108*/];
  assign T1172 = T1173;
  assign T1173 = T1174;
  assign T1174 = T1178[T1175];
  assign T1175 = T1176;
  assign T1176 = T1177;
  assign T1177 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1178 = T1179;
  assign T1179 = io_ipin_in[8'h83/* 131*/:7'h78/* 120*/];
  assign T1180 = T1181;
  assign T1181 = T1182;
  assign T1182 = T1186[T1183];
  assign T1183 = T1184;
  assign T1184 = T1185;
  assign T1185 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1186 = T1187;
  assign T1187 = io_ipin_in[8'h8f/* 143*/:8'h84/* 132*/];
  assign T1188 = T1189;
  assign T1189 = T1190;
  assign T1190 = T1194[T1191];
  assign T1191 = T1192;
  assign T1192 = T1193;
  assign T1193 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1194 = T1195;
  assign T1195 = io_ipin_in[8'h9b/* 155*/:8'h90/* 144*/];
  assign T1196 = T1197;
  assign T1197 = T1198;
  assign T1198 = T1202[T1199];
  assign T1199 = T1200;
  assign T1200 = T1201;
  assign T1201 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1202 = T1203;
  assign T1203 = io_ipin_in[8'ha7/* 167*/:8'h9c/* 156*/];
  assign T1204 = T1205;
  assign T1205 = T1206;
  assign T1206 = T1210[T1207];
  assign T1207 = T1208;
  assign T1208 = T1209;
  assign T1209 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1210 = T1211;
  assign T1211 = io_ipin_in[8'hb3/* 179*/:8'ha8/* 168*/];
  assign T1212 = T1213;
  assign T1213 = T1214;
  assign T1214 = T1218[T1215];
  assign T1215 = T1216;
  assign T1216 = T1217;
  assign T1217 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1218 = T1219;
  assign T1219 = io_ipin_in[8'hbf/* 191*/:8'hb4/* 180*/];
  assign T1220 = T1221;
  assign T1221 = T1222;
  assign T1222 = T1226[T1223];
  assign T1223 = T1224;
  assign T1224 = T1225;
  assign T1225 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1226 = T1227;
  assign T1227 = io_ipin_in[8'hcb/* 203*/:8'hc0/* 192*/];
  assign T1228 = T1229;
  assign T1229 = T1230;
  assign T1230 = T1234[T1231];
  assign T1231 = T1232;
  assign T1232 = T1233;
  assign T1233 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1234 = T1235;
  assign T1235 = io_ipin_in[8'hd7/* 215*/:8'hcc/* 204*/];
  assign T1236 = T1237;
  assign T1237 = T1238;
  assign T1238 = T1242[T1239];
  assign T1239 = T1240;
  assign T1240 = T1241;
  assign T1241 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1242 = T1243;
  assign T1243 = io_ipin_in[8'he3/* 227*/:8'hd8/* 216*/];
  assign T1244 = T1245;
  assign T1245 = T1246;
  assign T1246 = T1250[T1247];
  assign T1247 = T1248;
  assign T1248 = T1249;
  assign T1249 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1250 = T1251;
  assign T1251 = io_ipin_in[8'hef/* 239*/:8'he4/* 228*/];
  assign T1252 = T1253;
  assign T1253 = T1254;
  assign T1254 = T1258[T1255];
  assign T1255 = T1256;
  assign T1256 = T1257;
  assign T1257 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1258 = T1259;
  assign T1259 = io_ipin_in[8'hfb/* 251*/:8'hf0/* 240*/];
  assign T1260 = T1261;
  assign T1261 = T1262;
  assign T1262 = T1266[T1263];
  assign T1263 = T1264;
  assign T1264 = T1265;
  assign T1265 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1266 = T1267;
  assign T1267 = io_ipin_in[9'h107/* 263*/:8'hfc/* 252*/];
  assign T1268 = T1269;
  assign T1269 = T1270;
  assign T1270 = T1274[T1271];
  assign T1271 = T1272;
  assign T1272 = T1273;
  assign T1273 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1274 = T1275;
  assign T1275 = io_ipin_in[9'h113/* 275*/:9'h108/* 264*/];
endmodule

module lut_tile_sp_28(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_29(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_30(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_31(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_32(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h6/* 6*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_33(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h7/* 7*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_34(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'h8/* 8*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_35(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [25:0] io_configs_en,
    input [275:0] io_ipin_in,
    input [572:0] io_chanxy_in,
    output[104:0] io_chanxy_out,
    output[7:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[263:0] T0;
  wire[831:0] this_config_io_configs_out;
  wire[91:0] T1;
  wire[199:0] T2;
  wire[30:0] T3;
  wire[22:0] this_sbcb_io_ipin_out;
  wire[7:0] this_clb_io_clb_out;
  wire[7:0] T4;
  wire[255:0] T5;
  wire[39:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[104:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[10'h333/* 819*/:10'h22c/* 556*/];
  assign T1 = this_config_io_configs_out[10'h22b/* 555*/:9'h1d0/* 464*/];
  assign T2 = this_config_io_configs_out[9'h1cf/* 463*/:9'h108/* 264*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[9'h107/* 263*/:9'h100/* 256*/];
  assign T5 = this_config_io_configs_out[8'hff/* 255*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {4'h0/* 0*/, 4'ha/* 10*/};
  assign io_x_loc = T7;
  assign T7 = {4'h0/* 0*/, 4'h9/* 9*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_26 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_13 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


