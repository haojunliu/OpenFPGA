module fpga(
    input [39:0] top_in,
    input [39:0] bot_in,
    input [39:0] left_in,
    input [39:0] right_in,
    output [39:0] top_out,
    output [39:0] bot_out,
    output [39:0] left_out,
    output [39:0] right_out,
    input [223:0] configs_in,
    input [244:0] configs_en,
    input ff_en, clock, rst
);

    // Interconnection Wire Declaration
    wire wire_25;
    wire wire_28;
    wire wire_31;
    wire wire_34;
    wire wire_37;
    wire wire_40;
    wire wire_43;
    wire wire_46;
    wire wire_73;
    wire wire_76;
    wire wire_79;
    wire wire_82;
    wire wire_85;
    wire wire_88;
    wire wire_91;
    wire wire_94;
    wire wire_121;
    wire wire_124;
    wire wire_127;
    wire wire_130;
    wire wire_133;
    wire wire_136;
    wire wire_139;
    wire wire_142;
    wire wire_169;
    wire wire_172;
    wire wire_175;
    wire wire_178;
    wire wire_181;
    wire wire_184;
    wire wire_187;
    wire wire_190;
    wire wire_217;
    wire wire_220;
    wire wire_223;
    wire wire_226;
    wire wire_229;
    wire wire_232;
    wire wire_235;
    wire wire_238;
    wire wire_265;
    wire wire_268;
    wire wire_271;
    wire wire_274;
    wire wire_277;
    wire wire_280;
    wire wire_283;
    wire wire_286;
    wire wire_333;
    wire wire_334;
    wire wire_335;
    wire wire_336;
    wire wire_337;
    wire wire_338;
    wire wire_339;
    wire wire_340;
    wire wire_341;
    wire wire_342;
    wire wire_389;
    wire wire_390;
    wire wire_391;
    wire wire_392;
    wire wire_393;
    wire wire_394;
    wire wire_395;
    wire wire_396;
    wire wire_397;
    wire wire_398;
    wire wire_445;
    wire wire_446;
    wire wire_447;
    wire wire_448;
    wire wire_449;
    wire wire_450;
    wire wire_451;
    wire wire_452;
    wire wire_453;
    wire wire_454;
    wire wire_501;
    wire wire_502;
    wire wire_503;
    wire wire_504;
    wire wire_505;
    wire wire_506;
    wire wire_507;
    wire wire_508;
    wire wire_509;
    wire wire_510;
    wire wire_557;
    wire wire_558;
    wire wire_559;
    wire wire_560;
    wire wire_561;
    wire wire_562;
    wire wire_563;
    wire wire_564;
    wire wire_565;
    wire wire_566;
    wire wire_593;
    wire wire_596;
    wire wire_599;
    wire wire_602;
    wire wire_605;
    wire wire_608;
    wire wire_611;
    wire wire_614;
    wire wire_641;
    wire wire_644;
    wire wire_647;
    wire wire_650;
    wire wire_653;
    wire wire_656;
    wire wire_659;
    wire wire_662;
    wire wire_709;
    wire wire_710;
    wire wire_711;
    wire wire_712;
    wire wire_713;
    wire wire_714;
    wire wire_715;
    wire wire_716;
    wire wire_717;
    wire wire_718;
    wire wire_765;
    wire wire_766;
    wire wire_767;
    wire wire_768;
    wire wire_769;
    wire wire_770;
    wire wire_771;
    wire wire_772;
    wire wire_773;
    wire wire_774;
    wire wire_821;
    wire wire_822;
    wire wire_823;
    wire wire_824;
    wire wire_825;
    wire wire_826;
    wire wire_827;
    wire wire_828;
    wire wire_829;
    wire wire_830;
    wire wire_877;
    wire wire_878;
    wire wire_879;
    wire wire_880;
    wire wire_881;
    wire wire_882;
    wire wire_883;
    wire wire_884;
    wire wire_885;
    wire wire_886;
    wire wire_933;
    wire wire_934;
    wire wire_935;
    wire wire_936;
    wire wire_937;
    wire wire_938;
    wire wire_939;
    wire wire_940;
    wire wire_941;
    wire wire_942;
    wire wire_969;
    wire wire_972;
    wire wire_975;
    wire wire_978;
    wire wire_981;
    wire wire_984;
    wire wire_987;
    wire wire_990;
    wire wire_1017;
    wire wire_1020;
    wire wire_1023;
    wire wire_1026;
    wire wire_1029;
    wire wire_1032;
    wire wire_1035;
    wire wire_1038;
    wire wire_1085;
    wire wire_1086;
    wire wire_1087;
    wire wire_1088;
    wire wire_1089;
    wire wire_1090;
    wire wire_1091;
    wire wire_1092;
    wire wire_1093;
    wire wire_1094;
    wire wire_1141;
    wire wire_1142;
    wire wire_1143;
    wire wire_1144;
    wire wire_1145;
    wire wire_1146;
    wire wire_1147;
    wire wire_1148;
    wire wire_1149;
    wire wire_1150;
    wire wire_1197;
    wire wire_1198;
    wire wire_1199;
    wire wire_1200;
    wire wire_1201;
    wire wire_1202;
    wire wire_1203;
    wire wire_1204;
    wire wire_1205;
    wire wire_1206;
    wire wire_1253;
    wire wire_1254;
    wire wire_1255;
    wire wire_1256;
    wire wire_1257;
    wire wire_1258;
    wire wire_1259;
    wire wire_1260;
    wire wire_1261;
    wire wire_1262;
    wire wire_1309;
    wire wire_1310;
    wire wire_1311;
    wire wire_1312;
    wire wire_1313;
    wire wire_1314;
    wire wire_1315;
    wire wire_1316;
    wire wire_1317;
    wire wire_1318;
    wire wire_1345;
    wire wire_1348;
    wire wire_1351;
    wire wire_1354;
    wire wire_1357;
    wire wire_1360;
    wire wire_1363;
    wire wire_1366;
    wire wire_1393;
    wire wire_1396;
    wire wire_1399;
    wire wire_1402;
    wire wire_1405;
    wire wire_1408;
    wire wire_1411;
    wire wire_1414;
    wire wire_1461;
    wire wire_1462;
    wire wire_1463;
    wire wire_1464;
    wire wire_1465;
    wire wire_1466;
    wire wire_1467;
    wire wire_1468;
    wire wire_1469;
    wire wire_1470;
    wire wire_1517;
    wire wire_1518;
    wire wire_1519;
    wire wire_1520;
    wire wire_1521;
    wire wire_1522;
    wire wire_1523;
    wire wire_1524;
    wire wire_1525;
    wire wire_1526;
    wire wire_1573;
    wire wire_1574;
    wire wire_1575;
    wire wire_1576;
    wire wire_1577;
    wire wire_1578;
    wire wire_1579;
    wire wire_1580;
    wire wire_1581;
    wire wire_1582;
    wire wire_1629;
    wire wire_1630;
    wire wire_1631;
    wire wire_1632;
    wire wire_1633;
    wire wire_1634;
    wire wire_1635;
    wire wire_1636;
    wire wire_1637;
    wire wire_1638;
    wire wire_1685;
    wire wire_1686;
    wire wire_1687;
    wire wire_1688;
    wire wire_1689;
    wire wire_1690;
    wire wire_1691;
    wire wire_1692;
    wire wire_1693;
    wire wire_1694;
    wire wire_1721;
    wire wire_1724;
    wire wire_1727;
    wire wire_1730;
    wire wire_1733;
    wire wire_1736;
    wire wire_1739;
    wire wire_1742;
    wire wire_1769;
    wire wire_1772;
    wire wire_1775;
    wire wire_1778;
    wire wire_1781;
    wire wire_1784;
    wire wire_1787;
    wire wire_1790;
    wire wire_1837;
    wire wire_1838;
    wire wire_1839;
    wire wire_1840;
    wire wire_1841;
    wire wire_1842;
    wire wire_1843;
    wire wire_1844;
    wire wire_1845;
    wire wire_1846;
    wire wire_1893;
    wire wire_1894;
    wire wire_1895;
    wire wire_1896;
    wire wire_1897;
    wire wire_1898;
    wire wire_1899;
    wire wire_1900;
    wire wire_1901;
    wire wire_1902;
    wire wire_1949;
    wire wire_1950;
    wire wire_1951;
    wire wire_1952;
    wire wire_1953;
    wire wire_1954;
    wire wire_1955;
    wire wire_1956;
    wire wire_1957;
    wire wire_1958;
    wire wire_2005;
    wire wire_2006;
    wire wire_2007;
    wire wire_2008;
    wire wire_2009;
    wire wire_2010;
    wire wire_2011;
    wire wire_2012;
    wire wire_2013;
    wire wire_2014;
    wire wire_2061;
    wire wire_2062;
    wire wire_2063;
    wire wire_2064;
    wire wire_2065;
    wire wire_2066;
    wire wire_2067;
    wire wire_2068;
    wire wire_2069;
    wire wire_2070;
    wire wire_2097;
    wire wire_2100;
    wire wire_2103;
    wire wire_2106;
    wire wire_2109;
    wire wire_2112;
    wire wire_2115;
    wire wire_2118;
    wire wire_2145;
    wire wire_2148;
    wire wire_2151;
    wire wire_2154;
    wire wire_2157;
    wire wire_2160;
    wire wire_2163;
    wire wire_2166;
    wire wire_2193;
    wire wire_2196;
    wire wire_2199;
    wire wire_2202;
    wire wire_2205;
    wire wire_2208;
    wire wire_2211;
    wire wire_2214;
    wire wire_2241;
    wire wire_2244;
    wire wire_2247;
    wire wire_2250;
    wire wire_2253;
    wire wire_2256;
    wire wire_2259;
    wire wire_2262;
    wire wire_2289;
    wire wire_2292;
    wire wire_2295;
    wire wire_2298;
    wire wire_2301;
    wire wire_2304;
    wire wire_2307;
    wire wire_2310;
    wire wire_2337;
    wire wire_2340;
    wire wire_2343;
    wire wire_2346;
    wire wire_2349;
    wire wire_2352;
    wire wire_2355;
    wire wire_2358;
    wire wire_2360;
    wire wire_2361;
    wire wire_2362;
    wire wire_2363;
    wire wire_2364;
    wire wire_2365;
    wire wire_2366;
    wire wire_2367;
    wire wire_2368;
    wire wire_2369;
    wire wire_2370;
    wire wire_2371;
    wire wire_2372;
    wire wire_2373;
    wire wire_2374;
    wire wire_2375;
    wire wire_2376;
    wire wire_2377;
    wire wire_2378;
    wire wire_2379;
    wire wire_2380;
    wire wire_2381;
    wire wire_2382;
    wire wire_2383;
    wire wire_2384;
    wire wire_2385;
    wire wire_2386;
    wire wire_2387;
    wire wire_2388;
    wire wire_2389;
    wire wire_2390;
    wire wire_2391;
    wire wire_2392;
    wire wire_2393;
    wire wire_2394;
    wire wire_2395;
    wire wire_2396;
    wire wire_2397;
    wire wire_2398;
    wire wire_2399;
    wire wire_2400;
    wire wire_2401;
    wire wire_2402;
    wire wire_2403;
    wire wire_2404;
    wire wire_2405;
    wire wire_2406;
    wire wire_2407;
    wire wire_2408;
    wire wire_2409;
    wire wire_2410;
    wire wire_2411;
    wire wire_2412;
    wire wire_2413;
    wire wire_2414;
    wire wire_2415;
    wire wire_2416;
    wire wire_2417;
    wire wire_2418;
    wire wire_2419;
    wire wire_2420;
    wire wire_2421;
    wire wire_2422;
    wire wire_2423;
    wire wire_2424;
    wire wire_2425;
    wire wire_2426;
    wire wire_2427;
    wire wire_2428;
    wire wire_2429;
    wire wire_2430;
    wire wire_2431;
    wire wire_2432;
    wire wire_2433;
    wire wire_2434;
    wire wire_2435;
    wire wire_2436;
    wire wire_2437;
    wire wire_2438;
    wire wire_2439;
    wire wire_2440;
    wire wire_2441;
    wire wire_2442;
    wire wire_2443;
    wire wire_2444;
    wire wire_2445;
    wire wire_2446;
    wire wire_2447;
    wire wire_2448;
    wire wire_2449;
    wire wire_2450;
    wire wire_2451;
    wire wire_2452;
    wire wire_2453;
    wire wire_2454;
    wire wire_2455;
    wire wire_2456;
    wire wire_2457;
    wire wire_2458;
    wire wire_2459;
    wire wire_2460;
    wire wire_2461;
    wire wire_2462;
    wire wire_2463;
    wire wire_2464;
    wire wire_2465;
    wire wire_2466;
    wire wire_2467;
    wire wire_2468;
    wire wire_2469;
    wire wire_2470;
    wire wire_2471;
    wire wire_2472;
    wire wire_2473;
    wire wire_2474;
    wire wire_2475;
    wire wire_2476;
    wire wire_2477;
    wire wire_2478;
    wire wire_2479;
    wire wire_2480;
    wire wire_2481;
    wire wire_2482;
    wire wire_2483;
    wire wire_2484;
    wire wire_2485;
    wire wire_2486;
    wire wire_2487;
    wire wire_2488;
    wire wire_2489;
    wire wire_2490;
    wire wire_2491;
    wire wire_2492;
    wire wire_2493;
    wire wire_2494;
    wire wire_2495;
    wire wire_2496;
    wire wire_2497;
    wire wire_2498;
    wire wire_2499;
    wire wire_2500;
    wire wire_2501;
    wire wire_2502;
    wire wire_2503;
    wire wire_2504;
    wire wire_2505;
    wire wire_2506;
    wire wire_2507;
    wire wire_2508;
    wire wire_2509;
    wire wire_2510;
    wire wire_2511;
    wire wire_2512;
    wire wire_2513;
    wire wire_2514;
    wire wire_2515;
    wire wire_2516;
    wire wire_2517;
    wire wire_2518;
    wire wire_2519;
    wire wire_2520;
    wire wire_2521;
    wire wire_2522;
    wire wire_2523;
    wire wire_2524;
    wire wire_2525;
    wire wire_2526;
    wire wire_2527;
    wire wire_2528;
    wire wire_2529;
    wire wire_2530;
    wire wire_2531;
    wire wire_2532;
    wire wire_2533;
    wire wire_2534;
    wire wire_2535;
    wire wire_2536;
    wire wire_2537;
    wire wire_2538;
    wire wire_2539;
    wire wire_2540;
    wire wire_2541;
    wire wire_2542;
    wire wire_2543;
    wire wire_2544;
    wire wire_2545;
    wire wire_2546;
    wire wire_2547;
    wire wire_2548;
    wire wire_2549;
    wire wire_2550;
    wire wire_2551;
    wire wire_2552;
    wire wire_2553;
    wire wire_2554;
    wire wire_2555;
    wire wire_2556;
    wire wire_2557;
    wire wire_2558;
    wire wire_2559;
    wire wire_2560;
    wire wire_2561;
    wire wire_2562;
    wire wire_2563;
    wire wire_2564;
    wire wire_2565;
    wire wire_2566;
    wire wire_2567;
    wire wire_2568;
    wire wire_2569;
    wire wire_2570;
    wire wire_2571;
    wire wire_2572;
    wire wire_2573;
    wire wire_2574;
    wire wire_2575;
    wire wire_2576;
    wire wire_2577;
    wire wire_2578;
    wire wire_2579;
    wire wire_2580;
    wire wire_2581;
    wire wire_2582;
    wire wire_2583;
    wire wire_2584;
    wire wire_2585;
    wire wire_2586;
    wire wire_2587;
    wire wire_2588;
    wire wire_2589;
    wire wire_2590;
    wire wire_2591;
    wire wire_2592;
    wire wire_2593;
    wire wire_2594;
    wire wire_2595;
    wire wire_2596;
    wire wire_2597;
    wire wire_2598;
    wire wire_2599;
    wire wire_2600;
    wire wire_2601;
    wire wire_2602;
    wire wire_2603;
    wire wire_2604;
    wire wire_2605;
    wire wire_2606;
    wire wire_2607;
    wire wire_2608;
    wire wire_2609;
    wire wire_2610;
    wire wire_2611;
    wire wire_2612;
    wire wire_2613;
    wire wire_2614;
    wire wire_2615;
    wire wire_2616;
    wire wire_2617;
    wire wire_2618;
    wire wire_2619;
    wire wire_2620;
    wire wire_2621;
    wire wire_2622;
    wire wire_2623;
    wire wire_2624;
    wire wire_2625;
    wire wire_2626;
    wire wire_2627;
    wire wire_2628;
    wire wire_2629;
    wire wire_2630;
    wire wire_2631;
    wire wire_2632;
    wire wire_2633;
    wire wire_2634;
    wire wire_2635;
    wire wire_2636;
    wire wire_2637;
    wire wire_2638;
    wire wire_2639;
    wire wire_2640;
    wire wire_2641;
    wire wire_2642;
    wire wire_2643;
    wire wire_2644;
    wire wire_2645;
    wire wire_2646;
    wire wire_2647;
    wire wire_2648;
    wire wire_2649;
    wire wire_2650;
    wire wire_2651;
    wire wire_2652;
    wire wire_2653;
    wire wire_2654;
    wire wire_2655;
    wire wire_2656;
    wire wire_2657;
    wire wire_2658;
    wire wire_2659;
    wire wire_2660;
    wire wire_2661;
    wire wire_2662;
    wire wire_2663;
    wire wire_2664;
    wire wire_2665;
    wire wire_2666;
    wire wire_2667;
    wire wire_2668;
    wire wire_2669;
    wire wire_2670;
    wire wire_2671;
    wire wire_2672;
    wire wire_2673;
    wire wire_2674;
    wire wire_2675;
    wire wire_2676;
    wire wire_2677;
    wire wire_2678;
    wire wire_2679;
    wire wire_2680;
    wire wire_2681;
    wire wire_2682;
    wire wire_2683;
    wire wire_2684;
    wire wire_2685;
    wire wire_2686;
    wire wire_2687;
    wire wire_2688;
    wire wire_2689;
    wire wire_2690;
    wire wire_2691;
    wire wire_2692;
    wire wire_2693;
    wire wire_2694;
    wire wire_2695;
    wire wire_2696;
    wire wire_2697;
    wire wire_2698;
    wire wire_2699;
    wire wire_2700;
    wire wire_2701;
    wire wire_2702;
    wire wire_2703;
    wire wire_2704;
    wire wire_2705;
    wire wire_2706;
    wire wire_2707;
    wire wire_2708;
    wire wire_2709;
    wire wire_2710;
    wire wire_2711;
    wire wire_2712;
    wire wire_2713;
    wire wire_2714;
    wire wire_2715;
    wire wire_2716;
    wire wire_2717;
    wire wire_2718;
    wire wire_2719;
    wire wire_2720;
    wire wire_2721;
    wire wire_2722;
    wire wire_2723;
    wire wire_2724;
    wire wire_2725;
    wire wire_2726;
    wire wire_2727;
    wire wire_2728;
    wire wire_2729;
    wire wire_2730;
    wire wire_2731;
    wire wire_2732;
    wire wire_2733;
    wire wire_2734;
    wire wire_2735;
    wire wire_2736;
    wire wire_2737;
    wire wire_2738;
    wire wire_2739;
    wire wire_2740;
    wire wire_2741;
    wire wire_2742;
    wire wire_2743;
    wire wire_2744;
    wire wire_2745;
    wire wire_2746;
    wire wire_2747;
    wire wire_2748;
    wire wire_2749;
    wire wire_2750;
    wire wire_2751;
    wire wire_2752;
    wire wire_2753;
    wire wire_2754;
    wire wire_2755;
    wire wire_2756;
    wire wire_2757;
    wire wire_2758;
    wire wire_2759;
    wire wire_2760;
    wire wire_2761;
    wire wire_2762;
    wire wire_2763;
    wire wire_2764;
    wire wire_2765;
    wire wire_2766;
    wire wire_2767;
    wire wire_2768;
    wire wire_2769;
    wire wire_2770;
    wire wire_2771;
    wire wire_2772;
    wire wire_2773;
    wire wire_2774;
    wire wire_2775;
    wire wire_2776;
    wire wire_2777;
    wire wire_2778;
    wire wire_2779;
    wire wire_2780;
    wire wire_2781;
    wire wire_2782;
    wire wire_2783;
    wire wire_2784;
    wire wire_2785;
    wire wire_2786;
    wire wire_2787;
    wire wire_2788;
    wire wire_2789;
    wire wire_2790;
    wire wire_2791;
    wire wire_2792;
    wire wire_2793;
    wire wire_2794;
    wire wire_2795;
    wire wire_2796;
    wire wire_2797;
    wire wire_2798;
    wire wire_2799;
    wire wire_2800;
    wire wire_2801;
    wire wire_2802;
    wire wire_2803;
    wire wire_2804;
    wire wire_2805;
    wire wire_2806;
    wire wire_2807;
    wire wire_2808;
    wire wire_2809;
    wire wire_2810;
    wire wire_2811;
    wire wire_2812;
    wire wire_2813;
    wire wire_2814;
    wire wire_2815;
    wire wire_2816;
    wire wire_2817;
    wire wire_2818;
    wire wire_2819;
    wire wire_2820;
    wire wire_2821;
    wire wire_2822;
    wire wire_2823;
    wire wire_2824;
    wire wire_2825;
    wire wire_2826;
    wire wire_2827;
    wire wire_2828;
    wire wire_2829;
    wire wire_2830;
    wire wire_2831;
    wire wire_2832;
    wire wire_2833;
    wire wire_2834;
    wire wire_2835;
    wire wire_2836;
    wire wire_2837;
    wire wire_2838;
    wire wire_2839;
    wire wire_2840;
    wire wire_2841;
    wire wire_2842;
    wire wire_2843;
    wire wire_2844;
    wire wire_2845;
    wire wire_2846;
    wire wire_2847;
    wire wire_2848;
    wire wire_2849;
    wire wire_2850;
    wire wire_2851;
    wire wire_2852;
    wire wire_2853;
    wire wire_2854;
    wire wire_2855;
    wire wire_2856;
    wire wire_2857;
    wire wire_2858;
    wire wire_2859;
    wire wire_2860;
    wire wire_2861;
    wire wire_2862;
    wire wire_2863;
    wire wire_2864;
    wire wire_2865;
    wire wire_2866;
    wire wire_2867;
    wire wire_2868;
    wire wire_2869;
    wire wire_2870;
    wire wire_2871;
    wire wire_2872;
    wire wire_2873;
    wire wire_2874;
    wire wire_2875;
    wire wire_2876;
    wire wire_2877;
    wire wire_2878;
    wire wire_2879;
    wire wire_2880;
    wire wire_2881;
    wire wire_2882;
    wire wire_2883;
    wire wire_2884;
    wire wire_2885;
    wire wire_2886;
    wire wire_2887;
    wire wire_2888;
    wire wire_2889;
    wire wire_2890;
    wire wire_2891;
    wire wire_2892;
    wire wire_2893;
    wire wire_2894;
    wire wire_2895;
    wire wire_2896;
    wire wire_2897;
    wire wire_2898;
    wire wire_2899;
    wire wire_2900;
    wire wire_2901;
    wire wire_2902;
    wire wire_2903;
    wire wire_2904;
    wire wire_2905;
    wire wire_2906;
    wire wire_2907;
    wire wire_2908;
    wire wire_2909;
    wire wire_2910;
    wire wire_2911;
    wire wire_2912;
    wire wire_2913;
    wire wire_2914;
    wire wire_2915;
    wire wire_2916;
    wire wire_2917;
    wire wire_2918;
    wire wire_2919;
    wire wire_2920;
    wire wire_2921;
    wire wire_2922;
    wire wire_2923;
    wire wire_2924;
    wire wire_2925;
    wire wire_2926;
    wire wire_2927;
    wire wire_2928;
    wire wire_2929;
    wire wire_2930;
    wire wire_2931;
    wire wire_2932;
    wire wire_2933;
    wire wire_2934;
    wire wire_2935;
    wire wire_2936;
    wire wire_2937;
    wire wire_2938;
    wire wire_2939;
    wire wire_2940;
    wire wire_2941;
    wire wire_2942;
    wire wire_2943;
    wire wire_2944;
    wire wire_2945;
    wire wire_2946;
    wire wire_2947;
    wire wire_2948;
    wire wire_2949;
    wire wire_2950;
    wire wire_2951;
    wire wire_2952;
    wire wire_2953;
    wire wire_2954;
    wire wire_2955;
    wire wire_2956;
    wire wire_2957;
    wire wire_2958;
    wire wire_2959;
    wire wire_2960;
    wire wire_2961;
    wire wire_2962;
    wire wire_2963;
    wire wire_2964;
    wire wire_2965;
    wire wire_2966;
    wire wire_2967;
    wire wire_2968;
    wire wire_2969;
    wire wire_2970;
    wire wire_2971;
    wire wire_2972;
    wire wire_2973;
    wire wire_2974;
    wire wire_2975;
    wire wire_2976;
    wire wire_2977;
    wire wire_2978;
    wire wire_2979;
    wire wire_2980;
    wire wire_2981;
    wire wire_2982;
    wire wire_2983;
    wire wire_2984;
    wire wire_2985;
    wire wire_2986;
    wire wire_2987;
    wire wire_2988;
    wire wire_2989;
    wire wire_2990;
    wire wire_2991;
    wire wire_2992;
    wire wire_2993;
    wire wire_2994;
    wire wire_2995;
    wire wire_2996;
    wire wire_2997;
    wire wire_2998;
    wire wire_2999;
    wire wire_3000;
    wire wire_3001;
    wire wire_3002;
    wire wire_3003;
    wire wire_3004;
    wire wire_3005;
    wire wire_3006;
    wire wire_3007;
    wire wire_3008;
    wire wire_3009;
    wire wire_3010;
    wire wire_3011;
    wire wire_3012;
    wire wire_3013;
    wire wire_3014;
    wire wire_3015;
    wire wire_3016;
    wire wire_3017;
    wire wire_3018;
    wire wire_3019;
    wire wire_3020;
    wire wire_3021;
    wire wire_3022;
    wire wire_3023;
    wire wire_3024;
    wire wire_3025;
    wire wire_3026;
    wire wire_3027;
    wire wire_3028;
    wire wire_3029;
    wire wire_3030;
    wire wire_3031;
    wire wire_3032;
    wire wire_3033;
    wire wire_3034;
    wire wire_3035;
    wire wire_3036;
    wire wire_3037;
    wire wire_3038;
    wire wire_3039;
    wire wire_3040;
    wire wire_3041;
    wire wire_3042;
    wire wire_3043;
    wire wire_3044;
    wire wire_3045;
    wire wire_3046;
    wire wire_3047;
    wire wire_3048;
    wire wire_3049;
    wire wire_3050;
    wire wire_3051;
    wire wire_3052;
    wire wire_3053;
    wire wire_3054;
    wire wire_3055;
    wire wire_3056;
    wire wire_3057;
    wire wire_3058;
    wire wire_3059;
    wire wire_3060;
    wire wire_3061;
    wire wire_3062;
    wire wire_3063;
    wire wire_3064;
    wire wire_3065;
    wire wire_3066;
    wire wire_3067;
    wire wire_3068;
    wire wire_3069;
    wire wire_3070;
    wire wire_3071;
    wire wire_3072;
    wire wire_3073;
    wire wire_3074;
    wire wire_3075;
    wire wire_3076;
    wire wire_3077;
    wire wire_3078;
    wire wire_3079;
    wire wire_3080;
    wire wire_3081;
    wire wire_3082;
    wire wire_3083;
    wire wire_3084;
    wire wire_3085;
    wire wire_3086;
    wire wire_3087;
    wire wire_3088;
    wire wire_3089;
    wire wire_3090;
    wire wire_3091;
    wire wire_3092;
    wire wire_3093;
    wire wire_3094;
    wire wire_3095;
    wire wire_3096;
    wire wire_3097;
    wire wire_3098;
    wire wire_3099;
    wire wire_3100;
    wire wire_3101;
    wire wire_3102;
    wire wire_3103;
    wire wire_3104;
    wire wire_3105;
    wire wire_3106;
    wire wire_3107;
    wire wire_3108;
    wire wire_3109;
    wire wire_3110;
    wire wire_3111;
    wire wire_3112;
    wire wire_3113;
    wire wire_3114;
    wire wire_3115;
    wire wire_3116;
    wire wire_3117;
    wire wire_3118;
    wire wire_3119;
    wire wire_3120;
    wire wire_3121;
    wire wire_3122;
    wire wire_3123;
    wire wire_3124;
    wire wire_3125;
    wire wire_3126;
    wire wire_3127;
    wire wire_3128;
    wire wire_3129;
    wire wire_3130;
    wire wire_3131;
    wire wire_3132;
    wire wire_3133;
    wire wire_3134;
    wire wire_3135;
    wire wire_3136;
    wire wire_3137;
    wire wire_3138;
    wire wire_3139;
    wire wire_3140;
    wire wire_3141;
    wire wire_3142;
    wire wire_3143;
    wire wire_3144;
    wire wire_3145;
    wire wire_3146;
    wire wire_3147;
    wire wire_3148;
    wire wire_3149;
    wire wire_3150;
    wire wire_3151;
    wire wire_3152;
    wire wire_3153;
    wire wire_3154;
    wire wire_3155;
    wire wire_3156;
    wire wire_3157;
    wire wire_3158;
    wire wire_3159;
    wire wire_3160;
    wire wire_3161;
    wire wire_3162;
    wire wire_3163;
    wire wire_3164;
    wire wire_3165;
    wire wire_3166;
    wire wire_3167;
    wire wire_3168;
    wire wire_3169;
    wire wire_3170;
    wire wire_3171;
    wire wire_3172;
    wire wire_3173;
    wire wire_3174;
    wire wire_3175;
    wire wire_3176;
    wire wire_3177;
    wire wire_3178;
    wire wire_3179;
    wire wire_3180;
    wire wire_3181;
    wire wire_3182;
    wire wire_3183;
    wire wire_3184;
    wire wire_3185;
    wire wire_3186;
    wire wire_3187;
    wire wire_3188;
    wire wire_3189;
    wire wire_3190;
    wire wire_3191;
    wire wire_3192;
    wire wire_3193;
    wire wire_3194;
    wire wire_3195;
    wire wire_3196;
    wire wire_3197;
    wire wire_3198;
    wire wire_3199;
    wire wire_3200;
    wire wire_3201;
    wire wire_3202;
    wire wire_3203;
    wire wire_3204;
    wire wire_3205;
    wire wire_3206;
    wire wire_3207;
    wire wire_3208;
    wire wire_3209;
    wire wire_3210;
    wire wire_3211;
    wire wire_3212;
    wire wire_3213;
    wire wire_3214;
    wire wire_3215;
    wire wire_3216;
    wire wire_3217;
    wire wire_3218;
    wire wire_3219;
    wire wire_3220;
    wire wire_3221;
    wire wire_3222;
    wire wire_3223;
    wire wire_3224;
    wire wire_3225;
    wire wire_3226;
    wire wire_3227;
    wire wire_3228;
    wire wire_3229;
    wire wire_3230;
    wire wire_3231;
    wire wire_3232;
    wire wire_3233;
    wire wire_3234;
    wire wire_3235;
    wire wire_3236;
    wire wire_3237;
    wire wire_3238;
    wire wire_3239;
    wire wire_3240;
    wire wire_3241;
    wire wire_3242;
    wire wire_3243;
    wire wire_3244;
    wire wire_3245;
    wire wire_3246;
    wire wire_3247;
    wire wire_3248;
    wire wire_3249;
    wire wire_3250;
    wire wire_3251;
    wire wire_3252;
    wire wire_3253;
    wire wire_3254;
    wire wire_3255;
    wire wire_3256;
    wire wire_3257;
    wire wire_3258;
    wire wire_3259;
    wire wire_3260;
    wire wire_3261;
    wire wire_3262;
    wire wire_3263;
    wire wire_3264;
    wire wire_3265;
    wire wire_3266;
    wire wire_3267;
    wire wire_3268;
    wire wire_3269;
    wire wire_3270;
    wire wire_3271;
    wire wire_3272;
    wire wire_3273;
    wire wire_3274;
    wire wire_3275;
    wire wire_3276;
    wire wire_3277;
    wire wire_3278;
    wire wire_3279;
    wire wire_3280;
    wire wire_3281;
    wire wire_3282;
    wire wire_3283;
    wire wire_3284;
    wire wire_3285;
    wire wire_3286;
    wire wire_3287;
    wire wire_3288;
    wire wire_3289;
    wire wire_3290;
    wire wire_3291;
    wire wire_3292;
    wire wire_3293;
    wire wire_3294;
    wire wire_3295;
    wire wire_3296;
    wire wire_3297;
    wire wire_3298;
    wire wire_3299;
    wire wire_3300;
    wire wire_3301;
    wire wire_3302;
    wire wire_3303;
    wire wire_3304;
    wire wire_3305;
    wire wire_3306;
    wire wire_3307;
    wire wire_3308;
    wire wire_3309;
    wire wire_3310;
    wire wire_3311;
    wire wire_3312;
    wire wire_3313;
    wire wire_3314;
    wire wire_3315;
    wire wire_3316;
    wire wire_3317;
    wire wire_3318;
    wire wire_3319;
    wire wire_3320;
    wire wire_3321;
    wire wire_3322;
    wire wire_3323;
    wire wire_3324;
    wire wire_3325;
    wire wire_3326;
    wire wire_3327;
    wire wire_3328;
    wire wire_3329;
    wire wire_3330;
    wire wire_3331;
    wire wire_3332;
    wire wire_3333;
    wire wire_3334;
    wire wire_3335;
    wire wire_3336;
    wire wire_3337;
    wire wire_3338;
    wire wire_3339;
    wire wire_3340;
    wire wire_3341;
    wire wire_3342;
    wire wire_3343;
    wire wire_3344;
    wire wire_3345;
    wire wire_3346;
    wire wire_3347;
    wire wire_3348;
    wire wire_3349;
    wire wire_3350;
    wire wire_3351;
    wire wire_3352;
    wire wire_3353;
    wire wire_3354;
    wire wire_3355;
    wire wire_3356;
    wire wire_3357;
    wire wire_3358;
    wire wire_3359;
    wire wire_3360;
    wire wire_3361;
    wire wire_3362;
    wire wire_3363;
    wire wire_3364;
    wire wire_3365;
    wire wire_3366;
    wire wire_3367;
    wire wire_3368;
    wire wire_3369;
    wire wire_3370;
    wire wire_3371;
    wire wire_3372;
    wire wire_3373;
    wire wire_3374;
    wire wire_3375;
    wire wire_3376;
    wire wire_3377;
    wire wire_3378;
    wire wire_3379;
    wire wire_3380;
    wire wire_3381;
    wire wire_3382;
    wire wire_3383;
    wire wire_3384;
    wire wire_3385;
    wire wire_3386;
    wire wire_3387;
    wire wire_3388;
    wire wire_3389;
    wire wire_3390;
    wire wire_3391;
    wire wire_3392;
    wire wire_3393;
    wire wire_3394;
    wire wire_3395;
    wire wire_3396;
    wire wire_3397;
    wire wire_3398;
    wire wire_3399;
    wire wire_3400;
    wire wire_3401;
    wire wire_3402;
    wire wire_3403;
    wire wire_3404;
    wire wire_3405;
    wire wire_3406;
    wire wire_3407;
    wire wire_3408;
    wire wire_3409;
    wire wire_3410;
    wire wire_3411;
    wire wire_3412;
    wire wire_3413;
    wire wire_3414;
    wire wire_3415;
    wire wire_3416;
    wire wire_3417;
    wire wire_3418;
    wire wire_3419;
    wire wire_3420;
    wire wire_3421;
    wire wire_3422;
    wire wire_3423;
    wire wire_3424;
    wire wire_3425;
    wire wire_3426;
    wire wire_3427;
    wire wire_3428;
    wire wire_3429;
    wire wire_3430;
    wire wire_3431;
    wire wire_3432;
    wire wire_3433;
    wire wire_3434;
    wire wire_3435;
    wire wire_3436;
    wire wire_3437;
    wire wire_3438;
    wire wire_3439;
    wire wire_3440;
    wire wire_3441;
    wire wire_3442;
    wire wire_3443;
    wire wire_3444;
    wire wire_3445;
    wire wire_3446;
    wire wire_3447;
    wire wire_3448;
    wire wire_3449;
    wire wire_3450;
    wire wire_3451;
    wire wire_3452;
    wire wire_3453;
    wire wire_3454;
    wire wire_3455;
    wire wire_3456;
    wire wire_3457;
    wire wire_3458;
    wire wire_3459;
    wire wire_3460;
    wire wire_3461;
    wire wire_3462;
    wire wire_3463;
    wire wire_3464;
    wire wire_3465;
    wire wire_3466;
    wire wire_3467;
    wire wire_3468;
    wire wire_3469;
    wire wire_3470;
    wire wire_3471;
    wire wire_3472;
    wire wire_3473;
    wire wire_3474;
    wire wire_3475;
    wire wire_3476;
    wire wire_3477;
    wire wire_3478;
    wire wire_3479;
    wire wire_3480;
    wire wire_3481;
    wire wire_3482;
    wire wire_3483;
    wire wire_3484;
    wire wire_3485;
    wire wire_3486;
    wire wire_3487;
    wire wire_3488;
    wire wire_3489;
    wire wire_3490;
    wire wire_3491;
    wire wire_3492;
    wire wire_3493;
    wire wire_3494;
    wire wire_3495;
    wire wire_3496;
    wire wire_3497;
    wire wire_3498;
    wire wire_3499;
    wire wire_3500;
    wire wire_3501;
    wire wire_3502;
    wire wire_3503;
    wire wire_3504;
    wire wire_3505;
    wire wire_3506;
    wire wire_3507;
    wire wire_3508;
    wire wire_3509;
    wire wire_3510;
    wire wire_3511;
    wire wire_3512;
    wire wire_3513;
    wire wire_3514;
    wire wire_3515;
    wire wire_3516;
    wire wire_3517;
    wire wire_3518;
    wire wire_3519;
    wire wire_3520;
    wire wire_3521;
    wire wire_3522;
    wire wire_3523;
    wire wire_3524;
    wire wire_3525;
    wire wire_3526;
    wire wire_3527;
    wire wire_3528;
    wire wire_3529;
    wire wire_3530;
    wire wire_3531;
    wire wire_3532;
    wire wire_3533;
    wire wire_3534;
    wire wire_3535;
    wire wire_3536;
    wire wire_3537;
    wire wire_3538;
    wire wire_3539;
    wire wire_3540;
    wire wire_3541;
    wire wire_3542;
    wire wire_3543;
    wire wire_3544;
    wire wire_3545;
    wire wire_3546;
    wire wire_3547;
    wire wire_3548;
    wire wire_3549;
    wire wire_3550;
    wire wire_3551;
    wire wire_3552;
    wire wire_3553;
    wire wire_3554;
    wire wire_3555;
    wire wire_3556;
    wire wire_3557;
    wire wire_3558;
    wire wire_3559;
    wire wire_3560;
    wire wire_3561;
    wire wire_3562;
    wire wire_3563;
    wire wire_3564;
    wire wire_3565;
    wire wire_3566;
    wire wire_3567;
    wire wire_3568;
    wire wire_3569;
    wire wire_3570;
    wire wire_3571;
    wire wire_3572;
    wire wire_3573;
    wire wire_3574;
    wire wire_3575;
    wire wire_3576;
    wire wire_3577;
    wire wire_3578;
    wire wire_3579;
    wire wire_3580;
    wire wire_3581;
    wire wire_3582;
    wire wire_3583;
    wire wire_3584;
    wire wire_3585;
    wire wire_3586;
    wire wire_3587;
    wire wire_3588;
    wire wire_3589;
    wire wire_3590;
    wire wire_3591;
    wire wire_3592;
    wire wire_3593;
    wire wire_3594;
    wire wire_3595;
    wire wire_3596;
    wire wire_3597;
    wire wire_3598;
    wire wire_3599;
    wire wire_3600;
    wire wire_3601;
    wire wire_3602;
    wire wire_3603;
    wire wire_3604;
    wire wire_3605;
    wire wire_3606;
    wire wire_3607;
    wire wire_3608;
    wire wire_3609;
    wire wire_3610;
    wire wire_3611;
    wire wire_3612;
    wire wire_3613;
    wire wire_3614;
    wire wire_3615;
    wire wire_3616;
    wire wire_3617;
    wire wire_3618;
    wire wire_3619;
    wire wire_3620;
    wire wire_3621;
    wire wire_3622;
    wire wire_3623;
    wire wire_3624;
    wire wire_3625;
    wire wire_3626;
    wire wire_3627;
    wire wire_3628;
    wire wire_3629;
    wire wire_3630;
    wire wire_3631;
    wire wire_3632;
    wire wire_3633;
    wire wire_3634;
    wire wire_3635;
    wire wire_3636;
    wire wire_3637;
    wire wire_3638;
    wire wire_3639;
    wire wire_3640;
    wire wire_3641;
    wire wire_3642;
    wire wire_3643;
    wire wire_3644;
    wire wire_3645;
    wire wire_3646;
    wire wire_3647;
    wire wire_3648;
    wire wire_3649;
    wire wire_3650;
    wire wire_3651;
    wire wire_3652;
    wire wire_3653;
    wire wire_3654;
    wire wire_3655;
    wire wire_3656;
    wire wire_3657;
    wire wire_3658;
    wire wire_3659;
    wire wire_3660;
    wire wire_3661;
    wire wire_3662;
    wire wire_3663;
    wire wire_3664;
    wire wire_3665;
    wire wire_3666;
    wire wire_3667;
    wire wire_3668;
    wire wire_3669;
    wire wire_3670;
    wire wire_3671;
    wire wire_3672;
    wire wire_3673;
    wire wire_3674;
    wire wire_3675;
    wire wire_3676;
    wire wire_3677;
    wire wire_3678;
    wire wire_3679;
    wire wire_3680;
    wire wire_3681;
    wire wire_3682;
    wire wire_3683;
    wire wire_3684;
    wire wire_3685;
    wire wire_3686;
    wire wire_3687;
    wire wire_3688;
    wire wire_3689;
    wire wire_3690;
    wire wire_3691;
    wire wire_3692;
    wire wire_3693;
    wire wire_3694;
    wire wire_3695;
    wire wire_3696;
    wire wire_3697;
    wire wire_3698;
    wire wire_3699;
    wire wire_3700;
    wire wire_3701;
    wire wire_3702;
    wire wire_3703;
    wire wire_3704;
    wire wire_3705;
    wire wire_3706;
    wire wire_3707;
    wire wire_3708;
    wire wire_3709;
    wire wire_3710;
    wire wire_3711;
    wire wire_3712;
    wire wire_3713;
    wire wire_3714;
    wire wire_3715;
    wire wire_3716;
    wire wire_3717;
    wire wire_3718;
    wire wire_3719;
    wire wire_3720;
    wire wire_3721;
    wire wire_3722;
    wire wire_3723;
    wire wire_3724;
    wire wire_3725;
    wire wire_3726;
    wire wire_3727;
    wire wire_3728;
    wire wire_3729;
    wire wire_3730;
    wire wire_3731;
    wire wire_3732;
    wire wire_3733;
    wire wire_3734;
    wire wire_3735;
    wire wire_3736;
    wire wire_3737;
    wire wire_3738;
    wire wire_3739;
    wire wire_3740;
    wire wire_3741;
    wire wire_3742;
    wire wire_3743;
    wire wire_3744;
    wire wire_3745;
    wire wire_3746;
    wire wire_3747;
    wire wire_3748;
    wire wire_3749;
    wire wire_3750;
    wire wire_3751;
    wire wire_3752;
    wire wire_3753;
    wire wire_3754;
    wire wire_3755;
    wire wire_3756;
    wire wire_3757;
    wire wire_3758;
    wire wire_3759;
    wire wire_3760;
    wire wire_3761;
    wire wire_3762;
    wire wire_3763;
    wire wire_3764;
    wire wire_3765;
    wire wire_3766;
    wire wire_3767;
    wire wire_3768;
    wire wire_3769;
    wire wire_3770;
    wire wire_3771;
    wire wire_3772;
    wire wire_3773;
    wire wire_3774;
    wire wire_3775;
    wire wire_3776;
    wire wire_3777;
    wire wire_3778;
    wire wire_3779;
    wire wire_3780;
    wire wire_3781;
    wire wire_3782;
    wire wire_3783;
    wire wire_3784;
    wire wire_3785;
    wire wire_3786;
    wire wire_3787;
    wire wire_3788;
    wire wire_3789;
    wire wire_3790;
    wire wire_3791;
    wire wire_3792;
    wire wire_3793;
    wire wire_3794;
    wire wire_3795;
    wire wire_3796;
    wire wire_3797;
    wire wire_3798;
    wire wire_3799;
    wire wire_3800;
    wire wire_3801;
    wire wire_3802;
    wire wire_3803;
    wire wire_3804;
    wire wire_3805;
    wire wire_3806;
    wire wire_3807;
    wire wire_3808;
    wire wire_3809;
    wire wire_3810;
    wire wire_3811;
    wire wire_3812;
    wire wire_3813;
    wire wire_3814;
    wire wire_3815;
    wire wire_3816;
    wire wire_3817;
    wire wire_3818;
    wire wire_3819;
    wire wire_3820;
    wire wire_3821;
    wire wire_3822;
    wire wire_3823;
    wire wire_3824;
    wire wire_3825;
    wire wire_3826;
    wire wire_3827;
    wire wire_3828;
    wire wire_3829;
    wire wire_3830;
    wire wire_3831;
    wire wire_3832;
    wire wire_3833;
    wire wire_3834;
    wire wire_3835;
    wire wire_3836;
    wire wire_3837;
    wire wire_3838;
    wire wire_3839;
    wire wire_3840;
    wire wire_3841;
    wire wire_3842;
    wire wire_3843;
    wire wire_3844;
    wire wire_3845;
    wire wire_3846;
    wire wire_3847;
    wire wire_3848;
    wire wire_3849;
    wire wire_3850;
    wire wire_3851;
    wire wire_3852;
    wire wire_3853;
    wire wire_3854;
    wire wire_3855;
    wire wire_3856;
    wire wire_3857;
    wire wire_3858;
    wire wire_3859;
    wire wire_3860;
    wire wire_3861;
    wire wire_3862;
    wire wire_3863;
    wire wire_3864;
    wire wire_3865;
    wire wire_3866;
    wire wire_3867;
    wire wire_3868;
    wire wire_3869;
    wire wire_3870;
    wire wire_3871;
    wire wire_3872;
    wire wire_3873;
    wire wire_3874;
    wire wire_3875;
    wire wire_3876;
    wire wire_3877;
    wire wire_3878;
    wire wire_3879;
    wire wire_3880;
    wire wire_3881;
    wire wire_3882;
    wire wire_3883;
    wire wire_3884;
    wire wire_3885;
    wire wire_3886;
    wire wire_3887;
    wire wire_3888;
    wire wire_3889;
    wire wire_3890;
    wire wire_3891;
    wire wire_3892;
    wire wire_3893;
    wire wire_3894;
    wire wire_3895;
    wire wire_3896;
    wire wire_3897;
    wire wire_3898;
    wire wire_3899;
    wire wire_3900;
    wire wire_3901;
    wire wire_3902;
    wire wire_3903;
    wire wire_3904;
    wire wire_3905;
    wire wire_3906;
    wire wire_3907;
    wire wire_3908;
    wire wire_3909;
    wire wire_3910;
    wire wire_3911;
    wire wire_3912;
    wire wire_3913;
    wire wire_3914;
    wire wire_3915;
    wire wire_3916;
    wire wire_3917;
    wire wire_3918;
    wire wire_3919;
    wire wire_3920;
    wire wire_3921;
    wire wire_3922;
    wire wire_3923;
    wire wire_3924;
    wire wire_3925;
    wire wire_3926;
    wire wire_3927;
    wire wire_3928;
    wire wire_3929;
    wire wire_3930;
    wire wire_3931;
    wire wire_3932;
    wire wire_3933;
    wire wire_3934;
    wire wire_3935;
    wire wire_3936;
    wire wire_3937;
    wire wire_3938;
    wire wire_3939;
    wire wire_3940;
    wire wire_3941;
    wire wire_3942;
    wire wire_3943;
    wire wire_3944;
    wire wire_3945;
    wire wire_3946;
    wire wire_3947;
    wire wire_3948;
    wire wire_3949;
    wire wire_3950;
    wire wire_3951;
    wire wire_3952;
    wire wire_3953;
    wire wire_3954;
    wire wire_3955;
    wire wire_3956;
    wire wire_3957;
    wire wire_3958;
    wire wire_3959;
    wire wire_3960;
    wire wire_3961;
    wire wire_3962;
    wire wire_3963;
    wire wire_3964;
    wire wire_3965;
    wire wire_3966;
    wire wire_3967;
    wire wire_3968;
    wire wire_3969;
    wire wire_3970;
    wire wire_3971;
    wire wire_3972;
    wire wire_3973;
    wire wire_3974;
    wire wire_3975;
    wire wire_3976;
    wire wire_3977;
    wire wire_3978;
    wire wire_3979;
    wire wire_3980;
    wire wire_3981;
    wire wire_3982;
    wire wire_3983;
    wire wire_3984;
    wire wire_3985;
    wire wire_3986;
    wire wire_3987;
    wire wire_3988;
    wire wire_3989;
    wire wire_3990;
    wire wire_3991;
    wire wire_3992;
    wire wire_3993;
    wire wire_3994;
    wire wire_3995;
    wire wire_3996;
    wire wire_3997;
    wire wire_3998;
    wire wire_3999;
    wire wire_4000;
    wire wire_4001;
    wire wire_4002;
    wire wire_4003;
    wire wire_4004;
    wire wire_4005;
    wire wire_4006;
    wire wire_4007;
    wire wire_4008;
    wire wire_4009;
    wire wire_4010;
    wire wire_4011;
    wire wire_4012;
    wire wire_4013;
    wire wire_4014;
    wire wire_4015;
    wire wire_4016;
    wire wire_4017;
    wire wire_4018;
    wire wire_4019;
    wire wire_4020;
    wire wire_4021;
    wire wire_4022;
    wire wire_4023;
    wire wire_4024;
    wire wire_4025;
    wire wire_4026;
    wire wire_4027;
    wire wire_4028;
    wire wire_4029;
    wire wire_4030;
    wire wire_4031;
    wire wire_4032;
    wire wire_4033;
    wire wire_4034;
    wire wire_4035;
    wire wire_4036;
    wire wire_4037;
    wire wire_4038;
    wire wire_4039;
    wire wire_4040;
    wire wire_4041;
    wire wire_4042;
    wire wire_4043;
    wire wire_4044;
    wire wire_4045;
    wire wire_4046;
    wire wire_4047;
    wire wire_4048;
    wire wire_4049;
    wire wire_4050;
    wire wire_4051;
    wire wire_4052;
    wire wire_4053;
    wire wire_4054;
    wire wire_4055;
    wire wire_4056;
    wire wire_4057;
    wire wire_4058;
    wire wire_4059;
    wire wire_4060;
    wire wire_4061;
    wire wire_4062;
    wire wire_4063;
    wire wire_4064;
    wire wire_4065;
    wire wire_4066;
    wire wire_4067;
    wire wire_4068;
    wire wire_4069;
    wire wire_4070;
    wire wire_4071;
    wire wire_4072;
    wire wire_4073;
    wire wire_4074;
    wire wire_4075;
    wire wire_4076;
    wire wire_4077;
    wire wire_4078;
    wire wire_4079;
    wire wire_4080;
    wire wire_4081;
    wire wire_4082;
    wire wire_4083;
    wire wire_4084;
    wire wire_4085;
    wire wire_4086;
    wire wire_4087;
    wire wire_4088;
    wire wire_4089;
    wire wire_4090;
    wire wire_4091;
    wire wire_4092;
    wire wire_4093;
    wire wire_4094;
    wire wire_4095;
    wire wire_4096;
    wire wire_4097;
    wire wire_4098;
    wire wire_4099;
    wire wire_4100;
    wire wire_4101;
    wire wire_4102;
    wire wire_4103;
    wire wire_4104;
    wire wire_4105;
    wire wire_4106;
    wire wire_4107;
    wire wire_4108;
    wire wire_4109;
    wire wire_4110;
    wire wire_4111;
    wire wire_4112;
    wire wire_4113;
    wire wire_4114;
    wire wire_4115;
    wire wire_4116;
    wire wire_4117;
    wire wire_4118;
    wire wire_4119;
    wire wire_4120;
    wire wire_4121;
    wire wire_4122;
    wire wire_4123;
    wire wire_4124;
    wire wire_4125;
    wire wire_4126;
    wire wire_4127;
    wire wire_4128;
    wire wire_4129;
    wire wire_4130;
    wire wire_4131;
    wire wire_4132;
    wire wire_4133;
    wire wire_4134;
    wire wire_4135;
    wire wire_4136;
    wire wire_4137;
    wire wire_4138;
    wire wire_4139;
    wire wire_4140;
    wire wire_4141;
    wire wire_4142;
    wire wire_4143;
    wire wire_4144;
    wire wire_4145;
    wire wire_4146;
    wire wire_4147;
    wire wire_4148;
    wire wire_4149;
    wire wire_4150;
    wire wire_4151;
    wire wire_4152;
    wire wire_4153;
    wire wire_4154;
    wire wire_4155;
    wire wire_4156;
    wire wire_4157;
    wire wire_4158;
    wire wire_4159;
    wire wire_4160;
    wire wire_4161;
    wire wire_4162;
    wire wire_4163;
    wire wire_4164;
    wire wire_4165;
    wire wire_4166;
    wire wire_4167;
    wire wire_4168;
    wire wire_4169;
    wire wire_4170;
    wire wire_4171;
    wire wire_4172;
    wire wire_4173;
    wire wire_4174;
    wire wire_4175;
    wire wire_4176;
    wire wire_4177;
    wire wire_4178;
    wire wire_4179;
    wire wire_4180;
    wire wire_4181;
    wire wire_4182;
    wire wire_4183;
    wire wire_4184;
    wire wire_4185;
    wire wire_4186;
    wire wire_4187;
    wire wire_4188;
    wire wire_4189;
    wire wire_4190;
    wire wire_4191;
    wire wire_4192;
    wire wire_4193;
    wire wire_4194;
    wire wire_4195;
    wire wire_4196;
    wire wire_4197;
    wire wire_4198;
    wire wire_4199;
    wire wire_4200;
    wire wire_4201;
    wire wire_4202;
    wire wire_4203;
    wire wire_4204;
    wire wire_4205;
    wire wire_4206;
    wire wire_4207;
    wire wire_4208;
    wire wire_4209;
    wire wire_4210;
    wire wire_4211;
    wire wire_4212;
    wire wire_4213;
    wire wire_4214;
    wire wire_4215;
    wire wire_4216;
    wire wire_4217;
    wire wire_4218;
    wire wire_4219;
    wire wire_4220;
    wire wire_4221;
    wire wire_4222;
    wire wire_4223;
    wire wire_4224;
    wire wire_4225;
    wire wire_4226;
    wire wire_4227;
    wire wire_4228;
    wire wire_4229;
    wire wire_4230;
    wire wire_4231;
    wire wire_4232;
    wire wire_4233;
    wire wire_4234;
    wire wire_4235;
    wire wire_4236;
    wire wire_4237;
    wire wire_4238;
    wire wire_4239;
    wire wire_4240;
    wire wire_4241;
    wire wire_4242;
    wire wire_4243;
    wire wire_4244;
    wire wire_4245;
    wire wire_4246;
    wire wire_4247;
    wire wire_4248;
    wire wire_4249;
    wire wire_4250;
    wire wire_4251;
    wire wire_4252;
    wire wire_4253;
    wire wire_4254;
    wire wire_4255;
    wire wire_4256;
    wire wire_4257;
    wire wire_4258;
    wire wire_4259;
    wire wire_4260;
    wire wire_4261;
    wire wire_4262;
    wire wire_4263;
    wire wire_4264;
    wire wire_4265;
    wire wire_4266;
    wire wire_4267;
    wire wire_4268;
    wire wire_4269;
    wire wire_4270;
    wire wire_4271;
    wire wire_4272;
    wire wire_4273;
    wire wire_4274;
    wire wire_4275;
    wire wire_4276;
    wire wire_4277;
    wire wire_4278;
    wire wire_4279;
    wire wire_4280;
    wire wire_4281;
    wire wire_4282;
    wire wire_4283;
    wire wire_4284;
    wire wire_4285;
    wire wire_4286;
    wire wire_4287;
    wire wire_4288;
    wire wire_4289;
    wire wire_4290;
    wire wire_4291;
    wire wire_4292;
    wire wire_4293;
    wire wire_4294;
    wire wire_4295;
    wire wire_4296;
    wire wire_4297;
    wire wire_4298;
    wire wire_4299;
    wire wire_4300;
    wire wire_4301;
    wire wire_4302;
    wire wire_4303;
    wire wire_4304;
    wire wire_4305;
    wire wire_4306;
    wire wire_4307;
    wire wire_4308;
    wire wire_4309;
    wire wire_4310;
    wire wire_4311;
    wire wire_4312;
    wire wire_4313;
    wire wire_4314;
    wire wire_4315;
    wire wire_4316;
    wire wire_4317;
    wire wire_4318;
    wire wire_4319;
    wire wire_4320;
    wire wire_4321;
    wire wire_4322;
    wire wire_4323;
    wire wire_4324;
    wire wire_4325;
    wire wire_4326;
    wire wire_4327;
    wire wire_4328;
    wire wire_4329;
    wire wire_4330;
    wire wire_4331;
    wire wire_4332;
    wire wire_4333;
    wire wire_4334;
    wire wire_4335;
    wire wire_4336;
    wire wire_4337;
    wire wire_4338;
    wire wire_4339;
    wire wire_4340;
    wire wire_4341;
    wire wire_4342;
    wire wire_4343;
    wire wire_4344;
    wire wire_4345;
    wire wire_4346;
    wire wire_4347;
    wire wire_4348;
    wire wire_4349;
    wire wire_4350;
    wire wire_4351;
    wire wire_4352;
    wire wire_4353;
    wire wire_4354;
    wire wire_4355;
    wire wire_4356;
    wire wire_4357;
    wire wire_4358;
    wire wire_4359;
    wire wire_4360;
    wire wire_4361;
    wire wire_4362;
    wire wire_4363;
    wire wire_4364;
    wire wire_4365;
    wire wire_4366;
    wire wire_4367;
    wire wire_4368;
    wire wire_4369;
    wire wire_4370;
    wire wire_4371;
    wire wire_4372;
    wire wire_4373;
    wire wire_4374;
    wire wire_4375;
    wire wire_4376;
    wire wire_4377;
    wire wire_4378;
    wire wire_4379;
    wire wire_4380;
    wire wire_4381;
    wire wire_4382;
    wire wire_4383;
    wire wire_4384;
    wire wire_4385;
    wire wire_4386;
    wire wire_4387;
    wire wire_4388;
    wire wire_4389;
    wire wire_4390;
    wire wire_4391;
    wire wire_4392;
    wire wire_4393;
    wire wire_4394;
    wire wire_4395;
    wire wire_4396;
    wire wire_4397;
    wire wire_4398;
    wire wire_4399;
    wire wire_4400;
    wire wire_4401;
    wire wire_4402;
    wire wire_4403;
    wire wire_4404;
    wire wire_4405;
    wire wire_4406;
    wire wire_4407;
    wire wire_4408;
    wire wire_4409;
    wire wire_4410;
    wire wire_4411;
    wire wire_4412;
    wire wire_4413;
    wire wire_4414;
    wire wire_4415;
    wire wire_4416;
    wire wire_4417;
    wire wire_4418;
    wire wire_4419;
    wire wire_4420;
    wire wire_4421;
    wire wire_4422;
    wire wire_4423;
    wire wire_4424;
    wire wire_4425;
    wire wire_4426;
    wire wire_4427;
    wire wire_4428;
    wire wire_4429;
    wire wire_4430;
    wire wire_4431;
    wire wire_4432;
    wire wire_4433;
    wire wire_4434;
    wire wire_4435;
    wire wire_4436;
    wire wire_4437;
    wire wire_4438;
    wire wire_4439;
    wire wire_4440;
    wire wire_4441;
    wire wire_4442;
    wire wire_4443;
    wire wire_4444;
    wire wire_4445;
    wire wire_4446;
    wire wire_4447;
    wire wire_4448;
    wire wire_4449;
    wire wire_4450;
    wire wire_4451;
    wire wire_4452;
    wire wire_4453;
    wire wire_4454;
    wire wire_4455;
    wire wire_4456;
    wire wire_4457;
    wire wire_4458;
    wire wire_4459;
    wire wire_4460;
    wire wire_4461;
    wire wire_4462;
    wire wire_4463;
    wire wire_4464;
    wire wire_4465;
    wire wire_4466;
    wire wire_4467;
    wire wire_4468;
    wire wire_4469;
    wire wire_4470;
    wire wire_4471;
    wire wire_4472;
    wire wire_4473;
    wire wire_4474;
    wire wire_4475;
    wire wire_4476;
    wire wire_4477;
    wire wire_4478;
    wire wire_4479;
    wire wire_4480;
    wire wire_4481;
    wire wire_4482;
    wire wire_4483;
    wire wire_4484;
    wire wire_4485;
    wire wire_4486;
    wire wire_4487;
    wire wire_4488;
    wire wire_4489;
    wire wire_4490;
    wire wire_4491;
    wire wire_4492;
    wire wire_4493;
    wire wire_4494;
    wire wire_4495;
    wire wire_4496;
    wire wire_4497;
    wire wire_4498;
    wire wire_4499;
    wire wire_4500;
    wire wire_4501;
    wire wire_4502;
    wire wire_4503;
    wire wire_4504;
    wire wire_4505;
    wire wire_4506;
    wire wire_4507;
    wire wire_4508;
    wire wire_4509;
    wire wire_4510;
    wire wire_4511;
    wire wire_4512;
    wire wire_4513;
    wire wire_4514;
    wire wire_4515;
    wire wire_4516;
    wire wire_4517;
    wire wire_4518;
    wire wire_4519;
    wire wire_4520;
    wire wire_4521;
    wire wire_4522;
    wire wire_4523;
    wire wire_4524;
    wire wire_4525;
    wire wire_4526;
    wire wire_4527;
    wire wire_4528;
    wire wire_4529;
    wire wire_4530;
    wire wire_4531;
    wire wire_4532;
    wire wire_4533;
    wire wire_4534;
    wire wire_4535;
    wire wire_4536;
    wire wire_4537;
    wire wire_4538;
    wire wire_4539;
    wire wire_4540;
    wire wire_4541;
    wire wire_4542;
    wire wire_4543;
    wire wire_4544;
    wire wire_4545;
    wire wire_4546;
    wire wire_4547;
    wire wire_4548;
    wire wire_4549;
    wire wire_4550;
    wire wire_4551;
    wire wire_4552;
    wire wire_4553;
    wire wire_4554;
    wire wire_4555;
    wire wire_4556;
    wire wire_4557;
    wire wire_4558;
    wire wire_4559;
    wire wire_4560;
    wire wire_4561;
    wire wire_4562;
    wire wire_4563;
    wire wire_4564;
    wire wire_4565;
    wire wire_4566;
    wire wire_4567;
    wire wire_4568;
    wire wire_4569;
    wire wire_4570;
    wire wire_4571;
    wire wire_4572;
    wire wire_4573;
    wire wire_4574;
    wire wire_4575;
    wire wire_4576;
    wire wire_4577;
    wire wire_4578;
    wire wire_4579;
    wire wire_4580;
    wire wire_4581;
    wire wire_4582;
    wire wire_4583;
    wire wire_4584;
    wire wire_4585;
    wire wire_4586;
    wire wire_4587;
    wire wire_4588;
    wire wire_4589;
    wire wire_4590;
    wire wire_4591;
    wire wire_4592;
    wire wire_4593;
    wire wire_4594;
    wire wire_4595;
    wire wire_4596;
    wire wire_4597;
    wire wire_4598;
    wire wire_4599;
    wire wire_4600;
    wire wire_4601;
    wire wire_4602;
    wire wire_4603;
    wire wire_4604;
    wire wire_4605;
    wire wire_4606;
    wire wire_4607;
    wire wire_4608;
    wire wire_4609;
    wire wire_4610;
    wire wire_4611;
    wire wire_4612;
    wire wire_4613;
    wire wire_4614;
    wire wire_4615;
    wire wire_4616;
    wire wire_4617;
    wire wire_4618;
    wire wire_4619;
    wire wire_4620;
    wire wire_4621;
    wire wire_4622;
    wire wire_4623;
    wire wire_4624;
    wire wire_4625;
    wire wire_4626;
    wire wire_4627;
    wire wire_4628;
    wire wire_4629;
    wire wire_4630;
    wire wire_4631;
    wire wire_4632;
    wire wire_4633;
    wire wire_4634;
    wire wire_4635;
    wire wire_4636;
    wire wire_4637;
    wire wire_4638;
    wire wire_4639;
    wire wire_4640;
    wire wire_4641;
    wire wire_4642;
    wire wire_4643;
    wire wire_4644;
    wire wire_4645;
    wire wire_4646;
    wire wire_4647;
    wire wire_4648;
    wire wire_4649;
    wire wire_4650;
    wire wire_4651;
    wire wire_4652;
    wire wire_4653;
    wire wire_4654;
    wire wire_4655;
    wire wire_4656;
    wire wire_4657;
    wire wire_4658;
    wire wire_4659;
    wire wire_4660;
    wire wire_4661;
    wire wire_4662;
    wire wire_4663;
    wire wire_4664;
    wire wire_4665;
    wire wire_4666;
    wire wire_4667;
    wire wire_4668;
    wire wire_4669;
    wire wire_4670;
    wire wire_4671;
    wire wire_4672;
    wire wire_4673;
    wire wire_4674;
    wire wire_4675;
    wire wire_4676;
    wire wire_4677;
    wire wire_4678;
    wire wire_4679;
    wire wire_4680;
    wire wire_4681;
    wire wire_4682;
    wire wire_4683;
    wire wire_4684;
    wire wire_4685;
    wire wire_4686;
    wire wire_4687;
    wire wire_4688;
    wire wire_4689;
    wire wire_4690;
    wire wire_4691;
    wire wire_4692;
    wire wire_4693;
    wire wire_4694;
    wire wire_4695;
    wire wire_4696;
    wire wire_4697;
    wire wire_4698;
    wire wire_4699;
    wire wire_4700;
    wire wire_4701;
    wire wire_4702;
    wire wire_4703;
    wire wire_4704;
    wire wire_4705;
    wire wire_4706;
    wire wire_4707;
    wire wire_4708;
    wire wire_4709;
    wire wire_4710;
    wire wire_4711;
    wire wire_4712;
    wire wire_4713;
    wire wire_4714;
    wire wire_4715;
    wire wire_4716;
    wire wire_4717;
    wire wire_4718;
    wire wire_4719;
    wire wire_4720;
    wire wire_4721;
    wire wire_4722;
    wire wire_4723;
    wire wire_4724;
    wire wire_4725;
    wire wire_4726;
    wire wire_4727;
    wire wire_4728;
    wire wire_4729;
    wire wire_4730;
    wire wire_4731;
    wire wire_4732;
    wire wire_4733;
    wire wire_4734;
    wire wire_4735;
    wire wire_4736;
    wire wire_4737;
    wire wire_4738;
    wire wire_4739;
    wire wire_4740;
    wire wire_4741;
    wire wire_4742;
    wire wire_4743;
    wire wire_4744;
    wire wire_4745;
    wire wire_4746;
    wire wire_4747;
    wire wire_4748;
    wire wire_4749;
    wire wire_4750;
    wire wire_4751;
    wire wire_4752;
    wire wire_4753;
    wire wire_4754;
    wire wire_4755;
    wire wire_4756;
    wire wire_4757;
    wire wire_4758;
    wire wire_4759;
    wire wire_4760;
    wire wire_4761;
    wire wire_4762;
    wire wire_4763;
    wire wire_4764;
    wire wire_4765;
    wire wire_4766;
    wire wire_4767;
    wire wire_4768;
    wire wire_4769;
    wire wire_4770;
    wire wire_4771;
    wire wire_4772;
    wire wire_4773;
    wire wire_4774;
    wire wire_4775;
    wire wire_4776;
    wire wire_4777;
    wire wire_4778;
    wire wire_4779;
    wire wire_4780;
    wire wire_4781;
    wire wire_4782;
    wire wire_4783;
    wire wire_4784;
    wire wire_4785;
    wire wire_4786;
    wire wire_4787;
    wire wire_4788;
    wire wire_4789;
    wire wire_4790;
    wire wire_4791;
    wire wire_4792;
    wire wire_4793;
    wire wire_4794;
    wire wire_4795;
    wire wire_4796;
    wire wire_4797;
    wire wire_4798;
    wire wire_4799;
    wire wire_4800;
    wire wire_4801;
    wire wire_4802;
    wire wire_4803;
    wire wire_4804;
    wire wire_4805;
    wire wire_4806;
    wire wire_4807;
    wire wire_4808;
    wire wire_4809;
    wire wire_4810;
    wire wire_4811;
    wire wire_4812;
    wire wire_4813;
    wire wire_4814;
    wire wire_4815;
    wire wire_4816;
    wire wire_4817;
    wire wire_4818;
    wire wire_4819;
    wire wire_4820;
    wire wire_4821;
    wire wire_4822;
    wire wire_4823;
    wire wire_4824;
    wire wire_4825;
    wire wire_4826;
    wire wire_4827;
    wire wire_4828;
    wire wire_4829;
    wire wire_4830;
    wire wire_4831;
    wire wire_4832;
    wire wire_4833;
    wire wire_4834;
    wire wire_4835;
    wire wire_4836;
    wire wire_4837;
    wire wire_4838;
    wire wire_4839;
    wire wire_4840;
    wire wire_4841;
    wire wire_4842;
    wire wire_4843;
    wire wire_4844;
    wire wire_4845;
    wire wire_4846;
    wire wire_4847;
    wire wire_4848;
    wire wire_4849;
    wire wire_4850;
    wire wire_4851;
    wire wire_4852;
    wire wire_4853;
    wire wire_4854;
    wire wire_4855;
    wire wire_4856;
    wire wire_4857;
    wire wire_4858;
    wire wire_4859;
    wire wire_4860;
    wire wire_4861;
    wire wire_4862;
    wire wire_4863;
    wire wire_4864;
    wire wire_4865;
    wire wire_4866;
    wire wire_4867;
    wire wire_4868;
    wire wire_4869;
    wire wire_4870;
    wire wire_4871;
    wire wire_4872;
    wire wire_4873;
    wire wire_4874;
    wire wire_4875;
    wire wire_4876;
    wire wire_4877;
    wire wire_4878;
    wire wire_4879;
    wire wire_4880;
    wire wire_4881;
    wire wire_4882;
    wire wire_4883;
    wire wire_4884;
    wire wire_4885;
    wire wire_4886;
    wire wire_4887;
    wire wire_4888;
    wire wire_4889;
    wire wire_4890;
    wire wire_4891;
    wire wire_4892;
    wire wire_4893;
    wire wire_4894;
    wire wire_4895;
    wire wire_4896;
    wire wire_4897;
    wire wire_4898;
    wire wire_4899;
    wire wire_4900;
    wire wire_4901;
    wire wire_4902;
    wire wire_4903;
    wire wire_4904;
    wire wire_4905;
    wire wire_4906;
    wire wire_4907;
    wire wire_4908;
    wire wire_4909;
    wire wire_4910;
    wire wire_4911;
    wire wire_4912;
    wire wire_4913;
    wire wire_4914;
    wire wire_4915;
    wire wire_4916;
    wire wire_4917;
    wire wire_4918;
    wire wire_4919;
    wire wire_4920;
    wire wire_4921;
    wire wire_4922;
    wire wire_4923;
    wire wire_4924;
    wire wire_4925;
    wire wire_4926;
    wire wire_4927;
    wire wire_4928;
    wire wire_4929;
    wire wire_4930;
    wire wire_4931;
    wire wire_4932;
    wire wire_4933;
    wire wire_4934;
    wire wire_4935;
    wire wire_4936;
    wire wire_4937;
    wire wire_4938;
    wire wire_4939;
    wire wire_4940;
    wire wire_4941;
    wire wire_4942;
    wire wire_4943;
    wire wire_4944;
    wire wire_4945;
    wire wire_4946;
    wire wire_4947;
    wire wire_4948;
    wire wire_4949;
    wire wire_4950;
    wire wire_4951;
    wire wire_4952;
    wire wire_4953;
    wire wire_4954;
    wire wire_4955;
    wire wire_4956;
    wire wire_4957;
    wire wire_4958;
    wire wire_4959;
    wire wire_4960;
    wire wire_4961;
    wire wire_4962;
    wire wire_4963;
    wire wire_4964;
    wire wire_4965;
    wire wire_4966;
    wire wire_4967;
    wire wire_4968;
    wire wire_4969;
    wire wire_4970;
    wire wire_4971;
    wire wire_4972;
    wire wire_4973;
    wire wire_4974;
    wire wire_4975;
    wire wire_4976;
    wire wire_4977;
    wire wire_4978;
    wire wire_4979;
    wire wire_4980;
    wire wire_4981;
    wire wire_4982;
    wire wire_4983;
    wire wire_4984;
    wire wire_4985;
    wire wire_4986;
    wire wire_4987;
    wire wire_4988;
    wire wire_4989;
    wire wire_4990;
    wire wire_4991;
    wire wire_4992;
    wire wire_4993;
    wire wire_4994;
    wire wire_4995;
    wire wire_4996;
    wire wire_4997;
    wire wire_4998;
    wire wire_4999;
    wire wire_5000;
    wire wire_5001;
    wire wire_5002;
    wire wire_5003;
    wire wire_5004;
    wire wire_5005;
    wire wire_5006;
    wire wire_5007;
    wire wire_5008;
    wire wire_5009;
    wire wire_5010;
    wire wire_5011;
    wire wire_5012;
    wire wire_5013;
    wire wire_5014;
    wire wire_5015;
    wire wire_5016;
    wire wire_5017;
    wire wire_5018;
    wire wire_5019;
    wire wire_5020;
    wire wire_5021;
    wire wire_5022;
    wire wire_5023;
    wire wire_5024;
    wire wire_5025;
    wire wire_5026;
    wire wire_5027;
    wire wire_5028;
    wire wire_5029;
    wire wire_5030;
    wire wire_5031;
    wire wire_5032;
    wire wire_5033;
    wire wire_5034;
    wire wire_5035;
    wire wire_5036;
    wire wire_5037;
    wire wire_5038;
    wire wire_5039;
    wire wire_5040;
    wire wire_5041;
    wire wire_5042;
    wire wire_5043;
    wire wire_5044;
    wire wire_5045;
    wire wire_5046;
    wire wire_5047;
    wire wire_5048;
    wire wire_5049;
    wire wire_5050;
    wire wire_5051;
    wire wire_5052;
    wire wire_5053;
    wire wire_5054;
    wire wire_5055;
    wire wire_5056;
    wire wire_5057;
    wire wire_5058;
    wire wire_5059;
    wire wire_5060;
    wire wire_5061;
    wire wire_5062;
    wire wire_5063;
    wire wire_5064;
    wire wire_5065;
    wire wire_5066;
    wire wire_5067;
    wire wire_5068;
    wire wire_5069;
    wire wire_5070;
    wire wire_5071;
    wire wire_5072;
    wire wire_5073;
    wire wire_5074;
    wire wire_5075;
    wire wire_5076;
    wire wire_5077;
    wire wire_5078;
    wire wire_5079;
    wire wire_5080;
    wire wire_5081;
    wire wire_5082;
    wire wire_5083;
    wire wire_5084;
    wire wire_5085;
    wire wire_5086;
    wire wire_5087;
    wire wire_5088;
    wire wire_5089;
    wire wire_5090;
    wire wire_5091;
    wire wire_5092;
    wire wire_5093;
    wire wire_5094;
    wire wire_5095;
    wire wire_5096;
    wire wire_5097;
    wire wire_5098;
    wire wire_5099;
    wire wire_5100;
    wire wire_5101;
    wire wire_5102;
    wire wire_5103;
    wire wire_5104;
    wire wire_5105;
    wire wire_5106;
    wire wire_5107;
    wire wire_5108;
    wire wire_5109;
    wire wire_5110;
    wire wire_5111;
    wire wire_5112;
    wire wire_5113;
    wire wire_5114;
    wire wire_5115;
    wire wire_5116;
    wire wire_5117;
    wire wire_5118;
    wire wire_5119;
    wire wire_5120;
    wire wire_5121;
    wire wire_5122;
    wire wire_5123;
    wire wire_5124;
    wire wire_5125;
    wire wire_5126;
    wire wire_5127;
    wire wire_5128;
    wire wire_5129;
    wire wire_5130;
    wire wire_5131;
    wire wire_5132;
    wire wire_5133;
    wire wire_5134;
    wire wire_5135;
    wire wire_5136;
    wire wire_5137;
    wire wire_5138;
    wire wire_5139;
    wire wire_5140;
    wire wire_5141;
    wire wire_5142;
    wire wire_5143;
    wire wire_5144;
    wire wire_5145;
    wire wire_5146;
    wire wire_5147;
    wire wire_5148;
    wire wire_5149;
    wire wire_5150;
    wire wire_5151;
    wire wire_5152;
    wire wire_5153;
    wire wire_5154;
    wire wire_5155;
    wire wire_5156;
    wire wire_5157;
    wire wire_5158;
    wire wire_5159;
    wire wire_5160;
    wire wire_5161;
    wire wire_5162;
    wire wire_5163;
    wire wire_5164;
    wire wire_5165;
    wire wire_5166;
    wire wire_5167;
    wire wire_5168;
    wire wire_5169;
    wire wire_5170;
    wire wire_5171;
    wire wire_5172;
    wire wire_5173;
    wire wire_5174;
    wire wire_5175;
    wire wire_5176;
    wire wire_5177;
    wire wire_5178;
    wire wire_5179;
    wire wire_5180;
    wire wire_5181;
    wire wire_5182;
    wire wire_5183;
    wire wire_5184;
    wire wire_5185;
    wire wire_5186;
    wire wire_5187;
    wire wire_5188;
    wire wire_5189;
    wire wire_5190;
    wire wire_5191;
    wire wire_5192;
    wire wire_5193;
    wire wire_5194;
    wire wire_5195;
    wire wire_5196;
    wire wire_5197;
    wire wire_5198;
    wire wire_5199;
    wire wire_5200;
    wire wire_5201;
    wire wire_5202;
    wire wire_5203;
    wire wire_5204;
    wire wire_5205;
    wire wire_5206;
    wire wire_5207;
    wire wire_5208;
    wire wire_5209;
    wire wire_5210;
    wire wire_5211;
    wire wire_5212;
    wire wire_5213;
    wire wire_5214;
    wire wire_5215;
    wire wire_5216;
    wire wire_5217;
    wire wire_5218;
    wire wire_5219;
    wire wire_5220;
    wire wire_5221;
    wire wire_5222;
    wire wire_5223;
    wire wire_5224;
    wire wire_5225;
    wire wire_5226;
    wire wire_5227;
    wire wire_5228;
    wire wire_5229;
    wire wire_5230;
    wire wire_5231;
    wire wire_5232;
    wire wire_5233;
    wire wire_5234;
    wire wire_5235;
    wire wire_5236;
    wire wire_5237;
    wire wire_5238;
    wire wire_5239;
    wire wire_5240;
    wire wire_5241;
    wire wire_5242;
    wire wire_5243;
    wire wire_5244;
    wire wire_5245;
    wire wire_5246;
    wire wire_5247;
    wire wire_5248;
    wire wire_5249;
    wire wire_5250;
    wire wire_5251;
    wire wire_5252;
    wire wire_5253;
    wire wire_5254;
    wire wire_5255;
    wire wire_5256;
    wire wire_5257;
    wire wire_5258;
    wire wire_5259;
    wire wire_5260;
    wire wire_5261;
    wire wire_5262;
    wire wire_5263;
    wire wire_5264;
    wire wire_5265;
    wire wire_5266;
    wire wire_5267;
    wire wire_5268;
    wire wire_5269;
    wire wire_5270;
    wire wire_5271;
    wire wire_5272;
    wire wire_5273;
    wire wire_5274;
    wire wire_5275;
    wire wire_5276;
    wire wire_5277;
    wire wire_5278;
    wire wire_5279;
    wire wire_5280;
    wire wire_5281;
    wire wire_5282;
    wire wire_5283;
    wire wire_5284;
    wire wire_5285;
    wire wire_5286;
    wire wire_5287;
    wire wire_5288;
    wire wire_5289;
    wire wire_5290;
    wire wire_5291;
    wire wire_5292;
    wire wire_5293;
    wire wire_5294;
    wire wire_5295;
    wire wire_5296;
    wire wire_5297;
    wire wire_5298;
    wire wire_5299;
    wire wire_5300;
    wire wire_5301;
    wire wire_5302;
    wire wire_5303;
    wire wire_5304;
    wire wire_5305;
    wire wire_5306;
    wire wire_5307;
    wire wire_5308;
    wire wire_5309;
    wire wire_5310;
    wire wire_5311;
    wire wire_5312;
    wire wire_5313;
    wire wire_5314;
    wire wire_5315;
    wire wire_5316;
    wire wire_5317;
    wire wire_5318;
    wire wire_5319;
    wire wire_5320;
    wire wire_5321;
    wire wire_5322;
    wire wire_5323;
    wire wire_5324;
    wire wire_5325;
    wire wire_5326;
    wire wire_5327;
    wire wire_5328;
    wire wire_5329;
    wire wire_5330;
    wire wire_5331;
    wire wire_5332;
    wire wire_5333;
    wire wire_5334;
    wire wire_5335;
    wire wire_5336;
    wire wire_5337;
    wire wire_5338;
    wire wire_5339;
    wire wire_5340;
    wire wire_5341;
    wire wire_5342;
    wire wire_5343;
    wire wire_5344;
    wire wire_5345;
    wire wire_5346;
    wire wire_5347;
    wire wire_5348;
    wire wire_5349;
    wire wire_5350;
    wire wire_5351;
    wire wire_5352;
    wire wire_5353;
    wire wire_5354;
    wire wire_5355;
    wire wire_5356;
    wire wire_5357;
    wire wire_5358;
    wire wire_5359;
    wire wire_5360;
    wire wire_5361;
    wire wire_5362;
    wire wire_5363;
    wire wire_5364;
    wire wire_5365;
    wire wire_5366;
    wire wire_5367;
    wire wire_5368;
    wire wire_5369;
    wire wire_5370;
    wire wire_5371;
    wire wire_5372;
    wire wire_5373;
    wire wire_5374;
    wire wire_5375;
    wire wire_5376;
    wire wire_5377;
    wire wire_5378;
    wire wire_5379;
    wire wire_5380;
    wire wire_5381;
    wire wire_5382;
    wire wire_5383;
    wire wire_5384;
    wire wire_5385;
    wire wire_5386;
    wire wire_5387;
    wire wire_5388;
    wire wire_5389;
    wire wire_5390;
    wire wire_5391;
    wire wire_5392;
    wire wire_5393;
    wire wire_5394;
    wire wire_5395;
    wire wire_5396;
    wire wire_5397;
    wire wire_5398;
    wire wire_5399;
    wire wire_5400;
    wire wire_5401;
    wire wire_5402;
    wire wire_5403;
    wire wire_5404;
    wire wire_5405;
    wire wire_5406;
    wire wire_5407;
    wire wire_5408;
    wire wire_5409;
    wire wire_5410;
    wire wire_5411;
    wire wire_5412;
    wire wire_5413;
    wire wire_5414;
    wire wire_5415;
    wire wire_5416;
    wire wire_5417;
    wire wire_5418;
    wire wire_5419;
    wire wire_5420;
    wire wire_5421;
    wire wire_5422;
    wire wire_5423;
    wire wire_5424;
    wire wire_5425;
    wire wire_5426;
    wire wire_5427;
    wire wire_5428;
    wire wire_5429;
    wire wire_5430;
    wire wire_5431;
    wire wire_5432;
    wire wire_5433;
    wire wire_5434;
    wire wire_5435;
    wire wire_5436;
    wire wire_5437;
    wire wire_5438;
    wire wire_5439;
    wire wire_5440;
    wire wire_5441;
    wire wire_5442;
    wire wire_5443;
    wire wire_5444;
    wire wire_5445;
    wire wire_5446;
    wire wire_5447;
    wire wire_5448;
    wire wire_5449;
    wire wire_5450;
    wire wire_5451;
    wire wire_5452;
    wire wire_5453;
    wire wire_5454;
    wire wire_5455;
    wire wire_5456;
    wire wire_5457;
    wire wire_5458;
    wire wire_5459;
    wire wire_5460;
    wire wire_5461;
    wire wire_5462;
    wire wire_5463;
    wire wire_5464;
    wire wire_5465;
    wire wire_5466;
    wire wire_5467;
    wire wire_5468;
    wire wire_5469;
    wire wire_5470;
    wire wire_5471;
    wire wire_5472;
    wire wire_5473;
    wire wire_5474;
    wire wire_5475;
    wire wire_5476;
    wire wire_5477;
    wire wire_5478;
    wire wire_5479;
    wire wire_5480;
    wire wire_5481;
    wire wire_5482;
    wire wire_5483;
    wire wire_5484;
    wire wire_5485;
    wire wire_5486;
    wire wire_5487;
    wire wire_5488;
    wire wire_5489;
    wire wire_5490;
    wire wire_5491;
    wire wire_5492;
    wire wire_5493;
    wire wire_5494;
    wire wire_5495;
    wire wire_5496;
    wire wire_5497;
    wire wire_5498;
    wire wire_5499;
    wire wire_5500;
    wire wire_5501;
    wire wire_5502;
    wire wire_5503;
    wire wire_5504;
    wire wire_5505;
    wire wire_5506;
    wire wire_5507;
    wire wire_5508;
    wire wire_5509;
    wire wire_5510;
    wire wire_5511;
    wire wire_5512;
    wire wire_5513;
    wire wire_5514;
    wire wire_5515;
    wire wire_5516;
    wire wire_5517;
    wire wire_5518;
    wire wire_5519;
    wire wire_5520;
    wire wire_5521;
    wire wire_5522;
    wire wire_5523;
    wire wire_5524;
    wire wire_5525;
    wire wire_5526;
    wire wire_5527;
    wire wire_5528;
    wire wire_5529;
    wire wire_5530;
    wire wire_5531;
    wire wire_5532;
    wire wire_5533;
    wire wire_5534;
    wire wire_5535;
    wire wire_5536;
    wire wire_5537;
    wire wire_5538;
    wire wire_5539;
    wire wire_5540;
    wire wire_5541;
    wire wire_5542;
    wire wire_5543;
    wire wire_5544;
    wire wire_5545;
    wire wire_5546;
    wire wire_5547;
    wire wire_5548;
    wire wire_5549;
    wire wire_5550;
    wire wire_5551;
    wire wire_5552;
    wire wire_5553;
    wire wire_5554;
    wire wire_5555;
    wire wire_5556;
    wire wire_5557;
    wire wire_5558;
    wire wire_5559;
    wire wire_5560;
    wire wire_5561;
    wire wire_5562;
    wire wire_5563;
    wire wire_5564;
    wire wire_5565;
    wire wire_5566;
    wire wire_5567;
    wire wire_5568;
    wire wire_5569;
    wire wire_5570;
    wire wire_5571;
    wire wire_5572;
    wire wire_5573;
    wire wire_5574;
    wire wire_5575;
    wire wire_5576;
    wire wire_5577;
    wire wire_5578;
    wire wire_5579;
    wire wire_5580;
    wire wire_5581;
    wire wire_5582;
    wire wire_5583;
    wire wire_5584;
    wire wire_5585;
    wire wire_5586;
    wire wire_5587;
    wire wire_5588;
    wire wire_5589;
    wire wire_5590;
    wire wire_5591;
    wire wire_5592;
    wire wire_5593;
    wire wire_5594;
    wire wire_5595;
    wire wire_5596;
    wire wire_5597;
    wire wire_5598;
    wire wire_5599;
    wire wire_5600;
    wire wire_5601;
    wire wire_5602;
    wire wire_5603;
    wire wire_5604;
    wire wire_5605;
    wire wire_5606;
    wire wire_5607;
    wire wire_5608;
    wire wire_5609;
    wire wire_5610;
    wire wire_5611;
    wire wire_5612;
    wire wire_5613;
    wire wire_5614;
    wire wire_5615;
    wire wire_5616;
    wire wire_5617;
    wire wire_5618;
    wire wire_5619;
    wire wire_5620;
    wire wire_5621;
    wire wire_5622;
    wire wire_5623;
    wire wire_5624;
    wire wire_5625;
    wire wire_5626;
    wire wire_5627;
    wire wire_5628;
    wire wire_5629;
    wire wire_5630;
    wire wire_5631;
    wire wire_5632;
    wire wire_5633;
    wire wire_5634;
    wire wire_5635;
    wire wire_5636;
    wire wire_5637;
    wire wire_5638;
    wire wire_5639;
    wire wire_5640;
    wire wire_5641;
    wire wire_5642;
    wire wire_5643;
    wire wire_5644;
    wire wire_5645;
    wire wire_5646;
    wire wire_5647;
    wire wire_5648;
    wire wire_5649;
    wire wire_5650;
    wire wire_5651;
    wire wire_5652;
    wire wire_5653;
    wire wire_5654;
    wire wire_5655;
    wire wire_5656;
    wire wire_5657;
    wire wire_5658;
    wire wire_5659;
    wire wire_5660;
    wire wire_5661;
    wire wire_5662;
    wire wire_5663;
    wire wire_5664;
    wire wire_5665;
    wire wire_5666;
    wire wire_5667;
    wire wire_5668;
    wire wire_5669;
    wire wire_5670;
    wire wire_5671;
    wire wire_5672;
    wire wire_5673;
    wire wire_5674;
    wire wire_5675;
    wire wire_5676;
    wire wire_5677;
    wire wire_5678;
    wire wire_5679;
    wire wire_5680;
    wire wire_5681;
    wire wire_5682;
    wire wire_5683;
    wire wire_5684;
    wire wire_5685;
    wire wire_5686;
    wire wire_5687;
    wire wire_5688;
    wire wire_5689;
    wire wire_5690;
    wire wire_5691;
    wire wire_5692;
    wire wire_5693;
    wire wire_5694;
    wire wire_5695;
    wire wire_5696;
    wire wire_5697;
    wire wire_5698;
    wire wire_5699;
    wire wire_5700;
    wire wire_5701;
    wire wire_5702;
    wire wire_5703;
    wire wire_5704;
    wire wire_5705;
    wire wire_5706;
    wire wire_5707;
    wire wire_5708;
    wire wire_5709;
    wire wire_5710;
    wire wire_5711;
    wire wire_5712;
    wire wire_5713;
    wire wire_5714;
    wire wire_5715;
    wire wire_5716;
    wire wire_5717;
    wire wire_5718;
    wire wire_5719;
    wire wire_5720;
    wire wire_5721;
    wire wire_5722;
    wire wire_5723;
    wire wire_5724;
    wire wire_5725;
    wire wire_5726;
    wire wire_5727;
    wire wire_5728;
    wire wire_5729;
    wire wire_5730;
    wire wire_5731;
    wire wire_5732;
    wire wire_5733;
    wire wire_5734;
    wire wire_5735;
    wire wire_5736;
    wire wire_5737;
    wire wire_5738;
    wire wire_5739;
    wire wire_5740;
    wire wire_5741;
    wire wire_5742;
    wire wire_5743;
    wire wire_5744;
    wire wire_5745;
    wire wire_5746;
    wire wire_5747;
    wire wire_5748;
    wire wire_5749;
    wire wire_5750;
    wire wire_5751;
    wire wire_5752;
    wire wire_5753;
    wire wire_5754;
    wire wire_5755;
    wire wire_5756;
    wire wire_5757;
    wire wire_5758;
    wire wire_5759;
    wire wire_5760;
    wire wire_5761;
    wire wire_5762;
    wire wire_5763;
    wire wire_5764;
    wire wire_5765;
    wire wire_5766;
    wire wire_5767;
    wire wire_5768;
    wire wire_5769;
    wire wire_5770;
    wire wire_5771;
    wire wire_5772;
    wire wire_5773;
    wire wire_5774;
    wire wire_5775;
    wire wire_5776;
    wire wire_5777;
    wire wire_5778;
    wire wire_5779;
    wire wire_5780;
    wire wire_5781;
    wire wire_5782;
    wire wire_5783;
    wire wire_5784;
    wire wire_5785;
    wire wire_5786;
    wire wire_5787;
    wire wire_5788;
    wire wire_5789;
    wire wire_5790;
    wire wire_5791;
    wire wire_5792;
    wire wire_5793;
    wire wire_5794;
    wire wire_5795;
    wire wire_5796;
    wire wire_5797;
    wire wire_5798;
    wire wire_5799;
    wire wire_5800;
    wire wire_5801;
    wire wire_5802;
    wire wire_5803;
    wire wire_5804;
    wire wire_5805;
    wire wire_5806;
    wire wire_5807;
    wire wire_5808;
    wire wire_5809;
    wire wire_5810;
    wire wire_5811;
    wire wire_5812;
    wire wire_5813;
    wire wire_5814;
    wire wire_5815;
    wire wire_5816;
    wire wire_5817;
    wire wire_5818;
    wire wire_5819;
    wire wire_5820;
    wire wire_5821;
    wire wire_5822;
    wire wire_5823;
    wire wire_5824;
    wire wire_5825;
    wire wire_5826;
    wire wire_5827;
    wire wire_5828;
    wire wire_5829;
    wire wire_5830;
    wire wire_5831;
    wire wire_5832;
    wire wire_5833;
    wire wire_5834;
    wire wire_5835;
    wire wire_5836;
    wire wire_5837;
    wire wire_5838;
    wire wire_5839;
    wire wire_5840;
    wire wire_5841;
    wire wire_5842;
    wire wire_5843;
    wire wire_5844;
    wire wire_5845;
    wire wire_5846;
    wire wire_5847;
    wire wire_5848;
    wire wire_5849;
    wire wire_5850;
    wire wire_5851;
    wire wire_5852;
    wire wire_5853;
    wire wire_5854;
    wire wire_5855;
    wire wire_5856;
    wire wire_5857;
    wire wire_5858;
    wire wire_5859;
    wire wire_5860;
    wire wire_5861;
    wire wire_5862;
    wire wire_5863;
    wire wire_5864;
    wire wire_5865;
    wire wire_5866;
    wire wire_5867;
    wire wire_5868;
    wire wire_5869;
    wire wire_5870;
    wire wire_5871;
    wire wire_5872;
    wire wire_5873;
    wire wire_5874;
    wire wire_5875;
    wire wire_5876;
    wire wire_5877;
    wire wire_5878;
    wire wire_5879;
    wire wire_5880;
    wire wire_5881;
    wire wire_5882;
    wire wire_5883;
    wire wire_5884;
    wire wire_5885;
    wire wire_5886;
    wire wire_5887;
    wire wire_5888;
    wire wire_5889;
    wire wire_5890;
    wire wire_5891;
    wire wire_5892;
    wire wire_5893;
    wire wire_5894;
    wire wire_5895;
    wire wire_5896;
    wire wire_5897;
    wire wire_5898;
    wire wire_5899;
    wire wire_5900;
    wire wire_5901;
    wire wire_5902;
    wire wire_5903;
    wire wire_5904;
    wire wire_5905;
    wire wire_5906;
    wire wire_5907;
    wire wire_5908;
    wire wire_5909;
    wire wire_5910;
    wire wire_5911;
    wire wire_5912;
    wire wire_5913;
    wire wire_5914;
    wire wire_5915;
    wire wire_5916;
    wire wire_5917;
    wire wire_5918;
    wire wire_5919;
    wire wire_5920;
    wire wire_5921;
    wire wire_5922;
    wire wire_5923;
    wire wire_5924;
    wire wire_5925;
    wire wire_5926;
    wire wire_5927;
    wire wire_5928;
    wire wire_5929;
    wire wire_5930;
    wire wire_5931;
    wire wire_5932;
    wire wire_5933;
    wire wire_5934;
    wire wire_5935;
    wire wire_5936;
    wire wire_5937;
    wire wire_5938;
    wire wire_5939;
    wire wire_5940;
    wire wire_5941;
    wire wire_5942;
    wire wire_5943;
    wire wire_5944;
    wire wire_5945;
    wire wire_5946;
    wire wire_5947;
    wire wire_5948;
    wire wire_5949;
    wire wire_5950;
    wire wire_5951;
    wire wire_5952;
    wire wire_5953;
    wire wire_5954;
    wire wire_5955;
    wire wire_5956;
    wire wire_5957;
    wire wire_5958;
    wire wire_5959;
    wire wire_5960;
    wire wire_5961;
    wire wire_5962;
    wire wire_5963;
    wire wire_5964;
    wire wire_5965;
    wire wire_5966;
    wire wire_5967;
    wire wire_5968;
    wire wire_5969;
    wire wire_5970;
    wire wire_5971;
    wire wire_5972;
    wire wire_5973;
    wire wire_5974;
    wire wire_5975;
    wire wire_5976;
    wire wire_5977;
    wire wire_5978;
    wire wire_5979;
    wire wire_5980;
    wire wire_5981;
    wire wire_5982;
    wire wire_5983;
    wire wire_5984;
    wire wire_5985;
    wire wire_5986;
    wire wire_5987;
    wire wire_5988;
    wire wire_5989;
    wire wire_5990;
    wire wire_5991;
    wire wire_5992;
    wire wire_5993;
    wire wire_5994;
    wire wire_5995;
    wire wire_5996;
    wire wire_5997;
    wire wire_5998;
    wire wire_5999;
    wire wire_6000;
    wire wire_6001;
    wire wire_6002;
    wire wire_6003;
    wire wire_6004;
    wire wire_6005;
    wire wire_6006;
    wire wire_6007;
    wire wire_6008;
    wire wire_6009;
    wire wire_6010;
    wire wire_6011;
    wire wire_6012;
    wire wire_6013;
    wire wire_6014;
    wire wire_6015;
    wire wire_6016;
    wire wire_6017;
    wire wire_6018;
    wire wire_6019;
    wire wire_6020;
    wire wire_6021;
    wire wire_6022;
    wire wire_6023;
    wire wire_6024;
    wire wire_6025;
    wire wire_6026;
    wire wire_6027;
    wire wire_6028;
    wire wire_6029;
    wire wire_6030;
    wire wire_6031;
    wire wire_6032;
    wire wire_6033;
    wire wire_6034;
    wire wire_6035;
    wire wire_6036;
    wire wire_6037;
    wire wire_6038;
    wire wire_6039;
    wire wire_6040;
    wire wire_6041;
    wire wire_6042;
    wire wire_6043;
    wire wire_6044;
    wire wire_6045;
    wire wire_6046;
    wire wire_6047;
    wire wire_6048;
    wire wire_6049;
    wire wire_6050;
    wire wire_6051;
    wire wire_6052;
    wire wire_6053;
    wire wire_6054;
    wire wire_6055;
    wire wire_6056;
    wire wire_6057;
    wire wire_6058;
    wire wire_6059;
    wire wire_6060;
    wire wire_6061;
    wire wire_6062;
    wire wire_6063;
    wire wire_6064;
    wire wire_6065;
    wire wire_6066;
    wire wire_6067;
    wire wire_6068;
    wire wire_6069;
    wire wire_6070;
    wire wire_6071;
    wire wire_6072;
    wire wire_6073;
    wire wire_6074;
    wire wire_6075;
    wire wire_6076;
    wire wire_6077;
    wire wire_6078;
    wire wire_6079;
    wire wire_6080;
    wire wire_6081;
    wire wire_6082;
    wire wire_6083;
    wire wire_6084;
    wire wire_6085;
    wire wire_6086;
    wire wire_6087;
    wire wire_6088;
    wire wire_6089;
    wire wire_6090;
    wire wire_6091;
    wire wire_6092;
    wire wire_6093;
    wire wire_6094;
    wire wire_6095;
    wire wire_6096;
    wire wire_6097;
    wire wire_6098;
    wire wire_6099;
    wire wire_6100;
    wire wire_6101;
    wire wire_6102;
    wire wire_6103;
    wire wire_6104;
    wire wire_6105;
    wire wire_6106;
    wire wire_6107;
    wire wire_6108;
    wire wire_6109;
    wire wire_6110;
    wire wire_6111;
    wire wire_6112;
    wire wire_6113;
    wire wire_6114;
    wire wire_6115;
    wire wire_6116;
    wire wire_6117;
    wire wire_6118;
    wire wire_6119;
    wire wire_6120;
    wire wire_6121;
    wire wire_6122;
    wire wire_6123;
    wire wire_6124;
    wire wire_6125;
    wire wire_6126;
    wire wire_6127;
    wire wire_6128;
    wire wire_6129;
    wire wire_6130;
    wire wire_6131;
    wire wire_6132;
    wire wire_6133;
    wire wire_6134;
    wire wire_6135;
    wire wire_6136;
    wire wire_6137;
    wire wire_6138;
    wire wire_6139;
    wire wire_6140;
    wire wire_6141;
    wire wire_6142;
    wire wire_6143;
    wire wire_6144;
    wire wire_6145;
    wire wire_6146;
    wire wire_6147;
    wire wire_6148;
    wire wire_6149;
    wire wire_6150;
    wire wire_6151;
    wire wire_6152;
    wire wire_6153;
    wire wire_6154;
    wire wire_6155;
    wire wire_6156;
    wire wire_6157;
    wire wire_6158;
    wire wire_6159;
    wire wire_6160;
    wire wire_6161;
    wire wire_6162;
    wire wire_6163;
    wire wire_6164;
    wire wire_6165;
    wire wire_6166;
    wire wire_6167;
    wire wire_6168;
    wire wire_6169;
    wire wire_6170;
    wire wire_6171;
    wire wire_6172;
    wire wire_6173;
    wire wire_6174;
    wire wire_6175;
    wire wire_6176;
    wire wire_6177;
    wire wire_6178;
    wire wire_6179;
    wire wire_6180;
    wire wire_6181;
    wire wire_6182;
    wire wire_6183;
    wire wire_6184;
    wire wire_6185;
    wire wire_6186;
    wire wire_6187;
    wire wire_6188;
    wire wire_6189;
    wire wire_6190;
    wire wire_6191;
    wire wire_6192;
    wire wire_6193;
    wire wire_6194;
    wire wire_6195;
    wire wire_6196;
    wire wire_6197;
    wire wire_6198;
    wire wire_6199;


    // FPGA IO TILES DECLARE
    wire [339:0] io_tile_1_0_chanxy_in;
    wire [99:0] io_tile_1_0_chanxy_out;
    wire [127:0] io_tile_1_0_ipin_in;
    wire [7:0] io_tile_1_0_opin_out;
    io_tile_sp_0 io_tile_1_0(
            .io_chanxy_in(io_tile_1_0_chanxy_in),
            .io_chanxy_out(io_tile_1_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[12:7]),
            .io_io_input(left_in[7:0]),
            .io_io_output(left_out[7:0]),
            .io_ipin_in(io_tile_1_0_ipin_in),
            .io_opin_out(io_tile_1_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [359:0] io_tile_2_0_chanxy_in;
    wire [39:0] io_tile_2_0_chanxy_out;
    wire [127:0] io_tile_2_0_ipin_in;
    wire [7:0] io_tile_2_0_opin_out;
    io_tile_sp_1 io_tile_2_0(
            .io_chanxy_in(io_tile_2_0_chanxy_in),
            .io_chanxy_out(io_tile_2_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[61:56]),
            .io_io_input(left_in[15:8]),
            .io_io_output(left_out[15:8]),
            .io_ipin_in(io_tile_2_0_ipin_in),
            .io_opin_out(io_tile_2_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [359:0] io_tile_3_0_chanxy_in;
    wire [39:0] io_tile_3_0_chanxy_out;
    wire [127:0] io_tile_3_0_ipin_in;
    wire [7:0] io_tile_3_0_opin_out;
    io_tile_sp_2 io_tile_3_0(
            .io_chanxy_in(io_tile_3_0_chanxy_in),
            .io_chanxy_out(io_tile_3_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[108:103]),
            .io_io_input(left_in[23:16]),
            .io_io_output(left_out[23:16]),
            .io_ipin_in(io_tile_3_0_ipin_in),
            .io_opin_out(io_tile_3_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [359:0] io_tile_4_0_chanxy_in;
    wire [39:0] io_tile_4_0_chanxy_out;
    wire [127:0] io_tile_4_0_ipin_in;
    wire [7:0] io_tile_4_0_opin_out;
    io_tile_sp_3 io_tile_4_0(
            .io_chanxy_in(io_tile_4_0_chanxy_in),
            .io_chanxy_out(io_tile_4_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[155:150]),
            .io_io_input(left_in[31:24]),
            .io_io_output(left_out[31:24]),
            .io_ipin_in(io_tile_4_0_ipin_in),
            .io_opin_out(io_tile_4_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [339:0] io_tile_5_0_chanxy_in;
    wire [99:0] io_tile_5_0_chanxy_out;
    wire [127:0] io_tile_5_0_ipin_in;
    wire [7:0] io_tile_5_0_opin_out;
    io_tile_sp_4 io_tile_5_0(
            .io_chanxy_in(io_tile_5_0_chanxy_in),
            .io_chanxy_out(io_tile_5_0_chanxy_out),
            .io_configs_in(configs_in[31:0]),
            .io_configs_en(configs_en[202:197]),
            .io_io_input(left_in[39:32]),
            .io_io_output(left_out[39:32]),
            .io_ipin_in(io_tile_5_0_ipin_in),
            .io_opin_out(io_tile_5_0_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_1_6_ipin_in;
    wire [7:0] io_tile_1_6_opin_out;
    io_tile_sp_5 io_tile_1_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[7:7]),
            .io_io_input(right_in[7:0]),
            .io_io_output(right_out[7:0]),
            .io_ipin_in(io_tile_1_6_ipin_in),
            .io_opin_out(io_tile_1_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_2_6_ipin_in;
    wire [7:0] io_tile_2_6_opin_out;
    io_tile_sp_6 io_tile_2_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[56:56]),
            .io_io_input(right_in[15:8]),
            .io_io_output(right_out[15:8]),
            .io_ipin_in(io_tile_2_6_ipin_in),
            .io_opin_out(io_tile_2_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_3_6_ipin_in;
    wire [7:0] io_tile_3_6_opin_out;
    io_tile_sp_7 io_tile_3_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[103:103]),
            .io_io_input(right_in[23:16]),
            .io_io_output(right_out[23:16]),
            .io_ipin_in(io_tile_3_6_ipin_in),
            .io_opin_out(io_tile_3_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_4_6_ipin_in;
    wire [7:0] io_tile_4_6_opin_out;
    io_tile_sp_8 io_tile_4_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[150:150]),
            .io_io_input(right_in[31:24]),
            .io_io_output(right_out[31:24]),
            .io_ipin_in(io_tile_4_6_ipin_in),
            .io_opin_out(io_tile_4_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_5_6_ipin_in;
    wire [7:0] io_tile_5_6_opin_out;
    io_tile_sp_9 io_tile_5_6(
            .io_configs_in(configs_in[223:192]),
            .io_configs_en(configs_en[197:197]),
            .io_io_input(right_in[39:32]),
            .io_io_output(right_out[39:32]),
            .io_ipin_in(io_tile_5_6_ipin_in),
            .io_opin_out(io_tile_5_6_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [355:0] io_tile_0_1_chanxy_in;
    wire [99:0] io_tile_0_1_chanxy_out;
    wire [127:0] io_tile_0_1_ipin_in;
    wire [7:0] io_tile_0_1_opin_out;
    io_tile_sp_10 io_tile_0_1(
            .io_chanxy_in(io_tile_0_1_chanxy_in),
            .io_chanxy_out(io_tile_0_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[6:0]),
            .io_io_input(bot_in[7:0]),
            .io_io_output(bot_out[7:0]),
            .io_ipin_in(io_tile_0_1_ipin_in),
            .io_opin_out(io_tile_0_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [375:0] io_tile_0_2_chanxy_in;
    wire [39:0] io_tile_0_2_chanxy_out;
    wire [127:0] io_tile_0_2_ipin_in;
    wire [7:0] io_tile_0_2_opin_out;
    io_tile_sp_11 io_tile_0_2(
            .io_chanxy_in(io_tile_0_2_chanxy_in),
            .io_chanxy_out(io_tile_0_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[5:0]),
            .io_io_input(bot_in[15:8]),
            .io_io_output(bot_out[15:8]),
            .io_ipin_in(io_tile_0_2_ipin_in),
            .io_opin_out(io_tile_0_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [375:0] io_tile_0_3_chanxy_in;
    wire [39:0] io_tile_0_3_chanxy_out;
    wire [127:0] io_tile_0_3_ipin_in;
    wire [7:0] io_tile_0_3_opin_out;
    io_tile_sp_12 io_tile_0_3(
            .io_chanxy_in(io_tile_0_3_chanxy_in),
            .io_chanxy_out(io_tile_0_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[5:0]),
            .io_io_input(bot_in[23:16]),
            .io_io_output(bot_out[23:16]),
            .io_ipin_in(io_tile_0_3_ipin_in),
            .io_opin_out(io_tile_0_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [375:0] io_tile_0_4_chanxy_in;
    wire [39:0] io_tile_0_4_chanxy_out;
    wire [127:0] io_tile_0_4_ipin_in;
    wire [7:0] io_tile_0_4_opin_out;
    io_tile_sp_13 io_tile_0_4(
            .io_chanxy_in(io_tile_0_4_chanxy_in),
            .io_chanxy_out(io_tile_0_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[5:0]),
            .io_io_input(bot_in[31:24]),
            .io_io_output(bot_out[31:24]),
            .io_ipin_in(io_tile_0_4_ipin_in),
            .io_opin_out(io_tile_0_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [355:0] io_tile_0_5_chanxy_in;
    wire [99:0] io_tile_0_5_chanxy_out;
    wire [127:0] io_tile_0_5_ipin_in;
    wire [7:0] io_tile_0_5_opin_out;
    io_tile_sp_14 io_tile_0_5(
            .io_chanxy_in(io_tile_0_5_chanxy_in),
            .io_chanxy_out(io_tile_0_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[6:0]),
            .io_io_input(bot_in[39:32]),
            .io_io_output(bot_out[39:32]),
            .io_ipin_in(io_tile_0_5_ipin_in),
            .io_opin_out(io_tile_0_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_6_1_ipin_in;
    wire [7:0] io_tile_6_1_opin_out;
    io_tile_sp_15 io_tile_6_1(
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[244:244]),
            .io_io_input(top_in[7:0]),
            .io_io_output(top_out[7:0]),
            .io_ipin_in(io_tile_6_1_ipin_in),
            .io_opin_out(io_tile_6_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_6_2_ipin_in;
    wire [7:0] io_tile_6_2_opin_out;
    io_tile_sp_16 io_tile_6_2(
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[244:244]),
            .io_io_input(top_in[15:8]),
            .io_io_output(top_out[15:8]),
            .io_ipin_in(io_tile_6_2_ipin_in),
            .io_opin_out(io_tile_6_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_6_3_ipin_in;
    wire [7:0] io_tile_6_3_opin_out;
    io_tile_sp_17 io_tile_6_3(
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[244:244]),
            .io_io_input(top_in[23:16]),
            .io_io_output(top_out[23:16]),
            .io_ipin_in(io_tile_6_3_ipin_in),
            .io_opin_out(io_tile_6_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_6_4_ipin_in;
    wire [7:0] io_tile_6_4_opin_out;
    io_tile_sp_18 io_tile_6_4(
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[244:244]),
            .io_io_input(top_in[31:24]),
            .io_io_output(top_out[31:24]),
            .io_ipin_in(io_tile_6_4_ipin_in),
            .io_opin_out(io_tile_6_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );

    wire [127:0] io_tile_6_5_ipin_in;
    wire [7:0] io_tile_6_5_opin_out;
    io_tile_sp_19 io_tile_6_5(
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[244:244]),
            .io_io_input(top_in[39:32]),
            .io_io_output(top_out[39:32]),
            .io_ipin_in(io_tile_6_5_ipin_in),
            .io_opin_out(io_tile_6_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .clk(clock),
            .reset(rst)
        );



    // FPGA LUT TILES DECLARE
    wire [839:0] lut_tile_1_1_chanxy_in;
    wire [199:0] lut_tile_1_1_chanxy_out;
    wire [527:0] lut_tile_1_1_ipin_in;
    wire [9:0] lut_tile_1_1_opin_out;
    lut_tile_sp_0 lut_tile_1_1(
            .io_chanxy_in(lut_tile_1_1_chanxy_in),
            .io_chanxy_out(lut_tile_1_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[55:7]),
            .io_ipin_in(lut_tile_1_1_ipin_in),
            .io_opin_out(lut_tile_1_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_2_1_chanxy_in;
    wire [139:0] lut_tile_2_1_chanxy_out;
    wire [527:0] lut_tile_2_1_ipin_in;
    wire [9:0] lut_tile_2_1_opin_out;
    lut_tile_sp_1 lut_tile_2_1(
            .io_chanxy_in(lut_tile_2_1_chanxy_in),
            .io_chanxy_out(lut_tile_2_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[102:56]),
            .io_ipin_in(lut_tile_2_1_ipin_in),
            .io_opin_out(lut_tile_2_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_3_1_chanxy_in;
    wire [139:0] lut_tile_3_1_chanxy_out;
    wire [527:0] lut_tile_3_1_ipin_in;
    wire [9:0] lut_tile_3_1_opin_out;
    lut_tile_sp_2 lut_tile_3_1(
            .io_chanxy_in(lut_tile_3_1_chanxy_in),
            .io_chanxy_out(lut_tile_3_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[149:103]),
            .io_ipin_in(lut_tile_3_1_ipin_in),
            .io_opin_out(lut_tile_3_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_4_1_chanxy_in;
    wire [139:0] lut_tile_4_1_chanxy_out;
    wire [527:0] lut_tile_4_1_ipin_in;
    wire [9:0] lut_tile_4_1_opin_out;
    lut_tile_sp_3 lut_tile_4_1(
            .io_chanxy_in(lut_tile_4_1_chanxy_in),
            .io_chanxy_out(lut_tile_4_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[196:150]),
            .io_ipin_in(lut_tile_4_1_ipin_in),
            .io_opin_out(lut_tile_4_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [759:0] lut_tile_5_1_chanxy_in;
    wire [199:0] lut_tile_5_1_chanxy_out;
    wire [527:0] lut_tile_5_1_ipin_in;
    wire [9:0] lut_tile_5_1_opin_out;
    lut_tile_sp_4 lut_tile_5_1(
            .io_chanxy_in(lut_tile_5_1_chanxy_in),
            .io_chanxy_out(lut_tile_5_1_chanxy_out),
            .io_configs_in(configs_in[63:32]),
            .io_configs_en(configs_en[243:197]),
            .io_ipin_in(lut_tile_5_1_ipin_in),
            .io_opin_out(lut_tile_5_1_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [775:0] lut_tile_1_5_chanxy_in;
    wire [199:0] lut_tile_1_5_chanxy_out;
    wire [527:0] lut_tile_1_5_ipin_in;
    wire [9:0] lut_tile_1_5_opin_out;
    lut_tile_sp_5 lut_tile_1_5(
            .io_chanxy_in(lut_tile_1_5_chanxy_in),
            .io_chanxy_out(lut_tile_1_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[54:7]),
            .io_ipin_in(lut_tile_1_5_ipin_in),
            .io_opin_out(lut_tile_1_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [795:0] lut_tile_2_5_chanxy_in;
    wire [139:0] lut_tile_2_5_chanxy_out;
    wire [527:0] lut_tile_2_5_ipin_in;
    wire [9:0] lut_tile_2_5_opin_out;
    lut_tile_sp_6 lut_tile_2_5(
            .io_chanxy_in(lut_tile_2_5_chanxy_in),
            .io_chanxy_out(lut_tile_2_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[102:56]),
            .io_ipin_in(lut_tile_2_5_ipin_in),
            .io_opin_out(lut_tile_2_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [795:0] lut_tile_3_5_chanxy_in;
    wire [139:0] lut_tile_3_5_chanxy_out;
    wire [527:0] lut_tile_3_5_ipin_in;
    wire [9:0] lut_tile_3_5_opin_out;
    lut_tile_sp_7 lut_tile_3_5(
            .io_chanxy_in(lut_tile_3_5_chanxy_in),
            .io_chanxy_out(lut_tile_3_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[149:103]),
            .io_ipin_in(lut_tile_3_5_ipin_in),
            .io_opin_out(lut_tile_3_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [795:0] lut_tile_4_5_chanxy_in;
    wire [139:0] lut_tile_4_5_chanxy_out;
    wire [527:0] lut_tile_4_5_ipin_in;
    wire [9:0] lut_tile_4_5_opin_out;
    lut_tile_sp_8 lut_tile_4_5(
            .io_chanxy_in(lut_tile_4_5_chanxy_in),
            .io_chanxy_out(lut_tile_4_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[196:150]),
            .io_ipin_in(lut_tile_4_5_ipin_in),
            .io_opin_out(lut_tile_4_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [695:0] lut_tile_5_5_chanxy_in;
    wire [199:0] lut_tile_5_5_chanxy_out;
    wire [527:0] lut_tile_5_5_ipin_in;
    wire [9:0] lut_tile_5_5_opin_out;
    lut_tile_sp_9 lut_tile_5_5(
            .io_chanxy_in(lut_tile_5_5_chanxy_in),
            .io_chanxy_out(lut_tile_5_5_chanxy_out),
            .io_configs_in(configs_in[191:160]),
            .io_configs_en(configs_en[242:197]),
            .io_ipin_in(lut_tile_5_5_ipin_in),
            .io_opin_out(lut_tile_5_5_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_1_2_chanxy_in;
    wire [139:0] lut_tile_1_2_chanxy_out;
    wire [527:0] lut_tile_1_2_ipin_in;
    wire [9:0] lut_tile_1_2_opin_out;
    lut_tile_sp_10 lut_tile_1_2(
            .io_chanxy_in(lut_tile_1_2_chanxy_in),
            .io_chanxy_out(lut_tile_1_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[53:7]),
            .io_ipin_in(lut_tile_1_2_ipin_in),
            .io_opin_out(lut_tile_1_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_1_3_chanxy_in;
    wire [139:0] lut_tile_1_3_chanxy_out;
    wire [527:0] lut_tile_1_3_ipin_in;
    wire [9:0] lut_tile_1_3_opin_out;
    lut_tile_sp_11 lut_tile_1_3(
            .io_chanxy_in(lut_tile_1_3_chanxy_in),
            .io_chanxy_out(lut_tile_1_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[53:7]),
            .io_ipin_in(lut_tile_1_3_ipin_in),
            .io_opin_out(lut_tile_1_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [859:0] lut_tile_1_4_chanxy_in;
    wire [139:0] lut_tile_1_4_chanxy_out;
    wire [527:0] lut_tile_1_4_ipin_in;
    wire [9:0] lut_tile_1_4_opin_out;
    lut_tile_sp_12 lut_tile_1_4(
            .io_chanxy_in(lut_tile_1_4_chanxy_in),
            .io_chanxy_out(lut_tile_1_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[53:7]),
            .io_ipin_in(lut_tile_1_4_ipin_in),
            .io_opin_out(lut_tile_1_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [779:0] lut_tile_5_2_chanxy_in;
    wire [139:0] lut_tile_5_2_chanxy_out;
    wire [527:0] lut_tile_5_2_ipin_in;
    wire [9:0] lut_tile_5_2_opin_out;
    lut_tile_sp_13 lut_tile_5_2(
            .io_chanxy_in(lut_tile_5_2_chanxy_in),
            .io_chanxy_out(lut_tile_5_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[243:197]),
            .io_ipin_in(lut_tile_5_2_ipin_in),
            .io_opin_out(lut_tile_5_2_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [779:0] lut_tile_5_3_chanxy_in;
    wire [139:0] lut_tile_5_3_chanxy_out;
    wire [527:0] lut_tile_5_3_ipin_in;
    wire [9:0] lut_tile_5_3_opin_out;
    lut_tile_sp_14 lut_tile_5_3(
            .io_chanxy_in(lut_tile_5_3_chanxy_in),
            .io_chanxy_out(lut_tile_5_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[243:197]),
            .io_ipin_in(lut_tile_5_3_ipin_in),
            .io_opin_out(lut_tile_5_3_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [779:0] lut_tile_5_4_chanxy_in;
    wire [139:0] lut_tile_5_4_chanxy_out;
    wire [527:0] lut_tile_5_4_ipin_in;
    wire [9:0] lut_tile_5_4_opin_out;
    lut_tile_sp_15 lut_tile_5_4(
            .io_chanxy_in(lut_tile_5_4_chanxy_in),
            .io_chanxy_out(lut_tile_5_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[243:197]),
            .io_ipin_in(lut_tile_5_4_ipin_in),
            .io_opin_out(lut_tile_5_4_opin_out),
            .io_x_loc(),
            .io_y_loc(),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_2_2_chanxy_in;
    wire [79:0] lut_tile_2_2_chanxy_out;
    wire [527:0] lut_tile_2_2_ipin_in;
    wire [9:0] lut_tile_2_2_opin_out;
    lut_tile lut_tile_2_2(
            .io_chanxy_in(lut_tile_2_2_chanxy_in),
            .io_chanxy_out(lut_tile_2_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[101:56]),
            .io_ipin_in(lut_tile_2_2_ipin_in),
            .io_opin_out(lut_tile_2_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_2_3_chanxy_in;
    wire [79:0] lut_tile_2_3_chanxy_out;
    wire [527:0] lut_tile_2_3_ipin_in;
    wire [9:0] lut_tile_2_3_opin_out;
    lut_tile lut_tile_2_3(
            .io_chanxy_in(lut_tile_2_3_chanxy_in),
            .io_chanxy_out(lut_tile_2_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[101:56]),
            .io_ipin_in(lut_tile_2_3_ipin_in),
            .io_opin_out(lut_tile_2_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_2_4_chanxy_in;
    wire [79:0] lut_tile_2_4_chanxy_out;
    wire [527:0] lut_tile_2_4_ipin_in;
    wire [9:0] lut_tile_2_4_opin_out;
    lut_tile lut_tile_2_4(
            .io_chanxy_in(lut_tile_2_4_chanxy_in),
            .io_chanxy_out(lut_tile_2_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[101:56]),
            .io_ipin_in(lut_tile_2_4_ipin_in),
            .io_opin_out(lut_tile_2_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_3_2_chanxy_in;
    wire [79:0] lut_tile_3_2_chanxy_out;
    wire [527:0] lut_tile_3_2_ipin_in;
    wire [9:0] lut_tile_3_2_opin_out;
    lut_tile lut_tile_3_2(
            .io_chanxy_in(lut_tile_3_2_chanxy_in),
            .io_chanxy_out(lut_tile_3_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[148:103]),
            .io_ipin_in(lut_tile_3_2_ipin_in),
            .io_opin_out(lut_tile_3_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_3_3_chanxy_in;
    wire [79:0] lut_tile_3_3_chanxy_out;
    wire [527:0] lut_tile_3_3_ipin_in;
    wire [9:0] lut_tile_3_3_opin_out;
    lut_tile lut_tile_3_3(
            .io_chanxy_in(lut_tile_3_3_chanxy_in),
            .io_chanxy_out(lut_tile_3_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[148:103]),
            .io_ipin_in(lut_tile_3_3_ipin_in),
            .io_opin_out(lut_tile_3_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_3_4_chanxy_in;
    wire [79:0] lut_tile_3_4_chanxy_out;
    wire [527:0] lut_tile_3_4_ipin_in;
    wire [9:0] lut_tile_3_4_opin_out;
    lut_tile lut_tile_3_4(
            .io_chanxy_in(lut_tile_3_4_chanxy_in),
            .io_chanxy_out(lut_tile_3_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[148:103]),
            .io_ipin_in(lut_tile_3_4_ipin_in),
            .io_opin_out(lut_tile_3_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_4_2_chanxy_in;
    wire [79:0] lut_tile_4_2_chanxy_out;
    wire [527:0] lut_tile_4_2_ipin_in;
    wire [9:0] lut_tile_4_2_opin_out;
    lut_tile lut_tile_4_2(
            .io_chanxy_in(lut_tile_4_2_chanxy_in),
            .io_chanxy_out(lut_tile_4_2_chanxy_out),
            .io_configs_in(configs_in[95:64]),
            .io_configs_en(configs_en[195:150]),
            .io_ipin_in(lut_tile_4_2_ipin_in),
            .io_opin_out(lut_tile_4_2_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_4_3_chanxy_in;
    wire [79:0] lut_tile_4_3_chanxy_out;
    wire [527:0] lut_tile_4_3_ipin_in;
    wire [9:0] lut_tile_4_3_opin_out;
    lut_tile lut_tile_4_3(
            .io_chanxy_in(lut_tile_4_3_chanxy_in),
            .io_chanxy_out(lut_tile_4_3_chanxy_out),
            .io_configs_in(configs_in[127:96]),
            .io_configs_en(configs_en[195:150]),
            .io_ipin_in(lut_tile_4_3_ipin_in),
            .io_opin_out(lut_tile_4_3_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );

    wire [879:0] lut_tile_4_4_chanxy_in;
    wire [79:0] lut_tile_4_4_chanxy_out;
    wire [527:0] lut_tile_4_4_ipin_in;
    wire [9:0] lut_tile_4_4_opin_out;
    lut_tile lut_tile_4_4(
            .io_chanxy_in(lut_tile_4_4_chanxy_in),
            .io_chanxy_out(lut_tile_4_4_chanxy_out),
            .io_configs_in(configs_in[159:128]),
            .io_configs_en(configs_en[195:150]),
            .io_ipin_in(lut_tile_4_4_ipin_in),
            .io_opin_out(lut_tile_4_4_opin_out),
            .io_ff_en(ff_en),
            .clk(clock),
            .reset(rst)
        );



    // LUT TILE IPIN
    assign lut_tile_1_1_ipin_in = {wire_2837, wire_2836, wire_2817, wire_2816, wire_2797, wire_2796, wire_2777, wire_2776, wire_2757, wire_2756, wire_2737, wire_2736, wire_2717, wire_2716, wire_2697, wire_2696, wire_4439, wire_4438, wire_4419, wire_4418, wire_4399, wire_4398, wire_4379, wire_4378, wire_4359, wire_4358, wire_4339, wire_4338, wire_4319, wire_4318, wire_4299, wire_4298, wire_2519, wire_2518, wire_2499, wire_2498, wire_2479, wire_2478, wire_2459, wire_2458, wire_2439, wire_2438, wire_2419, wire_2418, wire_2399, wire_2398, wire_2379, wire_2378, wire_4755, wire_4754, wire_4743, wire_4742, wire_4715, wire_4714, wire_4703, wire_4702, wire_4675, wire_4674, wire_4663, wire_4662, wire_4635, wire_4634, wire_4623, wire_4622, wire_2835, wire_2834, wire_2823, wire_2822, wire_2795, wire_2794, wire_2783, wire_2782, wire_2755, wire_2754, wire_2743, wire_2742, wire_2715, wire_2714, wire_2703, wire_2702, wire_4437, wire_4436, wire_4417, wire_4416, wire_4397, wire_4396, wire_4377, wire_4376, wire_4357, wire_4356, wire_4337, wire_4336, wire_4317, wire_4316, wire_4297, wire_4296, wire_2515, wire_2514, wire_2495, wire_2494, wire_2475, wire_2474, wire_2455, wire_2454, wire_2435, wire_2434, wire_2415, wire_2414, wire_2395, wire_2394, wire_2375, wire_2374, wire_4753, wire_4752, wire_4733, wire_4732, wire_4713, wire_4712, wire_4693, wire_4692, wire_4673, wire_4672, wire_4653, wire_4652, wire_4633, wire_4632, wire_4613, wire_4612, wire_2833, wire_2832, wire_2813, wire_2812, wire_2793, wire_2792, wire_2773, wire_2772, wire_2753, wire_2752, wire_2733, wire_2732, wire_2713, wire_2712, wire_2693, wire_2692, wire_4433, wire_4432, wire_4413, wire_4412, wire_4393, wire_4392, wire_4373, wire_4372, wire_4353, wire_4352, wire_4333, wire_4332, wire_4313, wire_4312, wire_4293, wire_4292, wire_2513, wire_2512, wire_2493, wire_2492, wire_2473, wire_2472, wire_2453, wire_2452, wire_2433, wire_2432, wire_2413, wire_2412, wire_2393, wire_2392, wire_2373, wire_2372, wire_4759, wire_4758, wire_4731, wire_4730, wire_4719, wire_4718, wire_4691, wire_4690, wire_4679, wire_4678, wire_4651, wire_4650, wire_4639, wire_4638, wire_4611, wire_4610, wire_2839, wire_2838, wire_2811, wire_2810, wire_2799, wire_2798, wire_2771, wire_2770, wire_2759, wire_2758, wire_2731, wire_2730, wire_2719, wire_2718, wire_2691, wire_2690, wire_4431, wire_4430, wire_4411, wire_4410, wire_4391, wire_4390, wire_4371, wire_4370, wire_4351, wire_4350, wire_4331, wire_4330, wire_4311, wire_4310, wire_4291, wire_4290, wire_2511, wire_2510, wire_2491, wire_2490, wire_2471, wire_2470, wire_2451, wire_2450, wire_2431, wire_2430, wire_2411, wire_2410, wire_2391, wire_2390, wire_2371, wire_2370, wire_4749, wire_4748, wire_4729, wire_4728, wire_4709, wire_4708, wire_4689, wire_4688, wire_4669, wire_4668, wire_4649, wire_4648, wire_4629, wire_4628, wire_4609, wire_4608, wire_2827, wire_2826, wire_2815, wire_2814, wire_2787, wire_2786, wire_2775, wire_2774, wire_2747, wire_2746, wire_2735, wire_2734, wire_2707, wire_2706, wire_2695, wire_2694, wire_4429, wire_4428, wire_4409, wire_4408, wire_4389, wire_4388, wire_4369, wire_4368, wire_4349, wire_4348, wire_4329, wire_4328, wire_4309, wire_4308, wire_4289, wire_4288, wire_2509, wire_2508, wire_2489, wire_2488, wire_2469, wire_2468, wire_2449, wire_2448, wire_2429, wire_2428, wire_2409, wire_2408, wire_2389, wire_2388, wire_2369, wire_2368, wire_4745, wire_4744, wire_4725, wire_4724, wire_4705, wire_4704, wire_4685, wire_4684, wire_4665, wire_4664, wire_4645, wire_4644, wire_4625, wire_4624, wire_4605, wire_4604, wire_2825, wire_2824, wire_2805, wire_2804, wire_2785, wire_2784, wire_2765, wire_2764, wire_2745, wire_2744, wire_2725, wire_2724, wire_2705, wire_2704, wire_2685, wire_2684, wire_4427, wire_4426, wire_4407, wire_4406, wire_4387, wire_4386, wire_4367, wire_4366, wire_4347, wire_4346, wire_4327, wire_4326, wire_4307, wire_4306, wire_4287, wire_4286, wire_2507, wire_2506, wire_2487, wire_2486, wire_2467, wire_2466, wire_2447, wire_2446, wire_2427, wire_2426, wire_2407, wire_2406, wire_2387, wire_2386, wire_2367, wire_2366, wire_4751, wire_4750, wire_4723, wire_4722, wire_4711, wire_4710, wire_4683, wire_4682, wire_4671, wire_4670, wire_4643, wire_4642, wire_4631, wire_4630, wire_4603, wire_4602, wire_2831, wire_2830, wire_2803, wire_2802, wire_2791, wire_2790, wire_2763, wire_2762, wire_2751, wire_2750, wire_2723, wire_2722, wire_2711, wire_2710, wire_2683, wire_2682, wire_4425, wire_4424, wire_4405, wire_4404, wire_4385, wire_4384, wire_4365, wire_4364, wire_4345, wire_4344, wire_4325, wire_4324, wire_4305, wire_4304, wire_4285, wire_4284, wire_2503, wire_2502, wire_2483, wire_2482, wire_2463, wire_2462, wire_2443, wire_2442, wire_2423, wire_2422, wire_2403, wire_2402, wire_2383, wire_2382, wire_2363, wire_2362, wire_4741, wire_4740, wire_4721, wire_4720, wire_4701, wire_4700, wire_4681, wire_4680, wire_4661, wire_4660, wire_4641, wire_4640, wire_4621, wire_4620, wire_4601, wire_4600, wire_2821, wire_2820, wire_2801, wire_2800, wire_2781, wire_2780, wire_2761, wire_2760, wire_2741, wire_2740, wire_2721, wire_2720, wire_2701, wire_2700, wire_2681, wire_2680, wire_4421, wire_4420, wire_4401, wire_4400, wire_4381, wire_4380, wire_4361, wire_4360, wire_4341, wire_4340, wire_4321, wire_4320, wire_4301, wire_4300, wire_4281, wire_4280, wire_2501, wire_2500, wire_2481, wire_2480, wire_2461, wire_2460, wire_2441, wire_2440, wire_2421, wire_2420, wire_2401, wire_2400, wire_2381, wire_2380, wire_2361, wire_2360, wire_4739, wire_4738, wire_4727, wire_4726, wire_4699, wire_4698, wire_4687, wire_4686, wire_4659, wire_4658, wire_4647, wire_4646, wire_4619, wire_4618, wire_4607, wire_4606, wire_2819, wire_2818, wire_2807, wire_2806, wire_2779, wire_2778, wire_2767, wire_2766, wire_2739, wire_2738, wire_2727, wire_2726, wire_2699, wire_2698, wire_2687, wire_2686};
    // IPIN TOTAL: 528
    assign lut_tile_2_1_ipin_in = {wire_3155, wire_3154, wire_3143, wire_3142, wire_3115, wire_3114, wire_3103, wire_3102, wire_3075, wire_3074, wire_3063, wire_3062, wire_3035, wire_3034, wire_3023, wire_3022, wire_4437, wire_4436, wire_4417, wire_4416, wire_4397, wire_4396, wire_4377, wire_4376, wire_4357, wire_4356, wire_4337, wire_4336, wire_4317, wire_4316, wire_4297, wire_4296, wire_2837, wire_2836, wire_2817, wire_2816, wire_2797, wire_2796, wire_2777, wire_2776, wire_2757, wire_2756, wire_2737, wire_2736, wire_2717, wire_2716, wire_2697, wire_2696, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_4753, wire_4752, wire_4713, wire_4712, wire_4673, wire_4672, wire_4633, wire_4632, wire_3153, wire_3152, wire_3141, wire_3140, wire_3113, wire_3112, wire_3101, wire_3100, wire_3073, wire_3072, wire_3061, wire_3060, wire_3033, wire_3032, wire_3021, wire_3020, wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_4423, wire_4422, wire_4383, wire_4382, wire_4343, wire_4342, wire_4303, wire_4302, wire_2833, wire_2832, wire_2813, wire_2812, wire_2793, wire_2792, wire_2773, wire_2772, wire_2753, wire_2752, wire_2733, wire_2732, wire_2713, wire_2712, wire_2693, wire_2692, wire_4759, wire_4758, wire_4731, wire_4730, wire_4719, wire_4718, wire_4691, wire_4690, wire_4679, wire_4678, wire_4651, wire_4650, wire_4639, wire_4638, wire_4611, wire_4610, wire_3159, wire_3158, wire_3131, wire_3130, wire_3119, wire_3118, wire_3091, wire_3090, wire_3079, wire_3078, wire_3051, wire_3050, wire_3039, wire_3038, wire_3011, wire_3010, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_4439, wire_4438, wire_4399, wire_4398, wire_4359, wire_4358, wire_4319, wire_4318, wire_2839, wire_2838, wire_2811, wire_2810, wire_2799, wire_2798, wire_2771, wire_2770, wire_2759, wire_2758, wire_2731, wire_2730, wire_2719, wire_2718, wire_2691, wire_2690, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_4729, wire_4728, wire_4689, wire_4688, wire_4649, wire_4648, wire_4609, wire_4608, wire_3157, wire_3156, wire_3129, wire_3128, wire_3117, wire_3116, wire_3089, wire_3088, wire_3077, wire_3076, wire_3049, wire_3048, wire_3037, wire_3036, wire_3009, wire_3008, wire_4429, wire_4428, wire_4409, wire_4408, wire_4389, wire_4388, wire_4369, wire_4368, wire_4349, wire_4348, wire_4329, wire_4328, wire_4309, wire_4308, wire_4289, wire_4288, wire_2829, wire_2828, wire_2809, wire_2808, wire_2789, wire_2788, wire_2769, wire_2768, wire_2749, wire_2748, wire_2729, wire_2728, wire_2709, wire_2708, wire_2689, wire_2688, wire_4747, wire_4746, wire_4735, wire_4734, wire_4707, wire_4706, wire_4695, wire_4694, wire_4667, wire_4666, wire_4655, wire_4654, wire_4627, wire_4626, wire_4615, wire_4614, wire_3145, wire_3144, wire_3133, wire_3132, wire_3105, wire_3104, wire_3093, wire_3092, wire_3065, wire_3064, wire_3053, wire_3052, wire_3025, wire_3024, wire_3013, wire_3012, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_4415, wire_4414, wire_4375, wire_4374, wire_4335, wire_4334, wire_4295, wire_4294, wire_2827, wire_2826, wire_2815, wire_2814, wire_2787, wire_2786, wire_2775, wire_2774, wire_2747, wire_2746, wire_2735, wire_2734, wire_2707, wire_2706, wire_2695, wire_2694, wire_4751, wire_4750, wire_4723, wire_4722, wire_4711, wire_4710, wire_4683, wire_4682, wire_4671, wire_4670, wire_4643, wire_4642, wire_4631, wire_4630, wire_4603, wire_4602, wire_3151, wire_3150, wire_3123, wire_3122, wire_3111, wire_3110, wire_3083, wire_3082, wire_3071, wire_3070, wire_3043, wire_3042, wire_3031, wire_3030, wire_3003, wire_3002, wire_4425, wire_4424, wire_4405, wire_4404, wire_4385, wire_4384, wire_4365, wire_4364, wire_4345, wire_4344, wire_4325, wire_4324, wire_4305, wire_4304, wire_4285, wire_4284, wire_2825, wire_2824, wire_2805, wire_2804, wire_2785, wire_2784, wire_2765, wire_2764, wire_2745, wire_2744, wire_2725, wire_2724, wire_2705, wire_2704, wire_2685, wire_2684, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_4721, wire_4720, wire_4681, wire_4680, wire_4641, wire_4640, wire_4601, wire_4600, wire_3149, wire_3148, wire_3121, wire_3120, wire_3109, wire_3108, wire_3081, wire_3080, wire_3069, wire_3068, wire_3041, wire_3040, wire_3029, wire_3028, wire_3001, wire_3000, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440, wire_4431, wire_4430, wire_4391, wire_4390, wire_4351, wire_4350, wire_4311, wire_4310, wire_2821, wire_2820, wire_2801, wire_2800, wire_2781, wire_2780, wire_2761, wire_2760, wire_2741, wire_2740, wire_2721, wire_2720, wire_2701, wire_2700, wire_2681, wire_2680, wire_4739, wire_4738, wire_4727, wire_4726, wire_4699, wire_4698, wire_4687, wire_4686, wire_4659, wire_4658, wire_4647, wire_4646, wire_4619, wire_4618, wire_4607, wire_4606, wire_3139, wire_3138, wire_3127, wire_3126, wire_3099, wire_3098, wire_3087, wire_3086, wire_3059, wire_3058, wire_3047, wire_3046, wire_3019, wire_3018, wire_3007, wire_3006, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_4407, wire_4406, wire_4367, wire_4366, wire_4327, wire_4326, wire_4287, wire_4286, wire_2819, wire_2818, wire_2807, wire_2806, wire_2779, wire_2778, wire_2767, wire_2766, wire_2739, wire_2738, wire_2727, wire_2726, wire_2699, wire_2698, wire_2687, wire_2686, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_4737, wire_4736, wire_4697, wire_4696, wire_4657, wire_4656, wire_4617, wire_4616, wire_3137, wire_3136, wire_3125, wire_3124, wire_3097, wire_3096, wire_3085, wire_3084, wire_3057, wire_3056, wire_3045, wire_3044, wire_3017, wire_3016, wire_3005, wire_3004};
    // IPIN TOTAL: 528
    assign lut_tile_3_1_ipin_in = {wire_3473, wire_3472, wire_3461, wire_3460, wire_3433, wire_3432, wire_3421, wire_3420, wire_3393, wire_3392, wire_3381, wire_3380, wire_3353, wire_3352, wire_3341, wire_3340, wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_4423, wire_4422, wire_4383, wire_4382, wire_4343, wire_4342, wire_4303, wire_4302, wire_3155, wire_3154, wire_3143, wire_3142, wire_3115, wire_3114, wire_3103, wire_3102, wire_3075, wire_3074, wire_3063, wire_3062, wire_3035, wire_3034, wire_3023, wire_3022, wire_4839, wire_4838, wire_4829, wire_4828, wire_4819, wire_4818, wire_4809, wire_4808, wire_4739, wire_4738, wire_4699, wire_4698, wire_4659, wire_4658, wire_4619, wire_4618, wire_3479, wire_3478, wire_3459, wire_3458, wire_3439, wire_3438, wire_3419, wire_3418, wire_3399, wire_3398, wire_3379, wire_3378, wire_3359, wire_3358, wire_3339, wire_3338, wire_4515, wire_4514, wire_4505, wire_4504, wire_4495, wire_4494, wire_4485, wire_4484, wire_4433, wire_4432, wire_4393, wire_4392, wire_4353, wire_4352, wire_4313, wire_4312, wire_3159, wire_3158, wire_3131, wire_3130, wire_3119, wire_3118, wire_3091, wire_3090, wire_3079, wire_3078, wire_3051, wire_3050, wire_3039, wire_3038, wire_3011, wire_3010, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_4729, wire_4728, wire_4689, wire_4688, wire_4649, wire_4648, wire_4609, wire_4608, wire_3477, wire_3476, wire_3449, wire_3448, wire_3437, wire_3436, wire_3409, wire_3408, wire_3397, wire_3396, wire_3369, wire_3368, wire_3357, wire_3356, wire_3329, wire_3328, wire_4519, wire_4518, wire_4509, wire_4508, wire_4499, wire_4498, wire_4489, wire_4488, wire_4409, wire_4408, wire_4369, wire_4368, wire_4329, wire_4328, wire_4289, wire_4288, wire_3157, wire_3156, wire_3129, wire_3128, wire_3117, wire_3116, wire_3089, wire_3088, wire_3077, wire_3076, wire_3049, wire_3048, wire_3037, wire_3036, wire_3009, wire_3008, wire_4833, wire_4832, wire_4823, wire_4822, wire_4813, wire_4812, wire_4803, wire_4802, wire_4755, wire_4754, wire_4715, wire_4714, wire_4675, wire_4674, wire_4635, wire_4634, wire_3475, wire_3474, wire_3455, wire_3454, wire_3435, wire_3434, wire_3415, wire_3414, wire_3395, wire_3394, wire_3375, wire_3374, wire_3355, wire_3354, wire_3335, wire_3334, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_4415, wire_4414, wire_4375, wire_4374, wire_4335, wire_4334, wire_4295, wire_4294, wire_3147, wire_3146, wire_3135, wire_3134, wire_3107, wire_3106, wire_3095, wire_3094, wire_3067, wire_3066, wire_3055, wire_3054, wire_3027, wire_3026, wire_3015, wire_3014, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_4745, wire_4744, wire_4705, wire_4704, wire_4665, wire_4664, wire_4625, wire_4624, wire_3471, wire_3470, wire_3451, wire_3450, wire_3431, wire_3430, wire_3411, wire_3410, wire_3391, wire_3390, wire_3371, wire_3370, wire_3351, wire_3350, wire_3331, wire_3330, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_4425, wire_4424, wire_4385, wire_4384, wire_4345, wire_4344, wire_4305, wire_4304, wire_3145, wire_3144, wire_3133, wire_3132, wire_3105, wire_3104, wire_3093, wire_3092, wire_3065, wire_3064, wire_3053, wire_3052, wire_3025, wire_3024, wire_3013, wire_3012, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_4721, wire_4720, wire_4681, wire_4680, wire_4641, wire_4640, wire_4601, wire_4600, wire_3469, wire_3468, wire_3441, wire_3440, wire_3429, wire_3428, wire_3401, wire_3400, wire_3389, wire_3388, wire_3361, wire_3360, wire_3349, wire_3348, wire_3321, wire_3320, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440, wire_4431, wire_4430, wire_4391, wire_4390, wire_4351, wire_4350, wire_4311, wire_4310, wire_3151, wire_3150, wire_3123, wire_3122, wire_3111, wire_3110, wire_3083, wire_3082, wire_3071, wire_3070, wire_3043, wire_3042, wire_3031, wire_3030, wire_3003, wire_3002, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_4747, wire_4746, wire_4707, wire_4706, wire_4667, wire_4666, wire_4627, wire_4626, wire_3467, wire_3466, wire_3447, wire_3446, wire_3427, wire_3426, wire_3407, wire_3406, wire_3387, wire_3386, wire_3367, wire_3366, wire_3347, wire_3346, wire_3327, wire_3326, wire_4517, wire_4516, wire_4507, wire_4506, wire_4497, wire_4496, wire_4487, wire_4486, wire_4401, wire_4400, wire_4361, wire_4360, wire_4321, wire_4320, wire_4281, wire_4280, wire_3139, wire_3138, wire_3127, wire_3126, wire_3099, wire_3098, wire_3087, wire_3086, wire_3059, wire_3058, wire_3047, wire_3046, wire_3019, wire_3018, wire_3007, wire_3006, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_4737, wire_4736, wire_4697, wire_4696, wire_4657, wire_4656, wire_4617, wire_4616, wire_3457, wire_3456, wire_3445, wire_3444, wire_3417, wire_3416, wire_3405, wire_3404, wire_3377, wire_3376, wire_3365, wire_3364, wire_3337, wire_3336, wire_3325, wire_3324, wire_4511, wire_4510, wire_4501, wire_4500, wire_4491, wire_4490, wire_4481, wire_4480, wire_4417, wire_4416, wire_4377, wire_4376, wire_4337, wire_4336, wire_4297, wire_4296, wire_3137, wire_3136, wire_3125, wire_3124, wire_3097, wire_3096, wire_3085, wire_3084, wire_3057, wire_3056, wire_3045, wire_3044, wire_3017, wire_3016, wire_3005, wire_3004, wire_4835, wire_4834, wire_4825, wire_4824, wire_4815, wire_4814, wire_4805, wire_4804, wire_4723, wire_4722, wire_4683, wire_4682, wire_4643, wire_4642, wire_4603, wire_4602, wire_3463, wire_3462, wire_3443, wire_3442, wire_3423, wire_3422, wire_3403, wire_3402, wire_3383, wire_3382, wire_3363, wire_3362, wire_3343, wire_3342, wire_3323, wire_3322};
    // IPIN TOTAL: 528
    assign lut_tile_4_1_ipin_in = {wire_3799, wire_3798, wire_3779, wire_3778, wire_3759, wire_3758, wire_3739, wire_3738, wire_3719, wire_3718, wire_3699, wire_3698, wire_3679, wire_3678, wire_3659, wire_3658, wire_4515, wire_4514, wire_4505, wire_4504, wire_4495, wire_4494, wire_4485, wire_4484, wire_4433, wire_4432, wire_4393, wire_4392, wire_4353, wire_4352, wire_4313, wire_4312, wire_3473, wire_3472, wire_3461, wire_3460, wire_3433, wire_3432, wire_3421, wire_3420, wire_3393, wire_3392, wire_3381, wire_3380, wire_3353, wire_3352, wire_3341, wire_3340, wire_4875, wire_4874, wire_4865, wire_4864, wire_4855, wire_4854, wire_4845, wire_4844, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_3797, wire_3796, wire_3777, wire_3776, wire_3757, wire_3756, wire_3737, wire_3736, wire_3717, wire_3716, wire_3697, wire_3696, wire_3677, wire_3676, wire_3657, wire_3656, wire_4559, wire_4558, wire_4549, wire_4548, wire_4539, wire_4538, wire_4529, wire_4528, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_3477, wire_3476, wire_3449, wire_3448, wire_3437, wire_3436, wire_3409, wire_3408, wire_3397, wire_3396, wire_3369, wire_3368, wire_3357, wire_3356, wire_3329, wire_3328, wire_4833, wire_4832, wire_4823, wire_4822, wire_4813, wire_4812, wire_4803, wire_4802, wire_4755, wire_4754, wire_4715, wire_4714, wire_4675, wire_4674, wire_4635, wire_4634, wire_3795, wire_3794, wire_3775, wire_3774, wire_3755, wire_3754, wire_3735, wire_3734, wire_3715, wire_3714, wire_3695, wire_3694, wire_3675, wire_3674, wire_3655, wire_3654, wire_4553, wire_4552, wire_4543, wire_4542, wire_4533, wire_4532, wire_4523, wire_4522, wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_3475, wire_3474, wire_3455, wire_3454, wire_3435, wire_3434, wire_3415, wire_3414, wire_3395, wire_3394, wire_3375, wire_3374, wire_3355, wire_3354, wire_3335, wire_3334, wire_4879, wire_4878, wire_4869, wire_4868, wire_4859, wire_4858, wire_4849, wire_4848, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_3793, wire_3792, wire_3773, wire_3772, wire_3753, wire_3752, wire_3733, wire_3732, wire_3713, wire_3712, wire_3693, wire_3692, wire_3673, wire_3672, wire_3653, wire_3652, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_4425, wire_4424, wire_4385, wire_4384, wire_4345, wire_4344, wire_4305, wire_4304, wire_3465, wire_3464, wire_3453, wire_3452, wire_3425, wire_3424, wire_3413, wire_3412, wire_3385, wire_3384, wire_3373, wire_3372, wire_3345, wire_3344, wire_3333, wire_3332, wire_4837, wire_4836, wire_4827, wire_4826, wire_4817, wire_4816, wire_4807, wire_4806, wire_4731, wire_4730, wire_4691, wire_4690, wire_4651, wire_4650, wire_4611, wire_4610, wire_3789, wire_3788, wire_3769, wire_3768, wire_3749, wire_3748, wire_3729, wire_3728, wire_3709, wire_3708, wire_3689, wire_3688, wire_3669, wire_3668, wire_3649, wire_3648, wire_4557, wire_4556, wire_4547, wire_4546, wire_4537, wire_4536, wire_4527, wire_4526, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_3471, wire_3470, wire_3451, wire_3450, wire_3431, wire_3430, wire_3411, wire_3410, wire_3391, wire_3390, wire_3371, wire_3370, wire_3351, wire_3350, wire_3331, wire_3330, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_4747, wire_4746, wire_4707, wire_4706, wire_4667, wire_4666, wire_4627, wire_4626, wire_3787, wire_3786, wire_3767, wire_3766, wire_3747, wire_3746, wire_3727, wire_3726, wire_3707, wire_3706, wire_3687, wire_3686, wire_3667, wire_3666, wire_3647, wire_3646, wire_4517, wire_4516, wire_4507, wire_4506, wire_4497, wire_4496, wire_4487, wire_4486, wire_4401, wire_4400, wire_4361, wire_4360, wire_4321, wire_4320, wire_4281, wire_4280, wire_3469, wire_3468, wire_3441, wire_3440, wire_3429, wire_3428, wire_3401, wire_3400, wire_3389, wire_3388, wire_3361, wire_3360, wire_3349, wire_3348, wire_3321, wire_3320, wire_4877, wire_4876, wire_4867, wire_4866, wire_4857, wire_4856, wire_4847, wire_4846, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_3785, wire_3784, wire_3765, wire_3764, wire_3745, wire_3744, wire_3725, wire_3724, wire_3705, wire_3704, wire_3685, wire_3684, wire_3665, wire_3664, wire_3645, wire_3644, wire_4551, wire_4550, wire_4541, wire_4540, wire_4531, wire_4530, wire_4521, wire_4520, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_3457, wire_3456, wire_3445, wire_3444, wire_3417, wire_3416, wire_3405, wire_3404, wire_3377, wire_3376, wire_3365, wire_3364, wire_3337, wire_3336, wire_3325, wire_3324, wire_4835, wire_4834, wire_4825, wire_4824, wire_4815, wire_4814, wire_4805, wire_4804, wire_4723, wire_4722, wire_4683, wire_4682, wire_4643, wire_4642, wire_4603, wire_4602, wire_3783, wire_3782, wire_3763, wire_3762, wire_3743, wire_3742, wire_3723, wire_3722, wire_3703, wire_3702, wire_3683, wire_3682, wire_3663, wire_3662, wire_3643, wire_3642, wire_4555, wire_4554, wire_4545, wire_4544, wire_4535, wire_4534, wire_4525, wire_4524, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440, wire_3463, wire_3462, wire_3443, wire_3442, wire_3423, wire_3422, wire_3403, wire_3402, wire_3383, wire_3382, wire_3363, wire_3362, wire_3343, wire_3342, wire_3323, wire_3322, wire_4871, wire_4870, wire_4861, wire_4860, wire_4851, wire_4850, wire_4841, wire_4840, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_3781, wire_3780, wire_3761, wire_3760, wire_3741, wire_3740, wire_3721, wire_3720, wire_3701, wire_3700, wire_3681, wire_3680, wire_3661, wire_3660, wire_3641, wire_3640};
    // IPIN TOTAL: 528
    assign lut_tile_5_1_ipin_in = {wire_4117, wire_4116, wire_4097, wire_4096, wire_4077, wire_4076, wire_4057, wire_4056, wire_4037, wire_4036, wire_4017, wire_4016, wire_3997, wire_3996, wire_3977, wire_3976, wire_4559, wire_4558, wire_4549, wire_4548, wire_4539, wire_4538, wire_4529, wire_4528, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_3799, wire_3798, wire_3779, wire_3778, wire_3759, wire_3758, wire_3739, wire_3738, wire_3719, wire_3718, wire_3699, wire_3698, wire_3679, wire_3678, wire_3659, wire_3658, wire_4919, wire_4918, wire_4909, wire_4908, wire_4899, wire_4898, wire_4889, wire_4888, wire_4835, wire_4834, wire_4825, wire_4824, wire_4815, wire_4814, wire_4805, wire_4804, wire_4115, wire_4114, wire_4103, wire_4102, wire_4075, wire_4074, wire_4063, wire_4062, wire_4035, wire_4034, wire_4023, wire_4022, wire_3995, wire_3994, wire_3983, wire_3982, wire_4595, wire_4594, wire_4585, wire_4584, wire_4575, wire_4574, wire_4565, wire_4564, wire_4519, wire_4518, wire_4509, wire_4508, wire_4499, wire_4498, wire_4489, wire_4488, wire_3795, wire_3794, wire_3775, wire_3774, wire_3755, wire_3754, wire_3735, wire_3734, wire_3715, wire_3714, wire_3695, wire_3694, wire_3675, wire_3674, wire_3655, wire_3654, wire_4879, wire_4878, wire_4869, wire_4868, wire_4859, wire_4858, wire_4849, wire_4848, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_4113, wire_4112, wire_4093, wire_4092, wire_4073, wire_4072, wire_4053, wire_4052, wire_4033, wire_4032, wire_4013, wire_4012, wire_3993, wire_3992, wire_3973, wire_3972, wire_4599, wire_4598, wire_4589, wire_4588, wire_4579, wire_4578, wire_4569, wire_4568, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_3793, wire_3792, wire_3773, wire_3772, wire_3753, wire_3752, wire_3733, wire_3732, wire_3713, wire_3712, wire_3693, wire_3692, wire_3673, wire_3672, wire_3653, wire_3652, wire_4913, wire_4912, wire_4903, wire_4902, wire_4893, wire_4892, wire_4883, wire_4882, wire_4839, wire_4838, wire_4829, wire_4828, wire_4819, wire_4818, wire_4809, wire_4808, wire_4119, wire_4118, wire_4091, wire_4090, wire_4079, wire_4078, wire_4051, wire_4050, wire_4039, wire_4038, wire_4011, wire_4010, wire_3999, wire_3998, wire_3971, wire_3970, wire_4557, wire_4556, wire_4547, wire_4546, wire_4537, wire_4536, wire_4527, wire_4526, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_3791, wire_3790, wire_3771, wire_3770, wire_3751, wire_3750, wire_3731, wire_3730, wire_3711, wire_3710, wire_3691, wire_3690, wire_3671, wire_3670, wire_3651, wire_3650, wire_4873, wire_4872, wire_4863, wire_4862, wire_4853, wire_4852, wire_4843, wire_4842, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_4107, wire_4106, wire_4095, wire_4094, wire_4067, wire_4066, wire_4055, wire_4054, wire_4027, wire_4026, wire_4015, wire_4014, wire_3987, wire_3986, wire_3975, wire_3974, wire_4593, wire_4592, wire_4583, wire_4582, wire_4573, wire_4572, wire_4563, wire_4562, wire_4517, wire_4516, wire_4507, wire_4506, wire_4497, wire_4496, wire_4487, wire_4486, wire_3789, wire_3788, wire_3769, wire_3768, wire_3749, wire_3748, wire_3729, wire_3728, wire_3709, wire_3708, wire_3689, wire_3688, wire_3669, wire_3668, wire_3649, wire_3648, wire_4877, wire_4876, wire_4867, wire_4866, wire_4857, wire_4856, wire_4847, wire_4846, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_4105, wire_4104, wire_4085, wire_4084, wire_4065, wire_4064, wire_4045, wire_4044, wire_4025, wire_4024, wire_4005, wire_4004, wire_3985, wire_3984, wire_3965, wire_3964, wire_4551, wire_4550, wire_4541, wire_4540, wire_4531, wire_4530, wire_4521, wire_4520, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_3787, wire_3786, wire_3767, wire_3766, wire_3747, wire_3746, wire_3727, wire_3726, wire_3707, wire_3706, wire_3687, wire_3686, wire_3667, wire_3666, wire_3647, wire_3646, wire_4911, wire_4910, wire_4901, wire_4900, wire_4891, wire_4890, wire_4881, wire_4880, wire_4837, wire_4836, wire_4827, wire_4826, wire_4817, wire_4816, wire_4807, wire_4806, wire_4111, wire_4110, wire_4083, wire_4082, wire_4071, wire_4070, wire_4043, wire_4042, wire_4031, wire_4030, wire_4003, wire_4002, wire_3991, wire_3990, wire_3963, wire_3962, wire_4597, wire_4596, wire_4587, wire_4586, wire_4577, wire_4576, wire_4567, wire_4566, wire_4511, wire_4510, wire_4501, wire_4500, wire_4491, wire_4490, wire_4481, wire_4480, wire_3783, wire_3782, wire_3763, wire_3762, wire_3743, wire_3742, wire_3723, wire_3722, wire_3703, wire_3702, wire_3683, wire_3682, wire_3663, wire_3662, wire_3643, wire_3642, wire_4871, wire_4870, wire_4861, wire_4860, wire_4851, wire_4850, wire_4841, wire_4840, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_4101, wire_4100, wire_4081, wire_4080, wire_4061, wire_4060, wire_4041, wire_4040, wire_4021, wire_4020, wire_4001, wire_4000, wire_3981, wire_3980, wire_3961, wire_3960, wire_4591, wire_4590, wire_4581, wire_4580, wire_4571, wire_4570, wire_4561, wire_4560, wire_4515, wire_4514, wire_4505, wire_4504, wire_4495, wire_4494, wire_4485, wire_4484, wire_3781, wire_3780, wire_3761, wire_3760, wire_3741, wire_3740, wire_3721, wire_3720, wire_3701, wire_3700, wire_3681, wire_3680, wire_3661, wire_3660, wire_3641, wire_3640, wire_4915, wire_4914, wire_4905, wire_4904, wire_4895, wire_4894, wire_4885, wire_4884, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_4099, wire_4098, wire_4087, wire_4086, wire_4059, wire_4058, wire_4047, wire_4046, wire_4019, wire_4018, wire_4007, wire_4006, wire_3979, wire_3978, wire_3967, wire_3966};
    // IPIN TOTAL: 528
    assign lut_tile_1_2_ipin_in = {wire_2835, wire_2834, wire_2823, wire_2822, wire_2795, wire_2794, wire_2783, wire_2782, wire_2755, wire_2754, wire_2743, wire_2742, wire_2715, wire_2714, wire_2703, wire_2702, wire_4757, wire_4756, wire_4737, wire_4736, wire_4717, wire_4716, wire_4697, wire_4696, wire_4677, wire_4676, wire_4657, wire_4656, wire_4637, wire_4636, wire_4617, wire_4616, wire_2517, wire_2516, wire_2497, wire_2496, wire_2477, wire_2476, wire_2457, wire_2456, wire_2437, wire_2436, wire_2417, wire_2416, wire_2397, wire_2396, wire_2377, wire_2376, wire_5073, wire_5072, wire_5061, wire_5060, wire_5033, wire_5032, wire_5021, wire_5020, wire_4993, wire_4992, wire_4981, wire_4980, wire_4953, wire_4952, wire_4941, wire_4940, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_2833, wire_2832, wire_2793, wire_2792, wire_2753, wire_2752, wire_2713, wire_2712, wire_4755, wire_4754, wire_4743, wire_4742, wire_4715, wire_4714, wire_4703, wire_4702, wire_4675, wire_4674, wire_4663, wire_4662, wire_4635, wire_4634, wire_4623, wire_4622, wire_2513, wire_2512, wire_2493, wire_2492, wire_2473, wire_2472, wire_2453, wire_2452, wire_2433, wire_2432, wire_2413, wire_2412, wire_2393, wire_2392, wire_2373, wire_2372, wire_5079, wire_5078, wire_5051, wire_5050, wire_5039, wire_5038, wire_5011, wire_5010, wire_4999, wire_4998, wire_4971, wire_4970, wire_4959, wire_4958, wire_4931, wire_4930, wire_2839, wire_2838, wire_2811, wire_2810, wire_2799, wire_2798, wire_2771, wire_2770, wire_2759, wire_2758, wire_2731, wire_2730, wire_2719, wire_2718, wire_2691, wire_2690, wire_4759, wire_4758, wire_4731, wire_4730, wire_4719, wire_4718, wire_4691, wire_4690, wire_4679, wire_4678, wire_4651, wire_4650, wire_4639, wire_4638, wire_4611, wire_4610, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_2519, wire_2518, wire_2479, wire_2478, wire_2439, wire_2438, wire_2399, wire_2398, wire_5077, wire_5076, wire_5049, wire_5048, wire_5037, wire_5036, wire_5009, wire_5008, wire_4997, wire_4996, wire_4969, wire_4968, wire_4957, wire_4956, wire_4929, wire_4928, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_2809, wire_2808, wire_2769, wire_2768, wire_2729, wire_2728, wire_2689, wire_2688, wire_4749, wire_4748, wire_4729, wire_4728, wire_4709, wire_4708, wire_4689, wire_4688, wire_4669, wire_4668, wire_4649, wire_4648, wire_4629, wire_4628, wire_4609, wire_4608, wire_2509, wire_2508, wire_2489, wire_2488, wire_2469, wire_2468, wire_2449, wire_2448, wire_2429, wire_2428, wire_2409, wire_2408, wire_2389, wire_2388, wire_2369, wire_2368, wire_5067, wire_5066, wire_5055, wire_5054, wire_5027, wire_5026, wire_5015, wire_5014, wire_4987, wire_4986, wire_4975, wire_4974, wire_4947, wire_4946, wire_4935, wire_4934, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_2825, wire_2824, wire_2785, wire_2784, wire_2745, wire_2744, wire_2705, wire_2704, wire_4747, wire_4746, wire_4735, wire_4734, wire_4707, wire_4706, wire_4695, wire_4694, wire_4667, wire_4666, wire_4655, wire_4654, wire_4627, wire_4626, wire_4615, wire_4614, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_2495, wire_2494, wire_2455, wire_2454, wire_2415, wire_2414, wire_2375, wire_2374, wire_5071, wire_5070, wire_5043, wire_5042, wire_5031, wire_5030, wire_5003, wire_5002, wire_4991, wire_4990, wire_4963, wire_4962, wire_4951, wire_4950, wire_4923, wire_4922, wire_2831, wire_2830, wire_2803, wire_2802, wire_2791, wire_2790, wire_2763, wire_2762, wire_2751, wire_2750, wire_2723, wire_2722, wire_2711, wire_2710, wire_2683, wire_2682, wire_4745, wire_4744, wire_4725, wire_4724, wire_4705, wire_4704, wire_4685, wire_4684, wire_4665, wire_4664, wire_4645, wire_4644, wire_4625, wire_4624, wire_4605, wire_4604, wire_2505, wire_2504, wire_2485, wire_2484, wire_2465, wire_2464, wire_2445, wire_2444, wire_2425, wire_2424, wire_2405, wire_2404, wire_2385, wire_2384, wire_2365, wire_2364, wire_5069, wire_5068, wire_5041, wire_5040, wire_5029, wire_5028, wire_5001, wire_5000, wire_4989, wire_4988, wire_4961, wire_4960, wire_4949, wire_4948, wire_4921, wire_4920, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_2801, wire_2800, wire_2761, wire_2760, wire_2721, wire_2720, wire_2681, wire_2680, wire_4751, wire_4750, wire_4723, wire_4722, wire_4711, wire_4710, wire_4683, wire_4682, wire_4671, wire_4670, wire_4643, wire_4642, wire_4631, wire_4630, wire_4603, wire_4602, wire_2501, wire_2500, wire_2481, wire_2480, wire_2461, wire_2460, wire_2441, wire_2440, wire_2421, wire_2420, wire_2401, wire_2400, wire_2381, wire_2380, wire_2361, wire_2360, wire_5059, wire_5058, wire_5047, wire_5046, wire_5019, wire_5018, wire_5007, wire_5006, wire_4979, wire_4978, wire_4967, wire_4966, wire_4939, wire_4938, wire_4927, wire_4926, wire_2819, wire_2818, wire_2807, wire_2806, wire_2779, wire_2778, wire_2767, wire_2766, wire_2739, wire_2738, wire_2727, wire_2726, wire_2699, wire_2698, wire_2687, wire_2686, wire_4739, wire_4738, wire_4727, wire_4726, wire_4699, wire_4698, wire_4687, wire_4686, wire_4659, wire_4658, wire_4647, wire_4646, wire_4619, wire_4618, wire_4607, wire_4606, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_2487, wire_2486, wire_2447, wire_2446, wire_2407, wire_2406, wire_2367, wire_2366, wire_5057, wire_5056, wire_5045, wire_5044, wire_5017, wire_5016, wire_5005, wire_5004, wire_4977, wire_4976, wire_4965, wire_4964, wire_4937, wire_4936, wire_4925, wire_4924, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_2817, wire_2816, wire_2777, wire_2776, wire_2737, wire_2736, wire_2697, wire_2696};
    // IPIN TOTAL: 528
    assign lut_tile_2_2_ipin_in = {wire_3153, wire_3152, wire_3141, wire_3140, wire_3113, wire_3112, wire_3101, wire_3100, wire_3073, wire_3072, wire_3061, wire_3060, wire_3033, wire_3032, wire_3021, wire_3020, wire_4755, wire_4754, wire_4743, wire_4742, wire_4715, wire_4714, wire_4703, wire_4702, wire_4675, wire_4674, wire_4663, wire_4662, wire_4635, wire_4634, wire_4623, wire_4622, wire_2835, wire_2834, wire_2823, wire_2822, wire_2795, wire_2794, wire_2783, wire_2782, wire_2755, wire_2754, wire_2743, wire_2742, wire_2715, wire_2714, wire_2703, wire_2702, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_5059, wire_5058, wire_5019, wire_5018, wire_4979, wire_4978, wire_4939, wire_4938, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_3139, wire_3138, wire_3099, wire_3098, wire_3059, wire_3058, wire_3019, wire_3018, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_4753, wire_4752, wire_4713, wire_4712, wire_4673, wire_4672, wire_4633, wire_4632, wire_2839, wire_2838, wire_2811, wire_2810, wire_2799, wire_2798, wire_2771, wire_2770, wire_2759, wire_2758, wire_2731, wire_2730, wire_2719, wire_2718, wire_2691, wire_2690, wire_5077, wire_5076, wire_5049, wire_5048, wire_5037, wire_5036, wire_5009, wire_5008, wire_4997, wire_4996, wire_4969, wire_4968, wire_4957, wire_4956, wire_4929, wire_4928, wire_3157, wire_3156, wire_3129, wire_3128, wire_3117, wire_3116, wire_3089, wire_3088, wire_3077, wire_3076, wire_3049, wire_3048, wire_3037, wire_3036, wire_3009, wire_3008, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_4729, wire_4728, wire_4689, wire_4688, wire_4649, wire_4648, wire_4609, wire_4608, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_2809, wire_2808, wire_2769, wire_2768, wire_2729, wire_2728, wire_2689, wire_2688, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_5075, wire_5074, wire_5035, wire_5034, wire_4995, wire_4994, wire_4955, wire_4954, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_3155, wire_3154, wire_3115, wire_3114, wire_3075, wire_3074, wire_3035, wire_3034, wire_4747, wire_4746, wire_4735, wire_4734, wire_4707, wire_4706, wire_4695, wire_4694, wire_4667, wire_4666, wire_4655, wire_4654, wire_4627, wire_4626, wire_4615, wire_4614, wire_2827, wire_2826, wire_2815, wire_2814, wire_2787, wire_2786, wire_2775, wire_2774, wire_2747, wire_2746, wire_2735, wire_2734, wire_2707, wire_2706, wire_2695, wire_2694, wire_5065, wire_5064, wire_5053, wire_5052, wire_5025, wire_5024, wire_5013, wire_5012, wire_4985, wire_4984, wire_4973, wire_4972, wire_4945, wire_4944, wire_4933, wire_4932, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_3131, wire_3130, wire_3091, wire_3090, wire_3051, wire_3050, wire_3011, wire_3010, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_4745, wire_4744, wire_4705, wire_4704, wire_4665, wire_4664, wire_4625, wire_4624, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_2825, wire_2824, wire_2785, wire_2784, wire_2745, wire_2744, wire_2705, wire_2704, wire_5069, wire_5068, wire_5041, wire_5040, wire_5029, wire_5028, wire_5001, wire_5000, wire_4989, wire_4988, wire_4961, wire_4960, wire_4949, wire_4948, wire_4921, wire_4920, wire_3149, wire_3148, wire_3121, wire_3120, wire_3109, wire_3108, wire_3081, wire_3080, wire_3069, wire_3068, wire_3041, wire_3040, wire_3029, wire_3028, wire_3001, wire_3000, wire_4751, wire_4750, wire_4723, wire_4722, wire_4711, wire_4710, wire_4683, wire_4682, wire_4671, wire_4670, wire_4643, wire_4642, wire_4631, wire_4630, wire_4603, wire_4602, wire_2831, wire_2830, wire_2803, wire_2802, wire_2791, wire_2790, wire_2763, wire_2762, wire_2751, wire_2750, wire_2723, wire_2722, wire_2711, wire_2710, wire_2683, wire_2682, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_5067, wire_5066, wire_5027, wire_5026, wire_4987, wire_4986, wire_4947, wire_4946, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_3147, wire_3146, wire_3107, wire_3106, wire_3067, wire_3066, wire_3027, wire_3026, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_4721, wire_4720, wire_4681, wire_4680, wire_4641, wire_4640, wire_4601, wire_4600, wire_2819, wire_2818, wire_2807, wire_2806, wire_2779, wire_2778, wire_2767, wire_2766, wire_2739, wire_2738, wire_2727, wire_2726, wire_2699, wire_2698, wire_2687, wire_2686, wire_5057, wire_5056, wire_5045, wire_5044, wire_5017, wire_5016, wire_5005, wire_5004, wire_4977, wire_4976, wire_4965, wire_4964, wire_4937, wire_4936, wire_4925, wire_4924, wire_3137, wire_3136, wire_3125, wire_3124, wire_3097, wire_3096, wire_3085, wire_3084, wire_3057, wire_3056, wire_3045, wire_3044, wire_3017, wire_3016, wire_3005, wire_3004, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_4737, wire_4736, wire_4697, wire_4696, wire_4657, wire_4656, wire_4617, wire_4616, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_2817, wire_2816, wire_2777, wire_2776, wire_2737, wire_2736, wire_2697, wire_2696, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_5043, wire_5042, wire_5003, wire_5002, wire_4963, wire_4962, wire_4923, wire_4922, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_3123, wire_3122, wire_3083, wire_3082, wire_3043, wire_3042, wire_3003, wire_3002};
    // IPIN TOTAL: 528
    assign lut_tile_3_2_ipin_in = {wire_3479, wire_3478, wire_3459, wire_3458, wire_3439, wire_3438, wire_3419, wire_3418, wire_3399, wire_3398, wire_3379, wire_3378, wire_3359, wire_3358, wire_3339, wire_3338, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_4753, wire_4752, wire_4713, wire_4712, wire_4673, wire_4672, wire_4633, wire_4632, wire_3153, wire_3152, wire_3141, wire_3140, wire_3113, wire_3112, wire_3101, wire_3100, wire_3073, wire_3072, wire_3061, wire_3060, wire_3033, wire_3032, wire_3021, wire_3020, wire_5155, wire_5154, wire_5145, wire_5144, wire_5135, wire_5134, wire_5125, wire_5124, wire_5077, wire_5076, wire_5037, wire_5036, wire_4997, wire_4996, wire_4957, wire_4956, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_3477, wire_3476, wire_3437, wire_3436, wire_3397, wire_3396, wire_3357, wire_3356, wire_4839, wire_4838, wire_4829, wire_4828, wire_4819, wire_4818, wire_4809, wire_4808, wire_4739, wire_4738, wire_4699, wire_4698, wire_4659, wire_4658, wire_4619, wire_4618, wire_3157, wire_3156, wire_3129, wire_3128, wire_3117, wire_3116, wire_3089, wire_3088, wire_3077, wire_3076, wire_3049, wire_3048, wire_3037, wire_3036, wire_3009, wire_3008, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_5075, wire_5074, wire_5035, wire_5034, wire_4995, wire_4994, wire_4955, wire_4954, wire_3475, wire_3474, wire_3455, wire_3454, wire_3435, wire_3434, wire_3415, wire_3414, wire_3395, wire_3394, wire_3375, wire_3374, wire_3355, wire_3354, wire_3335, wire_3334, wire_4833, wire_4832, wire_4823, wire_4822, wire_4813, wire_4812, wire_4803, wire_4802, wire_4755, wire_4754, wire_4715, wire_4714, wire_4675, wire_4674, wire_4635, wire_4634, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_3155, wire_3154, wire_3115, wire_3114, wire_3075, wire_3074, wire_3035, wire_3034, wire_5159, wire_5158, wire_5149, wire_5148, wire_5139, wire_5138, wire_5129, wire_5128, wire_5053, wire_5052, wire_5013, wire_5012, wire_4973, wire_4972, wire_4933, wire_4932, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_3453, wire_3452, wire_3413, wire_3412, wire_3373, wire_3372, wire_3333, wire_3332, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_4745, wire_4744, wire_4705, wire_4704, wire_4665, wire_4664, wire_4625, wire_4624, wire_3145, wire_3144, wire_3133, wire_3132, wire_3105, wire_3104, wire_3093, wire_3092, wire_3065, wire_3064, wire_3053, wire_3052, wire_3025, wire_3024, wire_3013, wire_3012, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_5051, wire_5050, wire_5011, wire_5010, wire_4971, wire_4970, wire_4931, wire_4930, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_3469, wire_3468, wire_3429, wire_3428, wire_3389, wire_3388, wire_3349, wire_3348, wire_4837, wire_4836, wire_4827, wire_4826, wire_4817, wire_4816, wire_4807, wire_4806, wire_4731, wire_4730, wire_4691, wire_4690, wire_4651, wire_4650, wire_4611, wire_4610, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_3131, wire_3130, wire_3091, wire_3090, wire_3051, wire_3050, wire_3011, wire_3010, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_5067, wire_5066, wire_5027, wire_5026, wire_4987, wire_4986, wire_4947, wire_4946, wire_3467, wire_3466, wire_3447, wire_3446, wire_3427, wire_3426, wire_3407, wire_3406, wire_3387, wire_3386, wire_3367, wire_3366, wire_3347, wire_3346, wire_3327, wire_3326, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_4721, wire_4720, wire_4681, wire_4680, wire_4641, wire_4640, wire_4601, wire_4600, wire_3149, wire_3148, wire_3121, wire_3120, wire_3109, wire_3108, wire_3081, wire_3080, wire_3069, wire_3068, wire_3041, wire_3040, wire_3029, wire_3028, wire_3001, wire_3000, wire_5157, wire_5156, wire_5147, wire_5146, wire_5137, wire_5136, wire_5127, wire_5126, wire_5045, wire_5044, wire_5005, wire_5004, wire_4965, wire_4964, wire_4925, wire_4924, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_3445, wire_3444, wire_3405, wire_3404, wire_3365, wire_3364, wire_3325, wire_3324, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_4747, wire_4746, wire_4707, wire_4706, wire_4667, wire_4666, wire_4627, wire_4626, wire_3137, wire_3136, wire_3125, wire_3124, wire_3097, wire_3096, wire_3085, wire_3084, wire_3057, wire_3056, wire_3045, wire_3044, wire_3017, wire_3016, wire_3005, wire_3004, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_5043, wire_5042, wire_5003, wire_5002, wire_4963, wire_4962, wire_4923, wire_4922, wire_3463, wire_3462, wire_3443, wire_3442, wire_3423, wire_3422, wire_3403, wire_3402, wire_3383, wire_3382, wire_3363, wire_3362, wire_3343, wire_3342, wire_3323, wire_3322, wire_4835, wire_4834, wire_4825, wire_4824, wire_4815, wire_4814, wire_4805, wire_4804, wire_4723, wire_4722, wire_4683, wire_4682, wire_4643, wire_4642, wire_4603, wire_4602, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_3123, wire_3122, wire_3083, wire_3082, wire_3043, wire_3042, wire_3003, wire_3002, wire_5151, wire_5150, wire_5141, wire_5140, wire_5131, wire_5130, wire_5121, wire_5120, wire_5061, wire_5060, wire_5021, wire_5020, wire_4981, wire_4980, wire_4941, wire_4940, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_3461, wire_3460, wire_3421, wire_3420, wire_3381, wire_3380, wire_3341, wire_3340};
    // IPIN TOTAL: 528
    assign lut_tile_4_2_ipin_in = {wire_3797, wire_3796, wire_3777, wire_3776, wire_3757, wire_3756, wire_3737, wire_3736, wire_3717, wire_3716, wire_3697, wire_3696, wire_3677, wire_3676, wire_3657, wire_3656, wire_4839, wire_4838, wire_4829, wire_4828, wire_4819, wire_4818, wire_4809, wire_4808, wire_4739, wire_4738, wire_4699, wire_4698, wire_4659, wire_4658, wire_4619, wire_4618, wire_3479, wire_3478, wire_3459, wire_3458, wire_3439, wire_3438, wire_3419, wire_3418, wire_3399, wire_3398, wire_3379, wire_3378, wire_3359, wire_3358, wire_3339, wire_3338, wire_5199, wire_5198, wire_5189, wire_5188, wire_5179, wire_5178, wire_5169, wire_5168, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_3783, wire_3782, wire_3743, wire_3742, wire_3703, wire_3702, wire_3663, wire_3662, wire_4875, wire_4874, wire_4865, wire_4864, wire_4855, wire_4854, wire_4845, wire_4844, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_3475, wire_3474, wire_3455, wire_3454, wire_3435, wire_3434, wire_3415, wire_3414, wire_3395, wire_3394, wire_3375, wire_3374, wire_3355, wire_3354, wire_3335, wire_3334, wire_5159, wire_5158, wire_5149, wire_5148, wire_5139, wire_5138, wire_5129, wire_5128, wire_5053, wire_5052, wire_5013, wire_5012, wire_4973, wire_4972, wire_4933, wire_4932, wire_3793, wire_3792, wire_3773, wire_3772, wire_3753, wire_3752, wire_3733, wire_3732, wire_3713, wire_3712, wire_3693, wire_3692, wire_3673, wire_3672, wire_3653, wire_3652, wire_4879, wire_4878, wire_4869, wire_4868, wire_4859, wire_4858, wire_4849, wire_4848, wire_4793, wire_4792, wire_4783, wire_4782, wire_4773, wire_4772, wire_4763, wire_4762, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_3453, wire_3452, wire_3413, wire_3412, wire_3373, wire_3372, wire_3333, wire_3332, wire_5193, wire_5192, wire_5183, wire_5182, wire_5173, wire_5172, wire_5163, wire_5162, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_3799, wire_3798, wire_3759, wire_3758, wire_3719, wire_3718, wire_3679, wire_3678, wire_4837, wire_4836, wire_4827, wire_4826, wire_4817, wire_4816, wire_4807, wire_4806, wire_4731, wire_4730, wire_4691, wire_4690, wire_4651, wire_4650, wire_4611, wire_4610, wire_3471, wire_3470, wire_3451, wire_3450, wire_3431, wire_3430, wire_3411, wire_3410, wire_3391, wire_3390, wire_3371, wire_3370, wire_3351, wire_3350, wire_3331, wire_3330, wire_5153, wire_5152, wire_5143, wire_5142, wire_5133, wire_5132, wire_5123, wire_5122, wire_5069, wire_5068, wire_5029, wire_5028, wire_4989, wire_4988, wire_4949, wire_4948, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_3775, wire_3774, wire_3735, wire_3734, wire_3695, wire_3694, wire_3655, wire_3654, wire_4873, wire_4872, wire_4863, wire_4862, wire_4853, wire_4852, wire_4843, wire_4842, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_3469, wire_3468, wire_3429, wire_3428, wire_3389, wire_3388, wire_3349, wire_3348, wire_5157, wire_5156, wire_5147, wire_5146, wire_5137, wire_5136, wire_5127, wire_5126, wire_5045, wire_5044, wire_5005, wire_5004, wire_4965, wire_4964, wire_4925, wire_4924, wire_3785, wire_3784, wire_3765, wire_3764, wire_3745, wire_3744, wire_3725, wire_3724, wire_3705, wire_3704, wire_3685, wire_3684, wire_3665, wire_3664, wire_3645, wire_3644, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_4747, wire_4746, wire_4707, wire_4706, wire_4667, wire_4666, wire_4627, wire_4626, wire_3467, wire_3466, wire_3447, wire_3446, wire_3427, wire_3426, wire_3407, wire_3406, wire_3387, wire_3386, wire_3367, wire_3366, wire_3347, wire_3346, wire_3327, wire_3326, wire_5191, wire_5190, wire_5181, wire_5180, wire_5171, wire_5170, wire_5161, wire_5160, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_3791, wire_3790, wire_3751, wire_3750, wire_3711, wire_3710, wire_3671, wire_3670, wire_4877, wire_4876, wire_4867, wire_4866, wire_4857, wire_4856, wire_4847, wire_4846, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_3463, wire_3462, wire_3443, wire_3442, wire_3423, wire_3422, wire_3403, wire_3402, wire_3383, wire_3382, wire_3363, wire_3362, wire_3343, wire_3342, wire_3323, wire_3322, wire_5151, wire_5150, wire_5141, wire_5140, wire_5131, wire_5130, wire_5121, wire_5120, wire_5061, wire_5060, wire_5021, wire_5020, wire_4981, wire_4980, wire_4941, wire_4940, wire_3781, wire_3780, wire_3761, wire_3760, wire_3741, wire_3740, wire_3721, wire_3720, wire_3701, wire_3700, wire_3681, wire_3680, wire_3661, wire_3660, wire_3641, wire_3640, wire_4871, wire_4870, wire_4861, wire_4860, wire_4851, wire_4850, wire_4841, wire_4840, wire_4795, wire_4794, wire_4785, wire_4784, wire_4775, wire_4774, wire_4765, wire_4764, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_3461, wire_3460, wire_3421, wire_3420, wire_3381, wire_3380, wire_3341, wire_3340, wire_5195, wire_5194, wire_5185, wire_5184, wire_5175, wire_5174, wire_5165, wire_5164, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_3767, wire_3766, wire_3727, wire_3726, wire_3687, wire_3686, wire_3647, wire_3646};
    // IPIN TOTAL: 528
    assign lut_tile_5_2_ipin_in = {wire_4115, wire_4114, wire_4103, wire_4102, wire_4075, wire_4074, wire_4063, wire_4062, wire_4035, wire_4034, wire_4023, wire_4022, wire_3995, wire_3994, wire_3983, wire_3982, wire_4875, wire_4874, wire_4865, wire_4864, wire_4855, wire_4854, wire_4845, wire_4844, wire_4799, wire_4798, wire_4789, wire_4788, wire_4779, wire_4778, wire_4769, wire_4768, wire_3797, wire_3796, wire_3777, wire_3776, wire_3757, wire_3756, wire_3737, wire_3736, wire_3717, wire_3716, wire_3697, wire_3696, wire_3677, wire_3676, wire_3657, wire_3656, wire_5235, wire_5234, wire_5225, wire_5224, wire_5215, wire_5214, wire_5205, wire_5204, wire_5159, wire_5158, wire_5149, wire_5148, wire_5139, wire_5138, wire_5129, wire_5128, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_4113, wire_4112, wire_4073, wire_4072, wire_4033, wire_4032, wire_3993, wire_3992, wire_4919, wire_4918, wire_4909, wire_4908, wire_4899, wire_4898, wire_4889, wire_4888, wire_4835, wire_4834, wire_4825, wire_4824, wire_4815, wire_4814, wire_4805, wire_4804, wire_3793, wire_3792, wire_3773, wire_3772, wire_3753, wire_3752, wire_3733, wire_3732, wire_3713, wire_3712, wire_3693, wire_3692, wire_3673, wire_3672, wire_3653, wire_3652, wire_5193, wire_5192, wire_5183, wire_5182, wire_5173, wire_5172, wire_5163, wire_5162, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_4119, wire_4118, wire_4091, wire_4090, wire_4079, wire_4078, wire_4051, wire_4050, wire_4039, wire_4038, wire_4011, wire_4010, wire_3999, wire_3998, wire_3971, wire_3970, wire_4913, wire_4912, wire_4903, wire_4902, wire_4893, wire_4892, wire_4883, wire_4882, wire_4839, wire_4838, wire_4829, wire_4828, wire_4819, wire_4818, wire_4809, wire_4808, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_3799, wire_3798, wire_3759, wire_3758, wire_3719, wire_3718, wire_3679, wire_3678, wire_5239, wire_5238, wire_5229, wire_5228, wire_5219, wire_5218, wire_5209, wire_5208, wire_5153, wire_5152, wire_5143, wire_5142, wire_5133, wire_5132, wire_5123, wire_5122, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_4089, wire_4088, wire_4049, wire_4048, wire_4009, wire_4008, wire_3969, wire_3968, wire_4873, wire_4872, wire_4863, wire_4862, wire_4853, wire_4852, wire_4843, wire_4842, wire_4797, wire_4796, wire_4787, wire_4786, wire_4777, wire_4776, wire_4767, wire_4766, wire_3789, wire_3788, wire_3769, wire_3768, wire_3749, wire_3748, wire_3729, wire_3728, wire_3709, wire_3708, wire_3689, wire_3688, wire_3669, wire_3668, wire_3649, wire_3648, wire_5197, wire_5196, wire_5187, wire_5186, wire_5177, wire_5176, wire_5167, wire_5166, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_4105, wire_4104, wire_4065, wire_4064, wire_4025, wire_4024, wire_3985, wire_3984, wire_4917, wire_4916, wire_4907, wire_4906, wire_4897, wire_4896, wire_4887, wire_4886, wire_4833, wire_4832, wire_4823, wire_4822, wire_4813, wire_4812, wire_4803, wire_4802, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_3775, wire_3774, wire_3735, wire_3734, wire_3695, wire_3694, wire_3655, wire_3654, wire_5191, wire_5190, wire_5181, wire_5180, wire_5171, wire_5170, wire_5161, wire_5160, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_4111, wire_4110, wire_4083, wire_4082, wire_4071, wire_4070, wire_4043, wire_4042, wire_4031, wire_4030, wire_4003, wire_4002, wire_3991, wire_3990, wire_3963, wire_3962, wire_4877, wire_4876, wire_4867, wire_4866, wire_4857, wire_4856, wire_4847, wire_4846, wire_4791, wire_4790, wire_4781, wire_4780, wire_4771, wire_4770, wire_4761, wire_4760, wire_3785, wire_3784, wire_3765, wire_3764, wire_3745, wire_3744, wire_3725, wire_3724, wire_3705, wire_3704, wire_3685, wire_3684, wire_3665, wire_3664, wire_3645, wire_3644, wire_5237, wire_5236, wire_5227, wire_5226, wire_5217, wire_5216, wire_5207, wire_5206, wire_5151, wire_5150, wire_5141, wire_5140, wire_5131, wire_5130, wire_5121, wire_5120, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_4081, wire_4080, wire_4041, wire_4040, wire_4001, wire_4000, wire_3961, wire_3960, wire_4911, wire_4910, wire_4901, wire_4900, wire_4891, wire_4890, wire_4881, wire_4880, wire_4837, wire_4836, wire_4827, wire_4826, wire_4817, wire_4816, wire_4807, wire_4806, wire_3781, wire_3780, wire_3761, wire_3760, wire_3741, wire_3740, wire_3721, wire_3720, wire_3701, wire_3700, wire_3681, wire_3680, wire_3661, wire_3660, wire_3641, wire_3640, wire_5195, wire_5194, wire_5185, wire_5184, wire_5175, wire_5174, wire_5165, wire_5164, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_4099, wire_4098, wire_4087, wire_4086, wire_4059, wire_4058, wire_4047, wire_4046, wire_4019, wire_4018, wire_4007, wire_4006, wire_3979, wire_3978, wire_3967, wire_3966, wire_4915, wire_4914, wire_4905, wire_4904, wire_4895, wire_4894, wire_4885, wire_4884, wire_4831, wire_4830, wire_4821, wire_4820, wire_4811, wire_4810, wire_4801, wire_4800, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_3767, wire_3766, wire_3727, wire_3726, wire_3687, wire_3686, wire_3647, wire_3646, wire_5231, wire_5230, wire_5221, wire_5220, wire_5211, wire_5210, wire_5201, wire_5200, wire_5155, wire_5154, wire_5145, wire_5144, wire_5135, wire_5134, wire_5125, wire_5124, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_4097, wire_4096, wire_4057, wire_4056, wire_4017, wire_4016, wire_3977, wire_3976};
    // IPIN TOTAL: 528
    assign lut_tile_1_3_ipin_in = {wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_2833, wire_2832, wire_2793, wire_2792, wire_2753, wire_2752, wire_2713, wire_2712, wire_5075, wire_5074, wire_5063, wire_5062, wire_5035, wire_5034, wire_5023, wire_5022, wire_4995, wire_4994, wire_4983, wire_4982, wire_4955, wire_4954, wire_4943, wire_4942, wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_2503, wire_2502, wire_2463, wire_2462, wire_2423, wire_2422, wire_2383, wire_2382, wire_5399, wire_5398, wire_5379, wire_5378, wire_5359, wire_5358, wire_5339, wire_5338, wire_5319, wire_5318, wire_5299, wire_5298, wire_5279, wire_5278, wire_5259, wire_5258, wire_2919, wire_2918, wire_2909, wire_2908, wire_2899, wire_2898, wire_2889, wire_2888, wire_2819, wire_2818, wire_2779, wire_2778, wire_2739, wire_2738, wire_2699, wire_2698, wire_5073, wire_5072, wire_5061, wire_5060, wire_5033, wire_5032, wire_5021, wire_5020, wire_4993, wire_4992, wire_4981, wire_4980, wire_4953, wire_4952, wire_4941, wire_4940, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_2519, wire_2518, wire_2479, wire_2478, wire_2439, wire_2438, wire_2399, wire_2398, wire_5397, wire_5396, wire_5369, wire_5368, wire_5357, wire_5356, wire_5329, wire_5328, wire_5317, wire_5316, wire_5289, wire_5288, wire_5277, wire_5276, wire_5249, wire_5248, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_2809, wire_2808, wire_2769, wire_2768, wire_2729, wire_2728, wire_2689, wire_2688, wire_5077, wire_5076, wire_5049, wire_5048, wire_5037, wire_5036, wire_5009, wire_5008, wire_4997, wire_4996, wire_4969, wire_4968, wire_4957, wire_4956, wire_4929, wire_4928, wire_2599, wire_2598, wire_2589, wire_2588, wire_2579, wire_2578, wire_2569, wire_2568, wire_2489, wire_2488, wire_2449, wire_2448, wire_2409, wire_2408, wire_2369, wire_2368, wire_5395, wire_5394, wire_5375, wire_5374, wire_5355, wire_5354, wire_5335, wire_5334, wire_5315, wire_5314, wire_5295, wire_5294, wire_5275, wire_5274, wire_5255, wire_5254, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_2835, wire_2834, wire_2795, wire_2794, wire_2755, wire_2754, wire_2715, wire_2714, wire_5067, wire_5066, wire_5055, wire_5054, wire_5027, wire_5026, wire_5015, wire_5014, wire_4987, wire_4986, wire_4975, wire_4974, wire_4947, wire_4946, wire_4935, wire_4934, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_2495, wire_2494, wire_2455, wire_2454, wire_2415, wire_2414, wire_2375, wire_2374, wire_5385, wire_5384, wire_5373, wire_5372, wire_5345, wire_5344, wire_5333, wire_5332, wire_5305, wire_5304, wire_5293, wire_5292, wire_5265, wire_5264, wire_5253, wire_5252, wire_2917, wire_2916, wire_2907, wire_2906, wire_2897, wire_2896, wire_2887, wire_2886, wire_2811, wire_2810, wire_2771, wire_2770, wire_2731, wire_2730, wire_2691, wire_2690, wire_5065, wire_5064, wire_5053, wire_5052, wire_5025, wire_5024, wire_5013, wire_5012, wire_4985, wire_4984, wire_4973, wire_4972, wire_4945, wire_4944, wire_4933, wire_4932, wire_2593, wire_2592, wire_2583, wire_2582, wire_2573, wire_2572, wire_2563, wire_2562, wire_2505, wire_2504, wire_2465, wire_2464, wire_2425, wire_2424, wire_2385, wire_2384, wire_5389, wire_5388, wire_5361, wire_5360, wire_5349, wire_5348, wire_5321, wire_5320, wire_5309, wire_5308, wire_5281, wire_5280, wire_5269, wire_5268, wire_5241, wire_5240, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_2801, wire_2800, wire_2761, wire_2760, wire_2721, wire_2720, wire_2681, wire_2680, wire_5071, wire_5070, wire_5043, wire_5042, wire_5031, wire_5030, wire_5003, wire_5002, wire_4991, wire_4990, wire_4963, wire_4962, wire_4951, wire_4950, wire_4923, wire_4922, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_2511, wire_2510, wire_2471, wire_2470, wire_2431, wire_2430, wire_2391, wire_2390, wire_5387, wire_5386, wire_5367, wire_5366, wire_5347, wire_5346, wire_5327, wire_5326, wire_5307, wire_5306, wire_5287, wire_5286, wire_5267, wire_5266, wire_5247, wire_5246, wire_2911, wire_2910, wire_2901, wire_2900, wire_2891, wire_2890, wire_2881, wire_2880, wire_2827, wire_2826, wire_2787, wire_2786, wire_2747, wire_2746, wire_2707, wire_2706, wire_5069, wire_5068, wire_5041, wire_5040, wire_5029, wire_5028, wire_5001, wire_5000, wire_4989, wire_4988, wire_4961, wire_4960, wire_4949, wire_4948, wire_4921, wire_4920, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_2487, wire_2486, wire_2447, wire_2446, wire_2407, wire_2406, wire_2367, wire_2366, wire_5377, wire_5376, wire_5365, wire_5364, wire_5337, wire_5336, wire_5325, wire_5324, wire_5297, wire_5296, wire_5285, wire_5284, wire_5257, wire_5256, wire_5245, wire_5244, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_2817, wire_2816, wire_2777, wire_2776, wire_2737, wire_2736, wire_2697, wire_2696, wire_5057, wire_5056, wire_5045, wire_5044, wire_5017, wire_5016, wire_5005, wire_5004, wire_4977, wire_4976, wire_4965, wire_4964, wire_4937, wire_4936, wire_4925, wire_4924, wire_2591, wire_2590, wire_2581, wire_2580, wire_2571, wire_2570, wire_2561, wire_2560, wire_2497, wire_2496, wire_2457, wire_2456, wire_2417, wire_2416, wire_2377, wire_2376, wire_5383, wire_5382, wire_5363, wire_5362, wire_5343, wire_5342, wire_5323, wire_5322, wire_5303, wire_5302, wire_5283, wire_5282, wire_5263, wire_5262, wire_5243, wire_5242, wire_2915, wire_2914, wire_2905, wire_2904, wire_2895, wire_2894, wire_2885, wire_2884, wire_2803, wire_2802, wire_2763, wire_2762, wire_2723, wire_2722, wire_2683, wire_2682};
    // IPIN TOTAL: 528
    assign lut_tile_2_3_ipin_in = {wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_3139, wire_3138, wire_3099, wire_3098, wire_3059, wire_3058, wire_3019, wire_3018, wire_5073, wire_5072, wire_5061, wire_5060, wire_5033, wire_5032, wire_5021, wire_5020, wire_4993, wire_4992, wire_4981, wire_4980, wire_4953, wire_4952, wire_4941, wire_4940, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_2833, wire_2832, wire_2793, wire_2792, wire_2753, wire_2752, wire_2713, wire_2712, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_5397, wire_5396, wire_5357, wire_5356, wire_5317, wire_5316, wire_5277, wire_5276, wire_3235, wire_3234, wire_3225, wire_3224, wire_3215, wire_3214, wire_3205, wire_3204, wire_3157, wire_3156, wire_3117, wire_3116, wire_3077, wire_3076, wire_3037, wire_3036, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_5059, wire_5058, wire_5019, wire_5018, wire_4979, wire_4978, wire_4939, wire_4938, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_2809, wire_2808, wire_2769, wire_2768, wire_2729, wire_2728, wire_2689, wire_2688, wire_5395, wire_5394, wire_5375, wire_5374, wire_5355, wire_5354, wire_5335, wire_5334, wire_5315, wire_5314, wire_5295, wire_5294, wire_5275, wire_5274, wire_5255, wire_5254, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_3155, wire_3154, wire_3115, wire_3114, wire_3075, wire_3074, wire_3035, wire_3034, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_5075, wire_5074, wire_5035, wire_5034, wire_4995, wire_4994, wire_4955, wire_4954, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_2835, wire_2834, wire_2795, wire_2794, wire_2755, wire_2754, wire_2715, wire_2714, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_5373, wire_5372, wire_5333, wire_5332, wire_5293, wire_5292, wire_5253, wire_5252, wire_3239, wire_3238, wire_3229, wire_3228, wire_3219, wire_3218, wire_3209, wire_3208, wire_3133, wire_3132, wire_3093, wire_3092, wire_3053, wire_3052, wire_3013, wire_3012, wire_5065, wire_5064, wire_5053, wire_5052, wire_5025, wire_5024, wire_5013, wire_5012, wire_4985, wire_4984, wire_4973, wire_4972, wire_4945, wire_4944, wire_4933, wire_4932, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_2825, wire_2824, wire_2785, wire_2784, wire_2745, wire_2744, wire_2705, wire_2704, wire_5391, wire_5390, wire_5371, wire_5370, wire_5351, wire_5350, wire_5331, wire_5330, wire_5311, wire_5310, wire_5291, wire_5290, wire_5271, wire_5270, wire_5251, wire_5250, wire_3233, wire_3232, wire_3223, wire_3222, wire_3213, wire_3212, wire_3203, wire_3202, wire_3149, wire_3148, wire_3109, wire_3108, wire_3069, wire_3068, wire_3029, wire_3028, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_5051, wire_5050, wire_5011, wire_5010, wire_4971, wire_4970, wire_4931, wire_4930, wire_2917, wire_2916, wire_2907, wire_2906, wire_2897, wire_2896, wire_2887, wire_2886, wire_2811, wire_2810, wire_2771, wire_2770, wire_2731, wire_2730, wire_2691, wire_2690, wire_5387, wire_5386, wire_5367, wire_5366, wire_5347, wire_5346, wire_5327, wire_5326, wire_5307, wire_5306, wire_5287, wire_5286, wire_5267, wire_5266, wire_5247, wire_5246, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_3147, wire_3146, wire_3107, wire_3106, wire_3067, wire_3066, wire_3027, wire_3026, wire_5069, wire_5068, wire_5041, wire_5040, wire_5029, wire_5028, wire_5001, wire_5000, wire_4989, wire_4988, wire_4961, wire_4960, wire_4949, wire_4948, wire_4921, wire_4920, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_2801, wire_2800, wire_2761, wire_2760, wire_2721, wire_2720, wire_2681, wire_2680, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_5365, wire_5364, wire_5325, wire_5324, wire_5285, wire_5284, wire_5245, wire_5244, wire_3237, wire_3236, wire_3227, wire_3226, wire_3217, wire_3216, wire_3207, wire_3206, wire_3125, wire_3124, wire_3085, wire_3084, wire_3045, wire_3044, wire_3005, wire_3004, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_5067, wire_5066, wire_5027, wire_5026, wire_4987, wire_4986, wire_4947, wire_4946, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_2817, wire_2816, wire_2777, wire_2776, wire_2737, wire_2736, wire_2697, wire_2696, wire_5383, wire_5382, wire_5363, wire_5362, wire_5343, wire_5342, wire_5323, wire_5322, wire_5303, wire_5302, wire_5283, wire_5282, wire_5263, wire_5262, wire_5243, wire_5242, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_3123, wire_3122, wire_3083, wire_3082, wire_3043, wire_3042, wire_3003, wire_3002, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_5043, wire_5042, wire_5003, wire_5002, wire_4963, wire_4962, wire_4923, wire_4922, wire_2915, wire_2914, wire_2905, wire_2904, wire_2895, wire_2894, wire_2885, wire_2884, wire_2803, wire_2802, wire_2763, wire_2762, wire_2723, wire_2722, wire_2683, wire_2682, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_5381, wire_5380, wire_5341, wire_5340, wire_5301, wire_5300, wire_5261, wire_5260, wire_3231, wire_3230, wire_3221, wire_3220, wire_3211, wire_3210, wire_3201, wire_3200, wire_3141, wire_3140, wire_3101, wire_3100, wire_3061, wire_3060, wire_3021, wire_3020};
    // IPIN TOTAL: 528
    assign lut_tile_3_3_ipin_in = {wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_3477, wire_3476, wire_3437, wire_3436, wire_3397, wire_3396, wire_3357, wire_3356, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_5059, wire_5058, wire_5019, wire_5018, wire_4979, wire_4978, wire_4939, wire_4938, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_3139, wire_3138, wire_3099, wire_3098, wire_3059, wire_3058, wire_3019, wire_3018, wire_5479, wire_5478, wire_5469, wire_5468, wire_5459, wire_5458, wire_5449, wire_5448, wire_5383, wire_5382, wire_5343, wire_5342, wire_5303, wire_5302, wire_5263, wire_5262, wire_3559, wire_3558, wire_3549, wire_3548, wire_3539, wire_3538, wire_3529, wire_3528, wire_3463, wire_3462, wire_3423, wire_3422, wire_3383, wire_3382, wire_3343, wire_3342, wire_5155, wire_5154, wire_5145, wire_5144, wire_5135, wire_5134, wire_5125, wire_5124, wire_5077, wire_5076, wire_5037, wire_5036, wire_4997, wire_4996, wire_4957, wire_4956, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_3155, wire_3154, wire_3115, wire_3114, wire_3075, wire_3074, wire_3035, wire_3034, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_5373, wire_5372, wire_5333, wire_5332, wire_5293, wire_5292, wire_5253, wire_5252, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_3453, wire_3452, wire_3413, wire_3412, wire_3373, wire_3372, wire_3333, wire_3332, wire_5159, wire_5158, wire_5149, wire_5148, wire_5139, wire_5138, wire_5129, wire_5128, wire_5053, wire_5052, wire_5013, wire_5012, wire_4973, wire_4972, wire_4933, wire_4932, wire_3239, wire_3238, wire_3229, wire_3228, wire_3219, wire_3218, wire_3209, wire_3208, wire_3133, wire_3132, wire_3093, wire_3092, wire_3053, wire_3052, wire_3013, wire_3012, wire_5473, wire_5472, wire_5463, wire_5462, wire_5453, wire_5452, wire_5443, wire_5442, wire_5399, wire_5398, wire_5359, wire_5358, wire_5319, wire_5318, wire_5279, wire_5278, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_3479, wire_3478, wire_3439, wire_3438, wire_3399, wire_3398, wire_3359, wire_3358, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_5051, wire_5050, wire_5011, wire_5010, wire_4971, wire_4970, wire_4931, wire_4930, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_3131, wire_3130, wire_3091, wire_3090, wire_3051, wire_3050, wire_3011, wire_3010, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_5389, wire_5388, wire_5349, wire_5348, wire_5309, wire_5308, wire_5269, wire_5268, wire_3557, wire_3556, wire_3547, wire_3546, wire_3537, wire_3536, wire_3527, wire_3526, wire_3455, wire_3454, wire_3415, wire_3414, wire_3375, wire_3374, wire_3335, wire_3334, wire_5153, wire_5152, wire_5143, wire_5142, wire_5133, wire_5132, wire_5123, wire_5122, wire_5069, wire_5068, wire_5029, wire_5028, wire_4989, wire_4988, wire_4949, wire_4948, wire_3233, wire_3232, wire_3223, wire_3222, wire_3213, wire_3212, wire_3203, wire_3202, wire_3149, wire_3148, wire_3109, wire_3108, wire_3069, wire_3068, wire_3029, wire_3028, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_5365, wire_5364, wire_5325, wire_5324, wire_5285, wire_5284, wire_5245, wire_5244, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_3445, wire_3444, wire_3405, wire_3404, wire_3365, wire_3364, wire_3325, wire_3324, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_5067, wire_5066, wire_5027, wire_5026, wire_4987, wire_4986, wire_4947, wire_4946, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_3147, wire_3146, wire_3107, wire_3106, wire_3067, wire_3066, wire_3027, wire_3026, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_5391, wire_5390, wire_5351, wire_5350, wire_5311, wire_5310, wire_5271, wire_5270, wire_3551, wire_3550, wire_3541, wire_3540, wire_3531, wire_3530, wire_3521, wire_3520, wire_3471, wire_3470, wire_3431, wire_3430, wire_3391, wire_3390, wire_3351, wire_3350, wire_5157, wire_5156, wire_5147, wire_5146, wire_5137, wire_5136, wire_5127, wire_5126, wire_5045, wire_5044, wire_5005, wire_5004, wire_4965, wire_4964, wire_4925, wire_4924, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_3123, wire_3122, wire_3083, wire_3082, wire_3043, wire_3042, wire_3003, wire_3002, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_5381, wire_5380, wire_5341, wire_5340, wire_5301, wire_5300, wire_5261, wire_5260, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_3461, wire_3460, wire_3421, wire_3420, wire_3381, wire_3380, wire_3341, wire_3340, wire_5151, wire_5150, wire_5141, wire_5140, wire_5131, wire_5130, wire_5121, wire_5120, wire_5061, wire_5060, wire_5021, wire_5020, wire_4981, wire_4980, wire_4941, wire_4940, wire_3231, wire_3230, wire_3221, wire_3220, wire_3211, wire_3210, wire_3201, wire_3200, wire_3141, wire_3140, wire_3101, wire_3100, wire_3061, wire_3060, wire_3021, wire_3020, wire_5475, wire_5474, wire_5465, wire_5464, wire_5455, wire_5454, wire_5445, wire_5444, wire_5367, wire_5366, wire_5327, wire_5326, wire_5287, wire_5286, wire_5247, wire_5246, wire_3555, wire_3554, wire_3545, wire_3544, wire_3535, wire_3534, wire_3525, wire_3524, wire_3447, wire_3446, wire_3407, wire_3406, wire_3367, wire_3366, wire_3327, wire_3326};
    // IPIN TOTAL: 528
    assign lut_tile_4_3_ipin_in = {wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_3783, wire_3782, wire_3743, wire_3742, wire_3703, wire_3702, wire_3663, wire_3662, wire_5155, wire_5154, wire_5145, wire_5144, wire_5135, wire_5134, wire_5125, wire_5124, wire_5077, wire_5076, wire_5037, wire_5036, wire_4997, wire_4996, wire_4957, wire_4956, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_3477, wire_3476, wire_3437, wire_3436, wire_3397, wire_3396, wire_3357, wire_3356, wire_5515, wire_5514, wire_5505, wire_5504, wire_5495, wire_5494, wire_5485, wire_5484, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_3875, wire_3874, wire_3865, wire_3864, wire_3855, wire_3854, wire_3845, wire_3844, wire_3793, wire_3792, wire_3753, wire_3752, wire_3713, wire_3712, wire_3673, wire_3672, wire_5199, wire_5198, wire_5189, wire_5188, wire_5179, wire_5178, wire_5169, wire_5168, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_3453, wire_3452, wire_3413, wire_3412, wire_3373, wire_3372, wire_3333, wire_3332, wire_5473, wire_5472, wire_5463, wire_5462, wire_5453, wire_5452, wire_5443, wire_5442, wire_5399, wire_5398, wire_5359, wire_5358, wire_5319, wire_5318, wire_5279, wire_5278, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_3799, wire_3798, wire_3759, wire_3758, wire_3719, wire_3718, wire_3679, wire_3678, wire_5193, wire_5192, wire_5183, wire_5182, wire_5173, wire_5172, wire_5163, wire_5162, wire_5119, wire_5118, wire_5109, wire_5108, wire_5099, wire_5098, wire_5089, wire_5088, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_3479, wire_3478, wire_3439, wire_3438, wire_3399, wire_3398, wire_3359, wire_3358, wire_5519, wire_5518, wire_5509, wire_5508, wire_5499, wire_5498, wire_5489, wire_5488, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_3879, wire_3878, wire_3869, wire_3868, wire_3859, wire_3858, wire_3849, wire_3848, wire_3769, wire_3768, wire_3729, wire_3728, wire_3689, wire_3688, wire_3649, wire_3648, wire_5153, wire_5152, wire_5143, wire_5142, wire_5133, wire_5132, wire_5123, wire_5122, wire_5069, wire_5068, wire_5029, wire_5028, wire_4989, wire_4988, wire_4949, wire_4948, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_3469, wire_3468, wire_3429, wire_3428, wire_3389, wire_3388, wire_3349, wire_3348, wire_5477, wire_5476, wire_5467, wire_5466, wire_5457, wire_5456, wire_5447, wire_5446, wire_5375, wire_5374, wire_5335, wire_5334, wire_5295, wire_5294, wire_5255, wire_5254, wire_3873, wire_3872, wire_3863, wire_3862, wire_3853, wire_3852, wire_3843, wire_3842, wire_3785, wire_3784, wire_3745, wire_3744, wire_3705, wire_3704, wire_3665, wire_3664, wire_5197, wire_5196, wire_5187, wire_5186, wire_5177, wire_5176, wire_5167, wire_5166, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_3557, wire_3556, wire_3547, wire_3546, wire_3537, wire_3536, wire_3527, wire_3526, wire_3455, wire_3454, wire_3415, wire_3414, wire_3375, wire_3374, wire_3335, wire_3334, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_5391, wire_5390, wire_5351, wire_5350, wire_5311, wire_5310, wire_5271, wire_5270, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_3791, wire_3790, wire_3751, wire_3750, wire_3711, wire_3710, wire_3671, wire_3670, wire_5157, wire_5156, wire_5147, wire_5146, wire_5137, wire_5136, wire_5127, wire_5126, wire_5045, wire_5044, wire_5005, wire_5004, wire_4965, wire_4964, wire_4925, wire_4924, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_3445, wire_3444, wire_3405, wire_3404, wire_3365, wire_3364, wire_3325, wire_3324, wire_5517, wire_5516, wire_5507, wire_5506, wire_5497, wire_5496, wire_5487, wire_5486, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_3877, wire_3876, wire_3867, wire_3866, wire_3857, wire_3856, wire_3847, wire_3846, wire_3761, wire_3760, wire_3721, wire_3720, wire_3681, wire_3680, wire_3641, wire_3640, wire_5191, wire_5190, wire_5181, wire_5180, wire_5171, wire_5170, wire_5161, wire_5160, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_3461, wire_3460, wire_3421, wire_3420, wire_3381, wire_3380, wire_3341, wire_3340, wire_5475, wire_5474, wire_5465, wire_5464, wire_5455, wire_5454, wire_5445, wire_5444, wire_5367, wire_5366, wire_5327, wire_5326, wire_5287, wire_5286, wire_5247, wire_5246, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_3767, wire_3766, wire_3727, wire_3726, wire_3687, wire_3686, wire_3647, wire_3646, wire_5195, wire_5194, wire_5185, wire_5184, wire_5175, wire_5174, wire_5165, wire_5164, wire_5111, wire_5110, wire_5101, wire_5100, wire_5091, wire_5090, wire_5081, wire_5080, wire_3555, wire_3554, wire_3545, wire_3544, wire_3535, wire_3534, wire_3525, wire_3524, wire_3447, wire_3446, wire_3407, wire_3406, wire_3367, wire_3366, wire_3327, wire_3326, wire_5511, wire_5510, wire_5501, wire_5500, wire_5491, wire_5490, wire_5481, wire_5480, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_3871, wire_3870, wire_3861, wire_3860, wire_3851, wire_3850, wire_3841, wire_3840, wire_3777, wire_3776, wire_3737, wire_3736, wire_3697, wire_3696, wire_3657, wire_3656};
    // IPIN TOTAL: 528
    assign lut_tile_5_3_ipin_in = {wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_4113, wire_4112, wire_4073, wire_4072, wire_4033, wire_4032, wire_3993, wire_3992, wire_5199, wire_5198, wire_5189, wire_5188, wire_5179, wire_5178, wire_5169, wire_5168, wire_5115, wire_5114, wire_5105, wire_5104, wire_5095, wire_5094, wire_5085, wire_5084, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_3783, wire_3782, wire_3743, wire_3742, wire_3703, wire_3702, wire_3663, wire_3662, wire_5559, wire_5558, wire_5549, wire_5548, wire_5539, wire_5538, wire_5529, wire_5528, wire_5475, wire_5474, wire_5465, wire_5464, wire_5455, wire_5454, wire_5445, wire_5444, wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_4099, wire_4098, wire_4059, wire_4058, wire_4019, wire_4018, wire_3979, wire_3978, wire_5235, wire_5234, wire_5225, wire_5224, wire_5215, wire_5214, wire_5205, wire_5204, wire_5159, wire_5158, wire_5149, wire_5148, wire_5139, wire_5138, wire_5129, wire_5128, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_3799, wire_3798, wire_3759, wire_3758, wire_3719, wire_3718, wire_3679, wire_3678, wire_5519, wire_5518, wire_5509, wire_5508, wire_5499, wire_5498, wire_5489, wire_5488, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_4089, wire_4088, wire_4049, wire_4048, wire_4009, wire_4008, wire_3969, wire_3968, wire_5239, wire_5238, wire_5229, wire_5228, wire_5219, wire_5218, wire_5209, wire_5208, wire_5153, wire_5152, wire_5143, wire_5142, wire_5133, wire_5132, wire_5123, wire_5122, wire_3879, wire_3878, wire_3869, wire_3868, wire_3859, wire_3858, wire_3849, wire_3848, wire_3769, wire_3768, wire_3729, wire_3728, wire_3689, wire_3688, wire_3649, wire_3648, wire_5553, wire_5552, wire_5543, wire_5542, wire_5533, wire_5532, wire_5523, wire_5522, wire_5479, wire_5478, wire_5469, wire_5468, wire_5459, wire_5458, wire_5449, wire_5448, wire_4193, wire_4192, wire_4183, wire_4182, wire_4173, wire_4172, wire_4163, wire_4162, wire_4115, wire_4114, wire_4075, wire_4074, wire_4035, wire_4034, wire_3995, wire_3994, wire_5197, wire_5196, wire_5187, wire_5186, wire_5177, wire_5176, wire_5167, wire_5166, wire_5113, wire_5112, wire_5103, wire_5102, wire_5093, wire_5092, wire_5083, wire_5082, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_3775, wire_3774, wire_3735, wire_3734, wire_3695, wire_3694, wire_3655, wire_3654, wire_5513, wire_5512, wire_5503, wire_5502, wire_5493, wire_5492, wire_5483, wire_5482, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_4197, wire_4196, wire_4187, wire_4186, wire_4177, wire_4176, wire_4167, wire_4166, wire_4091, wire_4090, wire_4051, wire_4050, wire_4011, wire_4010, wire_3971, wire_3970, wire_5233, wire_5232, wire_5223, wire_5222, wire_5213, wire_5212, wire_5203, wire_5202, wire_5157, wire_5156, wire_5147, wire_5146, wire_5137, wire_5136, wire_5127, wire_5126, wire_3873, wire_3872, wire_3863, wire_3862, wire_3853, wire_3852, wire_3843, wire_3842, wire_3785, wire_3784, wire_3745, wire_3744, wire_3705, wire_3704, wire_3665, wire_3664, wire_5517, wire_5516, wire_5507, wire_5506, wire_5497, wire_5496, wire_5487, wire_5486, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_4081, wire_4080, wire_4041, wire_4040, wire_4001, wire_4000, wire_3961, wire_3960, wire_5191, wire_5190, wire_5181, wire_5180, wire_5171, wire_5170, wire_5161, wire_5160, wire_5117, wire_5116, wire_5107, wire_5106, wire_5097, wire_5096, wire_5087, wire_5086, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_3791, wire_3790, wire_3751, wire_3750, wire_3711, wire_3710, wire_3671, wire_3670, wire_5551, wire_5550, wire_5541, wire_5540, wire_5531, wire_5530, wire_5521, wire_5520, wire_5477, wire_5476, wire_5467, wire_5466, wire_5457, wire_5456, wire_5447, wire_5446, wire_4191, wire_4190, wire_4181, wire_4180, wire_4171, wire_4170, wire_4161, wire_4160, wire_4107, wire_4106, wire_4067, wire_4066, wire_4027, wire_4026, wire_3987, wire_3986, wire_5237, wire_5236, wire_5227, wire_5226, wire_5217, wire_5216, wire_5207, wire_5206, wire_5151, wire_5150, wire_5141, wire_5140, wire_5131, wire_5130, wire_5121, wire_5120, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_3767, wire_3766, wire_3727, wire_3726, wire_3687, wire_3686, wire_3647, wire_3646, wire_5511, wire_5510, wire_5501, wire_5500, wire_5491, wire_5490, wire_5481, wire_5480, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_4097, wire_4096, wire_4057, wire_4056, wire_4017, wire_4016, wire_3977, wire_3976, wire_5231, wire_5230, wire_5221, wire_5220, wire_5211, wire_5210, wire_5201, wire_5200, wire_5155, wire_5154, wire_5145, wire_5144, wire_5135, wire_5134, wire_5125, wire_5124, wire_3871, wire_3870, wire_3861, wire_3860, wire_3851, wire_3850, wire_3841, wire_3840, wire_3777, wire_3776, wire_3737, wire_3736, wire_3697, wire_3696, wire_3657, wire_3656, wire_5555, wire_5554, wire_5545, wire_5544, wire_5535, wire_5534, wire_5525, wire_5524, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_4083, wire_4082, wire_4043, wire_4042, wire_4003, wire_4002, wire_3963, wire_3962};
    // IPIN TOTAL: 528
    assign lut_tile_1_4_ipin_in = {wire_2919, wire_2918, wire_2909, wire_2908, wire_2899, wire_2898, wire_2889, wire_2888, wire_2819, wire_2818, wire_2779, wire_2778, wire_2739, wire_2738, wire_2699, wire_2698, wire_5393, wire_5392, wire_5381, wire_5380, wire_5353, wire_5352, wire_5341, wire_5340, wire_5313, wire_5312, wire_5301, wire_5300, wire_5273, wire_5272, wire_5261, wire_5260, wire_2595, wire_2594, wire_2585, wire_2584, wire_2575, wire_2574, wire_2565, wire_2564, wire_2513, wire_2512, wire_2473, wire_2472, wire_2433, wire_2432, wire_2393, wire_2392, wire_5717, wire_5716, wire_5697, wire_5696, wire_5677, wire_5676, wire_5657, wire_5656, wire_5637, wire_5636, wire_5617, wire_5616, wire_5597, wire_5596, wire_5577, wire_5576, wire_2955, wire_2954, wire_2945, wire_2944, wire_2935, wire_2934, wire_2925, wire_2924, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_5399, wire_5398, wire_5379, wire_5378, wire_5359, wire_5358, wire_5339, wire_5338, wire_5319, wire_5318, wire_5299, wire_5298, wire_5279, wire_5278, wire_5259, wire_5258, wire_2599, wire_2598, wire_2589, wire_2588, wire_2579, wire_2578, wire_2569, wire_2568, wire_2489, wire_2488, wire_2449, wire_2448, wire_2409, wire_2408, wire_2369, wire_2368, wire_5715, wire_5714, wire_5695, wire_5694, wire_5675, wire_5674, wire_5655, wire_5654, wire_5635, wire_5634, wire_5615, wire_5614, wire_5595, wire_5594, wire_5575, wire_5574, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_2835, wire_2834, wire_2795, wire_2794, wire_2755, wire_2754, wire_2715, wire_2714, wire_5395, wire_5394, wire_5375, wire_5374, wire_5355, wire_5354, wire_5335, wire_5334, wire_5315, wire_5314, wire_5295, wire_5294, wire_5275, wire_5274, wire_5255, wire_5254, wire_2633, wire_2632, wire_2623, wire_2622, wire_2613, wire_2612, wire_2603, wire_2602, wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_5713, wire_5712, wire_5693, wire_5692, wire_5673, wire_5672, wire_5653, wire_5652, wire_5633, wire_5632, wire_5613, wire_5612, wire_5593, wire_5592, wire_5573, wire_5572, wire_2959, wire_2958, wire_2949, wire_2948, wire_2939, wire_2938, wire_2929, wire_2928, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_5385, wire_5384, wire_5373, wire_5372, wire_5345, wire_5344, wire_5333, wire_5332, wire_5305, wire_5304, wire_5293, wire_5292, wire_5265, wire_5264, wire_5253, wire_5252, wire_2593, wire_2592, wire_2583, wire_2582, wire_2573, wire_2572, wire_2563, wire_2562, wire_2505, wire_2504, wire_2465, wire_2464, wire_2425, wire_2424, wire_2385, wire_2384, wire_5711, wire_5710, wire_5691, wire_5690, wire_5671, wire_5670, wire_5651, wire_5650, wire_5631, wire_5630, wire_5611, wire_5610, wire_5591, wire_5590, wire_5571, wire_5570, wire_2953, wire_2952, wire_2943, wire_2942, wire_2933, wire_2932, wire_2923, wire_2922, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_5391, wire_5390, wire_5371, wire_5370, wire_5351, wire_5350, wire_5331, wire_5330, wire_5311, wire_5310, wire_5291, wire_5290, wire_5271, wire_5270, wire_5251, wire_5250, wire_2637, wire_2636, wire_2627, wire_2626, wire_2617, wire_2616, wire_2607, wire_2606, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_5707, wire_5706, wire_5687, wire_5686, wire_5667, wire_5666, wire_5647, wire_5646, wire_5627, wire_5626, wire_5607, wire_5606, wire_5587, wire_5586, wire_5567, wire_5566, wire_2911, wire_2910, wire_2901, wire_2900, wire_2891, wire_2890, wire_2881, wire_2880, wire_2827, wire_2826, wire_2787, wire_2786, wire_2747, wire_2746, wire_2707, wire_2706, wire_5389, wire_5388, wire_5361, wire_5360, wire_5349, wire_5348, wire_5321, wire_5320, wire_5309, wire_5308, wire_5281, wire_5280, wire_5269, wire_5268, wire_5241, wire_5240, wire_2597, wire_2596, wire_2587, wire_2586, wire_2577, wire_2576, wire_2567, wire_2566, wire_2481, wire_2480, wire_2441, wire_2440, wire_2401, wire_2400, wire_2361, wire_2360, wire_5705, wire_5704, wire_5685, wire_5684, wire_5665, wire_5664, wire_5645, wire_5644, wire_5625, wire_5624, wire_5605, wire_5604, wire_5585, wire_5584, wire_5565, wire_5564, wire_2957, wire_2956, wire_2947, wire_2946, wire_2937, wire_2936, wire_2927, wire_2926, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_5387, wire_5386, wire_5367, wire_5366, wire_5347, wire_5346, wire_5327, wire_5326, wire_5307, wire_5306, wire_5287, wire_5286, wire_5267, wire_5266, wire_5247, wire_5246, wire_2591, wire_2590, wire_2581, wire_2580, wire_2571, wire_2570, wire_2561, wire_2560, wire_2497, wire_2496, wire_2457, wire_2456, wire_2417, wire_2416, wire_2377, wire_2376, wire_5703, wire_5702, wire_5683, wire_5682, wire_5663, wire_5662, wire_5643, wire_5642, wire_5623, wire_5622, wire_5603, wire_5602, wire_5583, wire_5582, wire_5563, wire_5562, wire_2915, wire_2914, wire_2905, wire_2904, wire_2895, wire_2894, wire_2885, wire_2884, wire_2803, wire_2802, wire_2763, wire_2762, wire_2723, wire_2722, wire_2683, wire_2682, wire_5383, wire_5382, wire_5363, wire_5362, wire_5343, wire_5342, wire_5323, wire_5322, wire_5303, wire_5302, wire_5283, wire_5282, wire_5263, wire_5262, wire_5243, wire_5242, wire_2635, wire_2634, wire_2625, wire_2624, wire_2615, wire_2614, wire_2605, wire_2604, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_5701, wire_5700, wire_5681, wire_5680, wire_5661, wire_5660, wire_5641, wire_5640, wire_5621, wire_5620, wire_5601, wire_5600, wire_5581, wire_5580, wire_5561, wire_5560, wire_2951, wire_2950, wire_2941, wire_2940, wire_2931, wire_2930, wire_2921, wire_2920, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844};
    // IPIN TOTAL: 528
    assign lut_tile_2_4_ipin_in = {wire_3235, wire_3234, wire_3225, wire_3224, wire_3215, wire_3214, wire_3205, wire_3204, wire_3157, wire_3156, wire_3117, wire_3116, wire_3077, wire_3076, wire_3037, wire_3036, wire_5399, wire_5398, wire_5379, wire_5378, wire_5359, wire_5358, wire_5339, wire_5338, wire_5319, wire_5318, wire_5299, wire_5298, wire_5279, wire_5278, wire_5259, wire_5258, wire_2919, wire_2918, wire_2909, wire_2908, wire_2899, wire_2898, wire_2889, wire_2888, wire_2819, wire_2818, wire_2779, wire_2778, wire_2739, wire_2738, wire_2699, wire_2698, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_5703, wire_5702, wire_5663, wire_5662, wire_5623, wire_5622, wire_5583, wire_5582, wire_3279, wire_3278, wire_3269, wire_3268, wire_3259, wire_3258, wire_3249, wire_3248, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_5397, wire_5396, wire_5357, wire_5356, wire_5317, wire_5316, wire_5277, wire_5276, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_2835, wire_2834, wire_2795, wire_2794, wire_2755, wire_2754, wire_2715, wire_2714, wire_5713, wire_5712, wire_5693, wire_5692, wire_5673, wire_5672, wire_5653, wire_5652, wire_5633, wire_5632, wire_5613, wire_5612, wire_5593, wire_5592, wire_5573, wire_5572, wire_3239, wire_3238, wire_3229, wire_3228, wire_3219, wire_3218, wire_3209, wire_3208, wire_3133, wire_3132, wire_3093, wire_3092, wire_3053, wire_3052, wire_3013, wire_3012, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_5373, wire_5372, wire_5333, wire_5332, wire_5293, wire_5292, wire_5253, wire_5252, wire_2959, wire_2958, wire_2949, wire_2948, wire_2939, wire_2938, wire_2929, wire_2928, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_5719, wire_5718, wire_5679, wire_5678, wire_5639, wire_5638, wire_5599, wire_5598, wire_3273, wire_3272, wire_3263, wire_3262, wire_3253, wire_3252, wire_3243, wire_3242, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_5391, wire_5390, wire_5371, wire_5370, wire_5351, wire_5350, wire_5331, wire_5330, wire_5311, wire_5310, wire_5291, wire_5290, wire_5271, wire_5270, wire_5251, wire_5250, wire_2917, wire_2916, wire_2907, wire_2906, wire_2897, wire_2896, wire_2887, wire_2886, wire_2811, wire_2810, wire_2771, wire_2770, wire_2731, wire_2730, wire_2691, wire_2690, wire_5709, wire_5708, wire_5689, wire_5688, wire_5669, wire_5668, wire_5649, wire_5648, wire_5629, wire_5628, wire_5609, wire_5608, wire_5589, wire_5588, wire_5569, wire_5568, wire_3277, wire_3276, wire_3267, wire_3266, wire_3257, wire_3256, wire_3247, wire_3246, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_5389, wire_5388, wire_5349, wire_5348, wire_5309, wire_5308, wire_5269, wire_5268, wire_2953, wire_2952, wire_2943, wire_2942, wire_2933, wire_2932, wire_2923, wire_2922, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_5705, wire_5704, wire_5685, wire_5684, wire_5665, wire_5664, wire_5645, wire_5644, wire_5625, wire_5624, wire_5605, wire_5604, wire_5585, wire_5584, wire_5565, wire_5564, wire_3237, wire_3236, wire_3227, wire_3226, wire_3217, wire_3216, wire_3207, wire_3206, wire_3125, wire_3124, wire_3085, wire_3084, wire_3045, wire_3044, wire_3005, wire_3004, wire_5387, wire_5386, wire_5367, wire_5366, wire_5347, wire_5346, wire_5327, wire_5326, wire_5307, wire_5306, wire_5287, wire_5286, wire_5267, wire_5266, wire_5247, wire_5246, wire_2911, wire_2910, wire_2901, wire_2900, wire_2891, wire_2890, wire_2881, wire_2880, wire_2827, wire_2826, wire_2787, wire_2786, wire_2747, wire_2746, wire_2707, wire_2706, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_5711, wire_5710, wire_5671, wire_5670, wire_5631, wire_5630, wire_5591, wire_5590, wire_3271, wire_3270, wire_3261, wire_3260, wire_3251, wire_3250, wire_3241, wire_3240, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_5365, wire_5364, wire_5325, wire_5324, wire_5285, wire_5284, wire_5245, wire_5244, wire_2915, wire_2914, wire_2905, wire_2904, wire_2895, wire_2894, wire_2885, wire_2884, wire_2803, wire_2802, wire_2763, wire_2762, wire_2723, wire_2722, wire_2683, wire_2682, wire_5701, wire_5700, wire_5681, wire_5680, wire_5661, wire_5660, wire_5641, wire_5640, wire_5621, wire_5620, wire_5601, wire_5600, wire_5581, wire_5580, wire_5561, wire_5560, wire_3231, wire_3230, wire_3221, wire_3220, wire_3211, wire_3210, wire_3201, wire_3200, wire_3141, wire_3140, wire_3101, wire_3100, wire_3061, wire_3060, wire_3021, wire_3020, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_5381, wire_5380, wire_5341, wire_5340, wire_5301, wire_5300, wire_5261, wire_5260, wire_2951, wire_2950, wire_2941, wire_2940, wire_2931, wire_2930, wire_2921, wire_2920, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_5687, wire_5686, wire_5647, wire_5646, wire_5607, wire_5606, wire_5567, wire_5566, wire_3275, wire_3274, wire_3265, wire_3264, wire_3255, wire_3254, wire_3245, wire_3244, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160};
    // IPIN TOTAL: 528
    assign lut_tile_3_4_ipin_in = {wire_3559, wire_3558, wire_3549, wire_3548, wire_3539, wire_3538, wire_3529, wire_3528, wire_3463, wire_3462, wire_3423, wire_3422, wire_3383, wire_3382, wire_3343, wire_3342, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_5397, wire_5396, wire_5357, wire_5356, wire_5317, wire_5316, wire_5277, wire_5276, wire_3235, wire_3234, wire_3225, wire_3224, wire_3215, wire_3214, wire_3205, wire_3204, wire_3157, wire_3156, wire_3117, wire_3116, wire_3077, wire_3076, wire_3037, wire_3036, wire_5795, wire_5794, wire_5785, wire_5784, wire_5775, wire_5774, wire_5765, wire_5764, wire_5713, wire_5712, wire_5673, wire_5672, wire_5633, wire_5632, wire_5593, wire_5592, wire_3595, wire_3594, wire_3585, wire_3584, wire_3575, wire_3574, wire_3565, wire_3564, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_5479, wire_5478, wire_5469, wire_5468, wire_5459, wire_5458, wire_5449, wire_5448, wire_5383, wire_5382, wire_5343, wire_5342, wire_5303, wire_5302, wire_5263, wire_5262, wire_3239, wire_3238, wire_3229, wire_3228, wire_3219, wire_3218, wire_3209, wire_3208, wire_3133, wire_3132, wire_3093, wire_3092, wire_3053, wire_3052, wire_3013, wire_3012, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_5719, wire_5718, wire_5679, wire_5678, wire_5639, wire_5638, wire_5599, wire_5598, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_3479, wire_3478, wire_3439, wire_3438, wire_3399, wire_3398, wire_3359, wire_3358, wire_5473, wire_5472, wire_5463, wire_5462, wire_5453, wire_5452, wire_5443, wire_5442, wire_5399, wire_5398, wire_5359, wire_5358, wire_5319, wire_5318, wire_5279, wire_5278, wire_3273, wire_3272, wire_3263, wire_3262, wire_3253, wire_3252, wire_3243, wire_3242, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_5799, wire_5798, wire_5789, wire_5788, wire_5779, wire_5778, wire_5769, wire_5768, wire_5689, wire_5688, wire_5649, wire_5648, wire_5609, wire_5608, wire_5569, wire_5568, wire_3599, wire_3598, wire_3589, wire_3588, wire_3579, wire_3578, wire_3569, wire_3568, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_5389, wire_5388, wire_5349, wire_5348, wire_5309, wire_5308, wire_5269, wire_5268, wire_3233, wire_3232, wire_3223, wire_3222, wire_3213, wire_3212, wire_3203, wire_3202, wire_3149, wire_3148, wire_3109, wire_3108, wire_3069, wire_3068, wire_3029, wire_3028, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_5695, wire_5694, wire_5655, wire_5654, wire_5615, wire_5614, wire_5575, wire_5574, wire_3593, wire_3592, wire_3583, wire_3582, wire_3573, wire_3572, wire_3563, wire_3562, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_5477, wire_5476, wire_5467, wire_5466, wire_5457, wire_5456, wire_5447, wire_5446, wire_5375, wire_5374, wire_5335, wire_5334, wire_5295, wire_5294, wire_5255, wire_5254, wire_3277, wire_3276, wire_3267, wire_3266, wire_3257, wire_3256, wire_3247, wire_3246, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_5711, wire_5710, wire_5671, wire_5670, wire_5631, wire_5630, wire_5591, wire_5590, wire_3551, wire_3550, wire_3541, wire_3540, wire_3531, wire_3530, wire_3521, wire_3520, wire_3471, wire_3470, wire_3431, wire_3430, wire_3391, wire_3390, wire_3351, wire_3350, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_5365, wire_5364, wire_5325, wire_5324, wire_5285, wire_5284, wire_5245, wire_5244, wire_3237, wire_3236, wire_3227, wire_3226, wire_3217, wire_3216, wire_3207, wire_3206, wire_3125, wire_3124, wire_3085, wire_3084, wire_3045, wire_3044, wire_3005, wire_3004, wire_5797, wire_5796, wire_5787, wire_5786, wire_5777, wire_5776, wire_5767, wire_5766, wire_5681, wire_5680, wire_5641, wire_5640, wire_5601, wire_5600, wire_5561, wire_5560, wire_3597, wire_3596, wire_3587, wire_3586, wire_3577, wire_3576, wire_3567, wire_3566, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_5391, wire_5390, wire_5351, wire_5350, wire_5311, wire_5310, wire_5271, wire_5270, wire_3231, wire_3230, wire_3221, wire_3220, wire_3211, wire_3210, wire_3201, wire_3200, wire_3141, wire_3140, wire_3101, wire_3100, wire_3061, wire_3060, wire_3021, wire_3020, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_5687, wire_5686, wire_5647, wire_5646, wire_5607, wire_5606, wire_5567, wire_5566, wire_3555, wire_3554, wire_3545, wire_3544, wire_3535, wire_3534, wire_3525, wire_3524, wire_3447, wire_3446, wire_3407, wire_3406, wire_3367, wire_3366, wire_3327, wire_3326, wire_5475, wire_5474, wire_5465, wire_5464, wire_5455, wire_5454, wire_5445, wire_5444, wire_5367, wire_5366, wire_5327, wire_5326, wire_5287, wire_5286, wire_5247, wire_5246, wire_3275, wire_3274, wire_3265, wire_3264, wire_3255, wire_3254, wire_3245, wire_3244, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_5791, wire_5790, wire_5781, wire_5780, wire_5771, wire_5770, wire_5761, wire_5760, wire_5697, wire_5696, wire_5657, wire_5656, wire_5617, wire_5616, wire_5577, wire_5576, wire_3591, wire_3590, wire_3581, wire_3580, wire_3571, wire_3570, wire_3561, wire_3560, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484};
    // IPIN TOTAL: 528
    assign lut_tile_4_4_ipin_in = {wire_3875, wire_3874, wire_3865, wire_3864, wire_3855, wire_3854, wire_3845, wire_3844, wire_3793, wire_3792, wire_3753, wire_3752, wire_3713, wire_3712, wire_3673, wire_3672, wire_5479, wire_5478, wire_5469, wire_5468, wire_5459, wire_5458, wire_5449, wire_5448, wire_5383, wire_5382, wire_5343, wire_5342, wire_5303, wire_5302, wire_5263, wire_5262, wire_3559, wire_3558, wire_3549, wire_3548, wire_3539, wire_3538, wire_3529, wire_3528, wire_3463, wire_3462, wire_3423, wire_3422, wire_3383, wire_3382, wire_3343, wire_3342, wire_5839, wire_5838, wire_5829, wire_5828, wire_5819, wire_5818, wire_5809, wire_5808, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_3919, wire_3918, wire_3909, wire_3908, wire_3899, wire_3898, wire_3889, wire_3888, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_5515, wire_5514, wire_5505, wire_5504, wire_5495, wire_5494, wire_5485, wire_5484, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_3479, wire_3478, wire_3439, wire_3438, wire_3399, wire_3398, wire_3359, wire_3358, wire_5799, wire_5798, wire_5789, wire_5788, wire_5779, wire_5778, wire_5769, wire_5768, wire_5689, wire_5688, wire_5649, wire_5648, wire_5609, wire_5608, wire_5569, wire_5568, wire_3879, wire_3878, wire_3869, wire_3868, wire_3859, wire_3858, wire_3849, wire_3848, wire_3769, wire_3768, wire_3729, wire_3728, wire_3689, wire_3688, wire_3649, wire_3648, wire_5519, wire_5518, wire_5509, wire_5508, wire_5499, wire_5498, wire_5489, wire_5488, wire_5433, wire_5432, wire_5423, wire_5422, wire_5413, wire_5412, wire_5403, wire_5402, wire_3599, wire_3598, wire_3589, wire_3588, wire_3579, wire_3578, wire_3569, wire_3568, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_5833, wire_5832, wire_5823, wire_5822, wire_5813, wire_5812, wire_5803, wire_5802, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_3913, wire_3912, wire_3903, wire_3902, wire_3893, wire_3892, wire_3883, wire_3882, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_5477, wire_5476, wire_5467, wire_5466, wire_5457, wire_5456, wire_5447, wire_5446, wire_5375, wire_5374, wire_5335, wire_5334, wire_5295, wire_5294, wire_5255, wire_5254, wire_3557, wire_3556, wire_3547, wire_3546, wire_3537, wire_3536, wire_3527, wire_3526, wire_3455, wire_3454, wire_3415, wire_3414, wire_3375, wire_3374, wire_3335, wire_3334, wire_5793, wire_5792, wire_5783, wire_5782, wire_5773, wire_5772, wire_5763, wire_5762, wire_5705, wire_5704, wire_5665, wire_5664, wire_5625, wire_5624, wire_5585, wire_5584, wire_3917, wire_3916, wire_3907, wire_3906, wire_3897, wire_3896, wire_3887, wire_3886, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_5513, wire_5512, wire_5503, wire_5502, wire_5493, wire_5492, wire_5483, wire_5482, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_3593, wire_3592, wire_3583, wire_3582, wire_3573, wire_3572, wire_3563, wire_3562, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_5797, wire_5796, wire_5787, wire_5786, wire_5777, wire_5776, wire_5767, wire_5766, wire_5681, wire_5680, wire_5641, wire_5640, wire_5601, wire_5600, wire_5561, wire_5560, wire_3877, wire_3876, wire_3867, wire_3866, wire_3857, wire_3856, wire_3847, wire_3846, wire_3761, wire_3760, wire_3721, wire_3720, wire_3681, wire_3680, wire_3641, wire_3640, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_5391, wire_5390, wire_5351, wire_5350, wire_5311, wire_5310, wire_5271, wire_5270, wire_3551, wire_3550, wire_3541, wire_3540, wire_3531, wire_3530, wire_3521, wire_3520, wire_3471, wire_3470, wire_3431, wire_3430, wire_3391, wire_3390, wire_3351, wire_3350, wire_5831, wire_5830, wire_5821, wire_5820, wire_5811, wire_5810, wire_5801, wire_5800, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_3911, wire_3910, wire_3901, wire_3900, wire_3891, wire_3890, wire_3881, wire_3880, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_5517, wire_5516, wire_5507, wire_5506, wire_5497, wire_5496, wire_5487, wire_5486, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_3555, wire_3554, wire_3545, wire_3544, wire_3535, wire_3534, wire_3525, wire_3524, wire_3447, wire_3446, wire_3407, wire_3406, wire_3367, wire_3366, wire_3327, wire_3326, wire_5791, wire_5790, wire_5781, wire_5780, wire_5771, wire_5770, wire_5761, wire_5760, wire_5697, wire_5696, wire_5657, wire_5656, wire_5617, wire_5616, wire_5577, wire_5576, wire_3871, wire_3870, wire_3861, wire_3860, wire_3851, wire_3850, wire_3841, wire_3840, wire_3777, wire_3776, wire_3737, wire_3736, wire_3697, wire_3696, wire_3657, wire_3656, wire_5511, wire_5510, wire_5501, wire_5500, wire_5491, wire_5490, wire_5481, wire_5480, wire_5435, wire_5434, wire_5425, wire_5424, wire_5415, wire_5414, wire_5405, wire_5404, wire_3591, wire_3590, wire_3581, wire_3580, wire_3571, wire_3570, wire_3561, wire_3560, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_5835, wire_5834, wire_5825, wire_5824, wire_5815, wire_5814, wire_5805, wire_5804, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_3915, wire_3914, wire_3905, wire_3904, wire_3895, wire_3894, wire_3885, wire_3884, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800};
    // IPIN TOTAL: 528
    assign lut_tile_5_4_ipin_in = {wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_4099, wire_4098, wire_4059, wire_4058, wire_4019, wire_4018, wire_3979, wire_3978, wire_5515, wire_5514, wire_5505, wire_5504, wire_5495, wire_5494, wire_5485, wire_5484, wire_5439, wire_5438, wire_5429, wire_5428, wire_5419, wire_5418, wire_5409, wire_5408, wire_3875, wire_3874, wire_3865, wire_3864, wire_3855, wire_3854, wire_3845, wire_3844, wire_3793, wire_3792, wire_3753, wire_3752, wire_3713, wire_3712, wire_3673, wire_3672, wire_5875, wire_5874, wire_5865, wire_5864, wire_5855, wire_5854, wire_5845, wire_5844, wire_5799, wire_5798, wire_5789, wire_5788, wire_5779, wire_5778, wire_5769, wire_5768, wire_4235, wire_4234, wire_4225, wire_4224, wire_4215, wire_4214, wire_4205, wire_4204, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_5559, wire_5558, wire_5549, wire_5548, wire_5539, wire_5538, wire_5529, wire_5528, wire_5475, wire_5474, wire_5465, wire_5464, wire_5455, wire_5454, wire_5445, wire_5444, wire_3879, wire_3878, wire_3869, wire_3868, wire_3859, wire_3858, wire_3849, wire_3848, wire_3769, wire_3768, wire_3729, wire_3728, wire_3689, wire_3688, wire_3649, wire_3648, wire_5833, wire_5832, wire_5823, wire_5822, wire_5813, wire_5812, wire_5803, wire_5802, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_4193, wire_4192, wire_4183, wire_4182, wire_4173, wire_4172, wire_4163, wire_4162, wire_4115, wire_4114, wire_4075, wire_4074, wire_4035, wire_4034, wire_3995, wire_3994, wire_5553, wire_5552, wire_5543, wire_5542, wire_5533, wire_5532, wire_5523, wire_5522, wire_5479, wire_5478, wire_5469, wire_5468, wire_5459, wire_5458, wire_5449, wire_5448, wire_3913, wire_3912, wire_3903, wire_3902, wire_3893, wire_3892, wire_3883, wire_3882, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_5879, wire_5878, wire_5869, wire_5868, wire_5859, wire_5858, wire_5849, wire_5848, wire_5793, wire_5792, wire_5783, wire_5782, wire_5773, wire_5772, wire_5763, wire_5762, wire_4239, wire_4238, wire_4229, wire_4228, wire_4219, wire_4218, wire_4209, wire_4208, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_5513, wire_5512, wire_5503, wire_5502, wire_5493, wire_5492, wire_5483, wire_5482, wire_5437, wire_5436, wire_5427, wire_5426, wire_5417, wire_5416, wire_5407, wire_5406, wire_3873, wire_3872, wire_3863, wire_3862, wire_3853, wire_3852, wire_3843, wire_3842, wire_3785, wire_3784, wire_3745, wire_3744, wire_3705, wire_3704, wire_3665, wire_3664, wire_5837, wire_5836, wire_5827, wire_5826, wire_5817, wire_5816, wire_5807, wire_5806, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_4233, wire_4232, wire_4223, wire_4222, wire_4213, wire_4212, wire_4203, wire_4202, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_5557, wire_5556, wire_5547, wire_5546, wire_5537, wire_5536, wire_5527, wire_5526, wire_5473, wire_5472, wire_5463, wire_5462, wire_5453, wire_5452, wire_5443, wire_5442, wire_3917, wire_3916, wire_3907, wire_3906, wire_3897, wire_3896, wire_3887, wire_3886, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_5831, wire_5830, wire_5821, wire_5820, wire_5811, wire_5810, wire_5801, wire_5800, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_4191, wire_4190, wire_4181, wire_4180, wire_4171, wire_4170, wire_4161, wire_4160, wire_4107, wire_4106, wire_4067, wire_4066, wire_4027, wire_4026, wire_3987, wire_3986, wire_5517, wire_5516, wire_5507, wire_5506, wire_5497, wire_5496, wire_5487, wire_5486, wire_5431, wire_5430, wire_5421, wire_5420, wire_5411, wire_5410, wire_5401, wire_5400, wire_3877, wire_3876, wire_3867, wire_3866, wire_3857, wire_3856, wire_3847, wire_3846, wire_3761, wire_3760, wire_3721, wire_3720, wire_3681, wire_3680, wire_3641, wire_3640, wire_5877, wire_5876, wire_5867, wire_5866, wire_5857, wire_5856, wire_5847, wire_5846, wire_5791, wire_5790, wire_5781, wire_5780, wire_5771, wire_5770, wire_5761, wire_5760, wire_4237, wire_4236, wire_4227, wire_4226, wire_4217, wire_4216, wire_4207, wire_4206, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_5551, wire_5550, wire_5541, wire_5540, wire_5531, wire_5530, wire_5521, wire_5520, wire_5477, wire_5476, wire_5467, wire_5466, wire_5457, wire_5456, wire_5447, wire_5446, wire_3871, wire_3870, wire_3861, wire_3860, wire_3851, wire_3850, wire_3841, wire_3840, wire_3777, wire_3776, wire_3737, wire_3736, wire_3697, wire_3696, wire_3657, wire_3656, wire_5835, wire_5834, wire_5825, wire_5824, wire_5815, wire_5814, wire_5805, wire_5804, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_4083, wire_4082, wire_4043, wire_4042, wire_4003, wire_4002, wire_3963, wire_3962, wire_5555, wire_5554, wire_5545, wire_5544, wire_5535, wire_5534, wire_5525, wire_5524, wire_5471, wire_5470, wire_5461, wire_5460, wire_5451, wire_5450, wire_5441, wire_5440, wire_3915, wire_3914, wire_3905, wire_3904, wire_3895, wire_3894, wire_3885, wire_3884, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_5871, wire_5870, wire_5861, wire_5860, wire_5851, wire_5850, wire_5841, wire_5840, wire_5795, wire_5794, wire_5785, wire_5784, wire_5775, wire_5774, wire_5765, wire_5764, wire_4231, wire_4230, wire_4221, wire_4220, wire_4211, wire_4210, wire_4201, wire_4200, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124};
    // IPIN TOTAL: 528
    assign lut_tile_1_5_ipin_in = {wire_2955, wire_2954, wire_2945, wire_2944, wire_2935, wire_2934, wire_2925, wire_2924, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_5719, wire_5718, wire_5699, wire_5698, wire_5679, wire_5678, wire_5659, wire_5658, wire_5639, wire_5638, wire_5619, wire_5618, wire_5599, wire_5598, wire_5579, wire_5578, wire_2639, wire_2638, wire_2629, wire_2628, wire_2619, wire_2618, wire_2609, wire_2608, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_6035, wire_6034, wire_6023, wire_6022, wire_5995, wire_5994, wire_5983, wire_5982, wire_5955, wire_5954, wire_5943, wire_5942, wire_5915, wire_5914, wire_5903, wire_5902, wire_2999, wire_2998, wire_2989, wire_2988, wire_2979, wire_2978, wire_2969, wire_2968, wire_2915, wire_2914, wire_2905, wire_2904, wire_2895, wire_2894, wire_2885, wire_2884, wire_5717, wire_5716, wire_5697, wire_5696, wire_5677, wire_5676, wire_5657, wire_5656, wire_5637, wire_5636, wire_5617, wire_5616, wire_5597, wire_5596, wire_5577, wire_5576, wire_2633, wire_2632, wire_2623, wire_2622, wire_2613, wire_2612, wire_2603, wire_2602, wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_6033, wire_6032, wire_6013, wire_6012, wire_5993, wire_5992, wire_5973, wire_5972, wire_5953, wire_5952, wire_5933, wire_5932, wire_5913, wire_5912, wire_5893, wire_5892, wire_2959, wire_2958, wire_2949, wire_2948, wire_2939, wire_2938, wire_2929, wire_2928, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_5713, wire_5712, wire_5693, wire_5692, wire_5673, wire_5672, wire_5653, wire_5652, wire_5633, wire_5632, wire_5613, wire_5612, wire_5593, wire_5592, wire_5573, wire_5572, wire_2679, wire_2678, wire_2669, wire_2668, wire_2659, wire_2658, wire_2649, wire_2648, wire_2593, wire_2592, wire_2583, wire_2582, wire_2573, wire_2572, wire_2563, wire_2562, wire_6039, wire_6038, wire_6011, wire_6010, wire_5999, wire_5998, wire_5971, wire_5970, wire_5959, wire_5958, wire_5931, wire_5930, wire_5919, wire_5918, wire_5891, wire_5890, wire_2993, wire_2992, wire_2983, wire_2982, wire_2973, wire_2972, wire_2963, wire_2962, wire_2919, wire_2918, wire_2909, wire_2908, wire_2899, wire_2898, wire_2889, wire_2888, wire_5711, wire_5710, wire_5691, wire_5690, wire_5671, wire_5670, wire_5651, wire_5650, wire_5631, wire_5630, wire_5611, wire_5610, wire_5591, wire_5590, wire_5571, wire_5570, wire_2637, wire_2636, wire_2627, wire_2626, wire_2617, wire_2616, wire_2607, wire_2606, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_6029, wire_6028, wire_6009, wire_6008, wire_5989, wire_5988, wire_5969, wire_5968, wire_5949, wire_5948, wire_5929, wire_5928, wire_5909, wire_5908, wire_5889, wire_5888, wire_2997, wire_2996, wire_2987, wire_2986, wire_2977, wire_2976, wire_2967, wire_2966, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_5709, wire_5708, wire_5689, wire_5688, wire_5669, wire_5668, wire_5649, wire_5648, wire_5629, wire_5628, wire_5609, wire_5608, wire_5589, wire_5588, wire_5569, wire_5568, wire_2673, wire_2672, wire_2663, wire_2662, wire_2653, wire_2652, wire_2643, wire_2642, wire_2597, wire_2596, wire_2587, wire_2586, wire_2577, wire_2576, wire_2567, wire_2566, wire_6025, wire_6024, wire_6005, wire_6004, wire_5985, wire_5984, wire_5965, wire_5964, wire_5945, wire_5944, wire_5925, wire_5924, wire_5905, wire_5904, wire_5885, wire_5884, wire_2957, wire_2956, wire_2947, wire_2946, wire_2937, wire_2936, wire_2927, wire_2926, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_5707, wire_5706, wire_5687, wire_5686, wire_5667, wire_5666, wire_5647, wire_5646, wire_5627, wire_5626, wire_5607, wire_5606, wire_5587, wire_5586, wire_5567, wire_5566, wire_2631, wire_2630, wire_2621, wire_2620, wire_2611, wire_2610, wire_2601, wire_2600, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_6031, wire_6030, wire_6003, wire_6002, wire_5991, wire_5990, wire_5963, wire_5962, wire_5951, wire_5950, wire_5923, wire_5922, wire_5911, wire_5910, wire_5883, wire_5882, wire_2991, wire_2990, wire_2981, wire_2980, wire_2971, wire_2970, wire_2961, wire_2960, wire_2917, wire_2916, wire_2907, wire_2906, wire_2897, wire_2896, wire_2887, wire_2886, wire_5705, wire_5704, wire_5685, wire_5684, wire_5665, wire_5664, wire_5645, wire_5644, wire_5625, wire_5624, wire_5605, wire_5604, wire_5585, wire_5584, wire_5565, wire_5564, wire_2635, wire_2634, wire_2625, wire_2624, wire_2615, wire_2614, wire_2605, wire_2604, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_6021, wire_6020, wire_6001, wire_6000, wire_5981, wire_5980, wire_5961, wire_5960, wire_5941, wire_5940, wire_5921, wire_5920, wire_5901, wire_5900, wire_5881, wire_5880, wire_2951, wire_2950, wire_2941, wire_2940, wire_2931, wire_2930, wire_2921, wire_2920, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_5701, wire_5700, wire_5681, wire_5680, wire_5661, wire_5660, wire_5641, wire_5640, wire_5621, wire_5620, wire_5601, wire_5600, wire_5581, wire_5580, wire_5561, wire_5560, wire_2671, wire_2670, wire_2661, wire_2660, wire_2651, wire_2650, wire_2641, wire_2640, wire_2595, wire_2594, wire_2585, wire_2584, wire_2575, wire_2574, wire_2565, wire_2564, wire_6019, wire_6018, wire_6007, wire_6006, wire_5979, wire_5978, wire_5967, wire_5966, wire_5939, wire_5938, wire_5927, wire_5926, wire_5899, wire_5898, wire_5887, wire_5886, wire_2995, wire_2994, wire_2985, wire_2984, wire_2975, wire_2974, wire_2965, wire_2964, wire_2911, wire_2910, wire_2901, wire_2900, wire_2891, wire_2890, wire_2881, wire_2880};
    // IPIN TOTAL: 528
    assign lut_tile_2_5_ipin_in = {wire_3279, wire_3278, wire_3269, wire_3268, wire_3259, wire_3258, wire_3249, wire_3248, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_5717, wire_5716, wire_5697, wire_5696, wire_5677, wire_5676, wire_5657, wire_5656, wire_5637, wire_5636, wire_5617, wire_5616, wire_5597, wire_5596, wire_5577, wire_5576, wire_2955, wire_2954, wire_2945, wire_2944, wire_2935, wire_2934, wire_2925, wire_2924, wire_2879, wire_2878, wire_2869, wire_2868, wire_2859, wire_2858, wire_2849, wire_2848, wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044, wire_6033, wire_6032, wire_5993, wire_5992, wire_5953, wire_5952, wire_5913, wire_5912, wire_3315, wire_3314, wire_3305, wire_3304, wire_3295, wire_3294, wire_3285, wire_3284, wire_3239, wire_3238, wire_3229, wire_3228, wire_3219, wire_3218, wire_3209, wire_3208, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_5703, wire_5702, wire_5663, wire_5662, wire_5623, wire_5622, wire_5583, wire_5582, wire_2959, wire_2958, wire_2949, wire_2948, wire_2939, wire_2938, wire_2929, wire_2928, wire_2873, wire_2872, wire_2863, wire_2862, wire_2853, wire_2852, wire_2843, wire_2842, wire_6039, wire_6038, wire_6011, wire_6010, wire_5999, wire_5998, wire_5971, wire_5970, wire_5959, wire_5958, wire_5931, wire_5930, wire_5919, wire_5918, wire_5891, wire_5890, wire_3273, wire_3272, wire_3263, wire_3262, wire_3253, wire_3252, wire_3243, wire_3242, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_5719, wire_5718, wire_5679, wire_5678, wire_5639, wire_5638, wire_5599, wire_5598, wire_2993, wire_2992, wire_2983, wire_2982, wire_2973, wire_2972, wire_2963, wire_2962, wire_2919, wire_2918, wire_2909, wire_2908, wire_2899, wire_2898, wire_2889, wire_2888, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_6009, wire_6008, wire_5969, wire_5968, wire_5929, wire_5928, wire_5889, wire_5888, wire_3319, wire_3318, wire_3309, wire_3308, wire_3299, wire_3298, wire_3289, wire_3288, wire_3233, wire_3232, wire_3223, wire_3222, wire_3213, wire_3212, wire_3203, wire_3202, wire_5709, wire_5708, wire_5689, wire_5688, wire_5669, wire_5668, wire_5649, wire_5648, wire_5629, wire_5628, wire_5609, wire_5608, wire_5589, wire_5588, wire_5569, wire_5568, wire_2953, wire_2952, wire_2943, wire_2942, wire_2933, wire_2932, wire_2923, wire_2922, wire_2877, wire_2876, wire_2867, wire_2866, wire_2857, wire_2856, wire_2847, wire_2846, wire_6027, wire_6026, wire_6015, wire_6014, wire_5987, wire_5986, wire_5975, wire_5974, wire_5947, wire_5946, wire_5935, wire_5934, wire_5907, wire_5906, wire_5895, wire_5894, wire_3313, wire_3312, wire_3303, wire_3302, wire_3293, wire_3292, wire_3283, wire_3282, wire_3237, wire_3236, wire_3227, wire_3226, wire_3217, wire_3216, wire_3207, wire_3206, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_5695, wire_5694, wire_5655, wire_5654, wire_5615, wire_5614, wire_5575, wire_5574, wire_2997, wire_2996, wire_2987, wire_2986, wire_2977, wire_2976, wire_2967, wire_2966, wire_2913, wire_2912, wire_2903, wire_2902, wire_2893, wire_2892, wire_2883, wire_2882, wire_6031, wire_6030, wire_6003, wire_6002, wire_5991, wire_5990, wire_5963, wire_5962, wire_5951, wire_5950, wire_5923, wire_5922, wire_5911, wire_5910, wire_5883, wire_5882, wire_3271, wire_3270, wire_3261, wire_3260, wire_3251, wire_3250, wire_3241, wire_3240, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_5705, wire_5704, wire_5685, wire_5684, wire_5665, wire_5664, wire_5645, wire_5644, wire_5625, wire_5624, wire_5605, wire_5604, wire_5585, wire_5584, wire_5565, wire_5564, wire_2957, wire_2956, wire_2947, wire_2946, wire_2937, wire_2936, wire_2927, wire_2926, wire_2871, wire_2870, wire_2861, wire_2860, wire_2851, wire_2850, wire_2841, wire_2840, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6001, wire_6000, wire_5961, wire_5960, wire_5921, wire_5920, wire_5881, wire_5880, wire_3317, wire_3316, wire_3307, wire_3306, wire_3297, wire_3296, wire_3287, wire_3286, wire_3231, wire_3230, wire_3221, wire_3220, wire_3211, wire_3210, wire_3201, wire_3200, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_5711, wire_5710, wire_5671, wire_5670, wire_5631, wire_5630, wire_5591, wire_5590, wire_2951, wire_2950, wire_2941, wire_2940, wire_2931, wire_2930, wire_2921, wire_2920, wire_2875, wire_2874, wire_2865, wire_2864, wire_2855, wire_2854, wire_2845, wire_2844, wire_6019, wire_6018, wire_6007, wire_6006, wire_5979, wire_5978, wire_5967, wire_5966, wire_5939, wire_5938, wire_5927, wire_5926, wire_5899, wire_5898, wire_5887, wire_5886, wire_3275, wire_3274, wire_3265, wire_3264, wire_3255, wire_3254, wire_3245, wire_3244, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_5687, wire_5686, wire_5647, wire_5646, wire_5607, wire_5606, wire_5567, wire_5566, wire_2995, wire_2994, wire_2985, wire_2984, wire_2975, wire_2974, wire_2965, wire_2964, wire_2911, wire_2910, wire_2901, wire_2900, wire_2891, wire_2890, wire_2881, wire_2880, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_6017, wire_6016, wire_5977, wire_5976, wire_5937, wire_5936, wire_5897, wire_5896, wire_3311, wire_3310, wire_3301, wire_3300, wire_3291, wire_3290, wire_3281, wire_3280, wire_3235, wire_3234, wire_3225, wire_3224, wire_3215, wire_3214, wire_3205, wire_3204};
    // IPIN TOTAL: 528
    assign lut_tile_3_5_ipin_in = {wire_3595, wire_3594, wire_3585, wire_3584, wire_3575, wire_3574, wire_3565, wire_3564, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_5703, wire_5702, wire_5663, wire_5662, wire_5623, wire_5622, wire_5583, wire_5582, wire_3279, wire_3278, wire_3269, wire_3268, wire_3259, wire_3258, wire_3249, wire_3248, wire_3195, wire_3194, wire_3185, wire_3184, wire_3175, wire_3174, wire_3165, wire_3164, wire_6119, wire_6118, wire_6109, wire_6108, wire_6099, wire_6098, wire_6089, wire_6088, wire_6019, wire_6018, wire_5979, wire_5978, wire_5939, wire_5938, wire_5899, wire_5898, wire_3639, wire_3638, wire_3629, wire_3628, wire_3619, wire_3618, wire_3609, wire_3608, wire_3555, wire_3554, wire_3545, wire_3544, wire_3535, wire_3534, wire_3525, wire_3524, wire_5795, wire_5794, wire_5785, wire_5784, wire_5775, wire_5774, wire_5765, wire_5764, wire_5713, wire_5712, wire_5673, wire_5672, wire_5633, wire_5632, wire_5593, wire_5592, wire_3273, wire_3272, wire_3263, wire_3262, wire_3253, wire_3252, wire_3243, wire_3242, wire_3199, wire_3198, wire_3189, wire_3188, wire_3179, wire_3178, wire_3169, wire_3168, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_6009, wire_6008, wire_5969, wire_5968, wire_5929, wire_5928, wire_5889, wire_5888, wire_3599, wire_3598, wire_3589, wire_3588, wire_3579, wire_3578, wire_3569, wire_3568, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_5799, wire_5798, wire_5789, wire_5788, wire_5779, wire_5778, wire_5769, wire_5768, wire_5689, wire_5688, wire_5649, wire_5648, wire_5609, wire_5608, wire_5569, wire_5568, wire_3319, wire_3318, wire_3309, wire_3308, wire_3299, wire_3298, wire_3289, wire_3288, wire_3233, wire_3232, wire_3223, wire_3222, wire_3213, wire_3212, wire_3203, wire_3202, wire_6113, wire_6112, wire_6103, wire_6102, wire_6093, wire_6092, wire_6083, wire_6082, wire_6035, wire_6034, wire_5995, wire_5994, wire_5955, wire_5954, wire_5915, wire_5914, wire_3633, wire_3632, wire_3623, wire_3622, wire_3613, wire_3612, wire_3603, wire_3602, wire_3559, wire_3558, wire_3549, wire_3548, wire_3539, wire_3538, wire_3529, wire_3528, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_5695, wire_5694, wire_5655, wire_5654, wire_5615, wire_5614, wire_5575, wire_5574, wire_3277, wire_3276, wire_3267, wire_3266, wire_3257, wire_3256, wire_3247, wire_3246, wire_3193, wire_3192, wire_3183, wire_3182, wire_3173, wire_3172, wire_3163, wire_3162, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_6025, wire_6024, wire_5985, wire_5984, wire_5945, wire_5944, wire_5905, wire_5904, wire_3637, wire_3636, wire_3627, wire_3626, wire_3617, wire_3616, wire_3607, wire_3606, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_5793, wire_5792, wire_5783, wire_5782, wire_5773, wire_5772, wire_5763, wire_5762, wire_5705, wire_5704, wire_5665, wire_5664, wire_5625, wire_5624, wire_5585, wire_5584, wire_3313, wire_3312, wire_3303, wire_3302, wire_3293, wire_3292, wire_3283, wire_3282, wire_3237, wire_3236, wire_3227, wire_3226, wire_3217, wire_3216, wire_3207, wire_3206, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6001, wire_6000, wire_5961, wire_5960, wire_5921, wire_5920, wire_5881, wire_5880, wire_3597, wire_3596, wire_3587, wire_3586, wire_3577, wire_3576, wire_3567, wire_3566, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_5711, wire_5710, wire_5671, wire_5670, wire_5631, wire_5630, wire_5591, wire_5590, wire_3271, wire_3270, wire_3261, wire_3260, wire_3251, wire_3250, wire_3241, wire_3240, wire_3197, wire_3196, wire_3187, wire_3186, wire_3177, wire_3176, wire_3167, wire_3166, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080, wire_6027, wire_6026, wire_5987, wire_5986, wire_5947, wire_5946, wire_5907, wire_5906, wire_3631, wire_3630, wire_3621, wire_3620, wire_3611, wire_3610, wire_3601, wire_3600, wire_3557, wire_3556, wire_3547, wire_3546, wire_3537, wire_3536, wire_3527, wire_3526, wire_5797, wire_5796, wire_5787, wire_5786, wire_5777, wire_5776, wire_5767, wire_5766, wire_5681, wire_5680, wire_5641, wire_5640, wire_5601, wire_5600, wire_5561, wire_5560, wire_3275, wire_3274, wire_3265, wire_3264, wire_3255, wire_3254, wire_3245, wire_3244, wire_3191, wire_3190, wire_3181, wire_3180, wire_3171, wire_3170, wire_3161, wire_3160, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_6017, wire_6016, wire_5977, wire_5976, wire_5937, wire_5936, wire_5897, wire_5896, wire_3591, wire_3590, wire_3581, wire_3580, wire_3571, wire_3570, wire_3561, wire_3560, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_5791, wire_5790, wire_5781, wire_5780, wire_5771, wire_5770, wire_5761, wire_5760, wire_5697, wire_5696, wire_5657, wire_5656, wire_5617, wire_5616, wire_5577, wire_5576, wire_3311, wire_3310, wire_3301, wire_3300, wire_3291, wire_3290, wire_3281, wire_3280, wire_3235, wire_3234, wire_3225, wire_3224, wire_3215, wire_3214, wire_3205, wire_3204, wire_6115, wire_6114, wire_6105, wire_6104, wire_6095, wire_6094, wire_6085, wire_6084, wire_6003, wire_6002, wire_5963, wire_5962, wire_5923, wire_5922, wire_5883, wire_5882, wire_3635, wire_3634, wire_3625, wire_3624, wire_3615, wire_3614, wire_3605, wire_3604, wire_3551, wire_3550, wire_3541, wire_3540, wire_3531, wire_3530, wire_3521, wire_3520};
    // IPIN TOTAL: 528
    assign lut_tile_4_5_ipin_in = {wire_3919, wire_3918, wire_3909, wire_3908, wire_3899, wire_3898, wire_3889, wire_3888, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_5795, wire_5794, wire_5785, wire_5784, wire_5775, wire_5774, wire_5765, wire_5764, wire_5713, wire_5712, wire_5673, wire_5672, wire_5633, wire_5632, wire_5593, wire_5592, wire_3595, wire_3594, wire_3585, wire_3584, wire_3575, wire_3574, wire_3565, wire_3564, wire_3519, wire_3518, wire_3509, wire_3508, wire_3499, wire_3498, wire_3489, wire_3488, wire_6155, wire_6154, wire_6145, wire_6144, wire_6135, wire_6134, wire_6125, wire_6124, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_3955, wire_3954, wire_3945, wire_3944, wire_3935, wire_3934, wire_3925, wire_3924, wire_3879, wire_3878, wire_3869, wire_3868, wire_3859, wire_3858, wire_3849, wire_3848, wire_5839, wire_5838, wire_5829, wire_5828, wire_5819, wire_5818, wire_5809, wire_5808, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_3599, wire_3598, wire_3589, wire_3588, wire_3579, wire_3578, wire_3569, wire_3568, wire_3513, wire_3512, wire_3503, wire_3502, wire_3493, wire_3492, wire_3483, wire_3482, wire_6113, wire_6112, wire_6103, wire_6102, wire_6093, wire_6092, wire_6083, wire_6082, wire_6035, wire_6034, wire_5995, wire_5994, wire_5955, wire_5954, wire_5915, wire_5914, wire_3913, wire_3912, wire_3903, wire_3902, wire_3893, wire_3892, wire_3883, wire_3882, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_5833, wire_5832, wire_5823, wire_5822, wire_5813, wire_5812, wire_5803, wire_5802, wire_5759, wire_5758, wire_5749, wire_5748, wire_5739, wire_5738, wire_5729, wire_5728, wire_3633, wire_3632, wire_3623, wire_3622, wire_3613, wire_3612, wire_3603, wire_3602, wire_3559, wire_3558, wire_3549, wire_3548, wire_3539, wire_3538, wire_3529, wire_3528, wire_6159, wire_6158, wire_6149, wire_6148, wire_6139, wire_6138, wire_6129, wire_6128, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_3959, wire_3958, wire_3949, wire_3948, wire_3939, wire_3938, wire_3929, wire_3928, wire_3873, wire_3872, wire_3863, wire_3862, wire_3853, wire_3852, wire_3843, wire_3842, wire_5793, wire_5792, wire_5783, wire_5782, wire_5773, wire_5772, wire_5763, wire_5762, wire_5705, wire_5704, wire_5665, wire_5664, wire_5625, wire_5624, wire_5585, wire_5584, wire_3593, wire_3592, wire_3583, wire_3582, wire_3573, wire_3572, wire_3563, wire_3562, wire_3517, wire_3516, wire_3507, wire_3506, wire_3497, wire_3496, wire_3487, wire_3486, wire_6117, wire_6116, wire_6107, wire_6106, wire_6097, wire_6096, wire_6087, wire_6086, wire_6011, wire_6010, wire_5971, wire_5970, wire_5931, wire_5930, wire_5891, wire_5890, wire_3953, wire_3952, wire_3943, wire_3942, wire_3933, wire_3932, wire_3923, wire_3922, wire_3877, wire_3876, wire_3867, wire_3866, wire_3857, wire_3856, wire_3847, wire_3846, wire_5837, wire_5836, wire_5827, wire_5826, wire_5817, wire_5816, wire_5807, wire_5806, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_3637, wire_3636, wire_3627, wire_3626, wire_3617, wire_3616, wire_3607, wire_3606, wire_3553, wire_3552, wire_3543, wire_3542, wire_3533, wire_3532, wire_3523, wire_3522, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080, wire_6027, wire_6026, wire_5987, wire_5986, wire_5947, wire_5946, wire_5907, wire_5906, wire_3911, wire_3910, wire_3901, wire_3900, wire_3891, wire_3890, wire_3881, wire_3880, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_5797, wire_5796, wire_5787, wire_5786, wire_5777, wire_5776, wire_5767, wire_5766, wire_5681, wire_5680, wire_5641, wire_5640, wire_5601, wire_5600, wire_5561, wire_5560, wire_3597, wire_3596, wire_3587, wire_3586, wire_3577, wire_3576, wire_3567, wire_3566, wire_3511, wire_3510, wire_3501, wire_3500, wire_3491, wire_3490, wire_3481, wire_3480, wire_6157, wire_6156, wire_6147, wire_6146, wire_6137, wire_6136, wire_6127, wire_6126, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_3957, wire_3956, wire_3947, wire_3946, wire_3937, wire_3936, wire_3927, wire_3926, wire_3871, wire_3870, wire_3861, wire_3860, wire_3851, wire_3850, wire_3841, wire_3840, wire_5831, wire_5830, wire_5821, wire_5820, wire_5811, wire_5810, wire_5801, wire_5800, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_3591, wire_3590, wire_3581, wire_3580, wire_3571, wire_3570, wire_3561, wire_3560, wire_3515, wire_3514, wire_3505, wire_3504, wire_3495, wire_3494, wire_3485, wire_3484, wire_6115, wire_6114, wire_6105, wire_6104, wire_6095, wire_6094, wire_6085, wire_6084, wire_6003, wire_6002, wire_5963, wire_5962, wire_5923, wire_5922, wire_5883, wire_5882, wire_3915, wire_3914, wire_3905, wire_3904, wire_3895, wire_3894, wire_3885, wire_3884, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_5835, wire_5834, wire_5825, wire_5824, wire_5815, wire_5814, wire_5805, wire_5804, wire_5751, wire_5750, wire_5741, wire_5740, wire_5731, wire_5730, wire_5721, wire_5720, wire_3635, wire_3634, wire_3625, wire_3624, wire_3615, wire_3614, wire_3605, wire_3604, wire_3551, wire_3550, wire_3541, wire_3540, wire_3531, wire_3530, wire_3521, wire_3520, wire_6151, wire_6150, wire_6141, wire_6140, wire_6131, wire_6130, wire_6121, wire_6120, wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044, wire_3951, wire_3950, wire_3941, wire_3940, wire_3931, wire_3930, wire_3921, wire_3920, wire_3875, wire_3874, wire_3865, wire_3864, wire_3855, wire_3854, wire_3845, wire_3844};
    // IPIN TOTAL: 528
    assign lut_tile_5_5_ipin_in = {wire_4235, wire_4234, wire_4225, wire_4224, wire_4215, wire_4214, wire_4205, wire_4204, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_5839, wire_5838, wire_5829, wire_5828, wire_5819, wire_5818, wire_5809, wire_5808, wire_5755, wire_5754, wire_5745, wire_5744, wire_5735, wire_5734, wire_5725, wire_5724, wire_3919, wire_3918, wire_3909, wire_3908, wire_3899, wire_3898, wire_3889, wire_3888, wire_3835, wire_3834, wire_3825, wire_3824, wire_3815, wire_3814, wire_3805, wire_3804, wire_6199, wire_6198, wire_6189, wire_6188, wire_6179, wire_6178, wire_6169, wire_6168, wire_6115, wire_6114, wire_6105, wire_6104, wire_6095, wire_6094, wire_6085, wire_6084, wire_4279, wire_4278, wire_4269, wire_4268, wire_4259, wire_4258, wire_4249, wire_4248, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_5875, wire_5874, wire_5865, wire_5864, wire_5855, wire_5854, wire_5845, wire_5844, wire_5799, wire_5798, wire_5789, wire_5788, wire_5779, wire_5778, wire_5769, wire_5768, wire_3913, wire_3912, wire_3903, wire_3902, wire_3893, wire_3892, wire_3883, wire_3882, wire_3839, wire_3838, wire_3829, wire_3828, wire_3819, wire_3818, wire_3809, wire_3808, wire_6159, wire_6158, wire_6149, wire_6148, wire_6139, wire_6138, wire_6129, wire_6128, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_4239, wire_4238, wire_4229, wire_4228, wire_4219, wire_4218, wire_4209, wire_4208, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_5879, wire_5878, wire_5869, wire_5868, wire_5859, wire_5858, wire_5849, wire_5848, wire_5793, wire_5792, wire_5783, wire_5782, wire_5773, wire_5772, wire_5763, wire_5762, wire_3959, wire_3958, wire_3949, wire_3948, wire_3939, wire_3938, wire_3929, wire_3928, wire_3873, wire_3872, wire_3863, wire_3862, wire_3853, wire_3852, wire_3843, wire_3842, wire_6193, wire_6192, wire_6183, wire_6182, wire_6173, wire_6172, wire_6163, wire_6162, wire_6119, wire_6118, wire_6109, wire_6108, wire_6099, wire_6098, wire_6089, wire_6088, wire_4273, wire_4272, wire_4263, wire_4262, wire_4253, wire_4252, wire_4243, wire_4242, wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_5837, wire_5836, wire_5827, wire_5826, wire_5817, wire_5816, wire_5807, wire_5806, wire_5753, wire_5752, wire_5743, wire_5742, wire_5733, wire_5732, wire_5723, wire_5722, wire_3917, wire_3916, wire_3907, wire_3906, wire_3897, wire_3896, wire_3887, wire_3886, wire_3833, wire_3832, wire_3823, wire_3822, wire_3813, wire_3812, wire_3803, wire_3802, wire_6153, wire_6152, wire_6143, wire_6142, wire_6133, wire_6132, wire_6123, wire_6122, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_4277, wire_4276, wire_4267, wire_4266, wire_4257, wire_4256, wire_4247, wire_4246, wire_4193, wire_4192, wire_4183, wire_4182, wire_4173, wire_4172, wire_4163, wire_4162, wire_5873, wire_5872, wire_5863, wire_5862, wire_5853, wire_5852, wire_5843, wire_5842, wire_5797, wire_5796, wire_5787, wire_5786, wire_5777, wire_5776, wire_5767, wire_5766, wire_3953, wire_3952, wire_3943, wire_3942, wire_3933, wire_3932, wire_3923, wire_3922, wire_3877, wire_3876, wire_3867, wire_3866, wire_3857, wire_3856, wire_3847, wire_3846, wire_6157, wire_6156, wire_6147, wire_6146, wire_6137, wire_6136, wire_6127, wire_6126, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_4237, wire_4236, wire_4227, wire_4226, wire_4217, wire_4216, wire_4207, wire_4206, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_5831, wire_5830, wire_5821, wire_5820, wire_5811, wire_5810, wire_5801, wire_5800, wire_5757, wire_5756, wire_5747, wire_5746, wire_5737, wire_5736, wire_5727, wire_5726, wire_3911, wire_3910, wire_3901, wire_3900, wire_3891, wire_3890, wire_3881, wire_3880, wire_3837, wire_3836, wire_3827, wire_3826, wire_3817, wire_3816, wire_3807, wire_3806, wire_6191, wire_6190, wire_6181, wire_6180, wire_6171, wire_6170, wire_6161, wire_6160, wire_6117, wire_6116, wire_6107, wire_6106, wire_6097, wire_6096, wire_6087, wire_6086, wire_4271, wire_4270, wire_4261, wire_4260, wire_4251, wire_4250, wire_4241, wire_4240, wire_4197, wire_4196, wire_4187, wire_4186, wire_4177, wire_4176, wire_4167, wire_4166, wire_5877, wire_5876, wire_5867, wire_5866, wire_5857, wire_5856, wire_5847, wire_5846, wire_5791, wire_5790, wire_5781, wire_5780, wire_5771, wire_5770, wire_5761, wire_5760, wire_3915, wire_3914, wire_3905, wire_3904, wire_3895, wire_3894, wire_3885, wire_3884, wire_3831, wire_3830, wire_3821, wire_3820, wire_3811, wire_3810, wire_3801, wire_3800, wire_6151, wire_6150, wire_6141, wire_6140, wire_6131, wire_6130, wire_6121, wire_6120, wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044, wire_4231, wire_4230, wire_4221, wire_4220, wire_4211, wire_4210, wire_4201, wire_4200, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_5871, wire_5870, wire_5861, wire_5860, wire_5851, wire_5850, wire_5841, wire_5840, wire_5795, wire_5794, wire_5785, wire_5784, wire_5775, wire_5774, wire_5765, wire_5764, wire_3951, wire_3950, wire_3941, wire_3940, wire_3931, wire_3930, wire_3921, wire_3920, wire_3875, wire_3874, wire_3865, wire_3864, wire_3855, wire_3854, wire_3845, wire_3844, wire_6195, wire_6194, wire_6185, wire_6184, wire_6175, wire_6174, wire_6165, wire_6164, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080, wire_4275, wire_4274, wire_4265, wire_4264, wire_4255, wire_4254, wire_4245, wire_4244, wire_4191, wire_4190, wire_4181, wire_4180, wire_4171, wire_4170, wire_4161, wire_4160};
    // IPIN TOTAL: 528


    // FPGA TILE OPIN
    assign wire_333 = lut_tile_1_1_opin_out[0];
    assign wire_334 = lut_tile_1_1_opin_out[1];
    assign wire_335 = lut_tile_1_1_opin_out[2];
    assign wire_336 = lut_tile_1_1_opin_out[3];
    assign wire_337 = lut_tile_1_1_opin_out[4];
    assign wire_338 = lut_tile_1_1_opin_out[5];
    assign wire_339 = lut_tile_1_1_opin_out[6];
    assign wire_340 = lut_tile_1_1_opin_out[7];
    assign wire_341 = lut_tile_1_1_opin_out[8];
    assign wire_342 = lut_tile_1_1_opin_out[9];
    assign wire_709 = lut_tile_1_2_opin_out[0];
    assign wire_710 = lut_tile_1_2_opin_out[1];
    assign wire_711 = lut_tile_1_2_opin_out[2];
    assign wire_712 = lut_tile_1_2_opin_out[3];
    assign wire_713 = lut_tile_1_2_opin_out[4];
    assign wire_714 = lut_tile_1_2_opin_out[5];
    assign wire_715 = lut_tile_1_2_opin_out[6];
    assign wire_716 = lut_tile_1_2_opin_out[7];
    assign wire_717 = lut_tile_1_2_opin_out[8];
    assign wire_718 = lut_tile_1_2_opin_out[9];
    assign wire_1085 = lut_tile_1_3_opin_out[0];
    assign wire_1086 = lut_tile_1_3_opin_out[1];
    assign wire_1087 = lut_tile_1_3_opin_out[2];
    assign wire_1088 = lut_tile_1_3_opin_out[3];
    assign wire_1089 = lut_tile_1_3_opin_out[4];
    assign wire_1090 = lut_tile_1_3_opin_out[5];
    assign wire_1091 = lut_tile_1_3_opin_out[6];
    assign wire_1092 = lut_tile_1_3_opin_out[7];
    assign wire_1093 = lut_tile_1_3_opin_out[8];
    assign wire_1094 = lut_tile_1_3_opin_out[9];
    assign wire_1461 = lut_tile_1_4_opin_out[0];
    assign wire_1462 = lut_tile_1_4_opin_out[1];
    assign wire_1463 = lut_tile_1_4_opin_out[2];
    assign wire_1464 = lut_tile_1_4_opin_out[3];
    assign wire_1465 = lut_tile_1_4_opin_out[4];
    assign wire_1466 = lut_tile_1_4_opin_out[5];
    assign wire_1467 = lut_tile_1_4_opin_out[6];
    assign wire_1468 = lut_tile_1_4_opin_out[7];
    assign wire_1469 = lut_tile_1_4_opin_out[8];
    assign wire_1470 = lut_tile_1_4_opin_out[9];
    assign wire_1837 = lut_tile_1_5_opin_out[0];
    assign wire_1838 = lut_tile_1_5_opin_out[1];
    assign wire_1839 = lut_tile_1_5_opin_out[2];
    assign wire_1840 = lut_tile_1_5_opin_out[3];
    assign wire_1841 = lut_tile_1_5_opin_out[4];
    assign wire_1842 = lut_tile_1_5_opin_out[5];
    assign wire_1843 = lut_tile_1_5_opin_out[6];
    assign wire_1844 = lut_tile_1_5_opin_out[7];
    assign wire_1845 = lut_tile_1_5_opin_out[8];
    assign wire_1846 = lut_tile_1_5_opin_out[9];
    assign wire_389 = lut_tile_2_1_opin_out[0];
    assign wire_390 = lut_tile_2_1_opin_out[1];
    assign wire_391 = lut_tile_2_1_opin_out[2];
    assign wire_392 = lut_tile_2_1_opin_out[3];
    assign wire_393 = lut_tile_2_1_opin_out[4];
    assign wire_394 = lut_tile_2_1_opin_out[5];
    assign wire_395 = lut_tile_2_1_opin_out[6];
    assign wire_396 = lut_tile_2_1_opin_out[7];
    assign wire_397 = lut_tile_2_1_opin_out[8];
    assign wire_398 = lut_tile_2_1_opin_out[9];
    assign wire_765 = lut_tile_2_2_opin_out[0];
    assign wire_766 = lut_tile_2_2_opin_out[1];
    assign wire_767 = lut_tile_2_2_opin_out[2];
    assign wire_768 = lut_tile_2_2_opin_out[3];
    assign wire_769 = lut_tile_2_2_opin_out[4];
    assign wire_770 = lut_tile_2_2_opin_out[5];
    assign wire_771 = lut_tile_2_2_opin_out[6];
    assign wire_772 = lut_tile_2_2_opin_out[7];
    assign wire_773 = lut_tile_2_2_opin_out[8];
    assign wire_774 = lut_tile_2_2_opin_out[9];
    assign wire_1141 = lut_tile_2_3_opin_out[0];
    assign wire_1142 = lut_tile_2_3_opin_out[1];
    assign wire_1143 = lut_tile_2_3_opin_out[2];
    assign wire_1144 = lut_tile_2_3_opin_out[3];
    assign wire_1145 = lut_tile_2_3_opin_out[4];
    assign wire_1146 = lut_tile_2_3_opin_out[5];
    assign wire_1147 = lut_tile_2_3_opin_out[6];
    assign wire_1148 = lut_tile_2_3_opin_out[7];
    assign wire_1149 = lut_tile_2_3_opin_out[8];
    assign wire_1150 = lut_tile_2_3_opin_out[9];
    assign wire_1517 = lut_tile_2_4_opin_out[0];
    assign wire_1518 = lut_tile_2_4_opin_out[1];
    assign wire_1519 = lut_tile_2_4_opin_out[2];
    assign wire_1520 = lut_tile_2_4_opin_out[3];
    assign wire_1521 = lut_tile_2_4_opin_out[4];
    assign wire_1522 = lut_tile_2_4_opin_out[5];
    assign wire_1523 = lut_tile_2_4_opin_out[6];
    assign wire_1524 = lut_tile_2_4_opin_out[7];
    assign wire_1525 = lut_tile_2_4_opin_out[8];
    assign wire_1526 = lut_tile_2_4_opin_out[9];
    assign wire_1893 = lut_tile_2_5_opin_out[0];
    assign wire_1894 = lut_tile_2_5_opin_out[1];
    assign wire_1895 = lut_tile_2_5_opin_out[2];
    assign wire_1896 = lut_tile_2_5_opin_out[3];
    assign wire_1897 = lut_tile_2_5_opin_out[4];
    assign wire_1898 = lut_tile_2_5_opin_out[5];
    assign wire_1899 = lut_tile_2_5_opin_out[6];
    assign wire_1900 = lut_tile_2_5_opin_out[7];
    assign wire_1901 = lut_tile_2_5_opin_out[8];
    assign wire_1902 = lut_tile_2_5_opin_out[9];
    assign wire_445 = lut_tile_3_1_opin_out[0];
    assign wire_446 = lut_tile_3_1_opin_out[1];
    assign wire_447 = lut_tile_3_1_opin_out[2];
    assign wire_448 = lut_tile_3_1_opin_out[3];
    assign wire_449 = lut_tile_3_1_opin_out[4];
    assign wire_450 = lut_tile_3_1_opin_out[5];
    assign wire_451 = lut_tile_3_1_opin_out[6];
    assign wire_452 = lut_tile_3_1_opin_out[7];
    assign wire_453 = lut_tile_3_1_opin_out[8];
    assign wire_454 = lut_tile_3_1_opin_out[9];
    assign wire_821 = lut_tile_3_2_opin_out[0];
    assign wire_822 = lut_tile_3_2_opin_out[1];
    assign wire_823 = lut_tile_3_2_opin_out[2];
    assign wire_824 = lut_tile_3_2_opin_out[3];
    assign wire_825 = lut_tile_3_2_opin_out[4];
    assign wire_826 = lut_tile_3_2_opin_out[5];
    assign wire_827 = lut_tile_3_2_opin_out[6];
    assign wire_828 = lut_tile_3_2_opin_out[7];
    assign wire_829 = lut_tile_3_2_opin_out[8];
    assign wire_830 = lut_tile_3_2_opin_out[9];
    assign wire_1197 = lut_tile_3_3_opin_out[0];
    assign wire_1198 = lut_tile_3_3_opin_out[1];
    assign wire_1199 = lut_tile_3_3_opin_out[2];
    assign wire_1200 = lut_tile_3_3_opin_out[3];
    assign wire_1201 = lut_tile_3_3_opin_out[4];
    assign wire_1202 = lut_tile_3_3_opin_out[5];
    assign wire_1203 = lut_tile_3_3_opin_out[6];
    assign wire_1204 = lut_tile_3_3_opin_out[7];
    assign wire_1205 = lut_tile_3_3_opin_out[8];
    assign wire_1206 = lut_tile_3_3_opin_out[9];
    assign wire_1573 = lut_tile_3_4_opin_out[0];
    assign wire_1574 = lut_tile_3_4_opin_out[1];
    assign wire_1575 = lut_tile_3_4_opin_out[2];
    assign wire_1576 = lut_tile_3_4_opin_out[3];
    assign wire_1577 = lut_tile_3_4_opin_out[4];
    assign wire_1578 = lut_tile_3_4_opin_out[5];
    assign wire_1579 = lut_tile_3_4_opin_out[6];
    assign wire_1580 = lut_tile_3_4_opin_out[7];
    assign wire_1581 = lut_tile_3_4_opin_out[8];
    assign wire_1582 = lut_tile_3_4_opin_out[9];
    assign wire_1949 = lut_tile_3_5_opin_out[0];
    assign wire_1950 = lut_tile_3_5_opin_out[1];
    assign wire_1951 = lut_tile_3_5_opin_out[2];
    assign wire_1952 = lut_tile_3_5_opin_out[3];
    assign wire_1953 = lut_tile_3_5_opin_out[4];
    assign wire_1954 = lut_tile_3_5_opin_out[5];
    assign wire_1955 = lut_tile_3_5_opin_out[6];
    assign wire_1956 = lut_tile_3_5_opin_out[7];
    assign wire_1957 = lut_tile_3_5_opin_out[8];
    assign wire_1958 = lut_tile_3_5_opin_out[9];
    assign wire_501 = lut_tile_4_1_opin_out[0];
    assign wire_502 = lut_tile_4_1_opin_out[1];
    assign wire_503 = lut_tile_4_1_opin_out[2];
    assign wire_504 = lut_tile_4_1_opin_out[3];
    assign wire_505 = lut_tile_4_1_opin_out[4];
    assign wire_506 = lut_tile_4_1_opin_out[5];
    assign wire_507 = lut_tile_4_1_opin_out[6];
    assign wire_508 = lut_tile_4_1_opin_out[7];
    assign wire_509 = lut_tile_4_1_opin_out[8];
    assign wire_510 = lut_tile_4_1_opin_out[9];
    assign wire_877 = lut_tile_4_2_opin_out[0];
    assign wire_878 = lut_tile_4_2_opin_out[1];
    assign wire_879 = lut_tile_4_2_opin_out[2];
    assign wire_880 = lut_tile_4_2_opin_out[3];
    assign wire_881 = lut_tile_4_2_opin_out[4];
    assign wire_882 = lut_tile_4_2_opin_out[5];
    assign wire_883 = lut_tile_4_2_opin_out[6];
    assign wire_884 = lut_tile_4_2_opin_out[7];
    assign wire_885 = lut_tile_4_2_opin_out[8];
    assign wire_886 = lut_tile_4_2_opin_out[9];
    assign wire_1253 = lut_tile_4_3_opin_out[0];
    assign wire_1254 = lut_tile_4_3_opin_out[1];
    assign wire_1255 = lut_tile_4_3_opin_out[2];
    assign wire_1256 = lut_tile_4_3_opin_out[3];
    assign wire_1257 = lut_tile_4_3_opin_out[4];
    assign wire_1258 = lut_tile_4_3_opin_out[5];
    assign wire_1259 = lut_tile_4_3_opin_out[6];
    assign wire_1260 = lut_tile_4_3_opin_out[7];
    assign wire_1261 = lut_tile_4_3_opin_out[8];
    assign wire_1262 = lut_tile_4_3_opin_out[9];
    assign wire_1629 = lut_tile_4_4_opin_out[0];
    assign wire_1630 = lut_tile_4_4_opin_out[1];
    assign wire_1631 = lut_tile_4_4_opin_out[2];
    assign wire_1632 = lut_tile_4_4_opin_out[3];
    assign wire_1633 = lut_tile_4_4_opin_out[4];
    assign wire_1634 = lut_tile_4_4_opin_out[5];
    assign wire_1635 = lut_tile_4_4_opin_out[6];
    assign wire_1636 = lut_tile_4_4_opin_out[7];
    assign wire_1637 = lut_tile_4_4_opin_out[8];
    assign wire_1638 = lut_tile_4_4_opin_out[9];
    assign wire_2005 = lut_tile_4_5_opin_out[0];
    assign wire_2006 = lut_tile_4_5_opin_out[1];
    assign wire_2007 = lut_tile_4_5_opin_out[2];
    assign wire_2008 = lut_tile_4_5_opin_out[3];
    assign wire_2009 = lut_tile_4_5_opin_out[4];
    assign wire_2010 = lut_tile_4_5_opin_out[5];
    assign wire_2011 = lut_tile_4_5_opin_out[6];
    assign wire_2012 = lut_tile_4_5_opin_out[7];
    assign wire_2013 = lut_tile_4_5_opin_out[8];
    assign wire_2014 = lut_tile_4_5_opin_out[9];
    assign wire_557 = lut_tile_5_1_opin_out[0];
    assign wire_558 = lut_tile_5_1_opin_out[1];
    assign wire_559 = lut_tile_5_1_opin_out[2];
    assign wire_560 = lut_tile_5_1_opin_out[3];
    assign wire_561 = lut_tile_5_1_opin_out[4];
    assign wire_562 = lut_tile_5_1_opin_out[5];
    assign wire_563 = lut_tile_5_1_opin_out[6];
    assign wire_564 = lut_tile_5_1_opin_out[7];
    assign wire_565 = lut_tile_5_1_opin_out[8];
    assign wire_566 = lut_tile_5_1_opin_out[9];
    assign wire_933 = lut_tile_5_2_opin_out[0];
    assign wire_934 = lut_tile_5_2_opin_out[1];
    assign wire_935 = lut_tile_5_2_opin_out[2];
    assign wire_936 = lut_tile_5_2_opin_out[3];
    assign wire_937 = lut_tile_5_2_opin_out[4];
    assign wire_938 = lut_tile_5_2_opin_out[5];
    assign wire_939 = lut_tile_5_2_opin_out[6];
    assign wire_940 = lut_tile_5_2_opin_out[7];
    assign wire_941 = lut_tile_5_2_opin_out[8];
    assign wire_942 = lut_tile_5_2_opin_out[9];
    assign wire_1309 = lut_tile_5_3_opin_out[0];
    assign wire_1310 = lut_tile_5_3_opin_out[1];
    assign wire_1311 = lut_tile_5_3_opin_out[2];
    assign wire_1312 = lut_tile_5_3_opin_out[3];
    assign wire_1313 = lut_tile_5_3_opin_out[4];
    assign wire_1314 = lut_tile_5_3_opin_out[5];
    assign wire_1315 = lut_tile_5_3_opin_out[6];
    assign wire_1316 = lut_tile_5_3_opin_out[7];
    assign wire_1317 = lut_tile_5_3_opin_out[8];
    assign wire_1318 = lut_tile_5_3_opin_out[9];
    assign wire_1685 = lut_tile_5_4_opin_out[0];
    assign wire_1686 = lut_tile_5_4_opin_out[1];
    assign wire_1687 = lut_tile_5_4_opin_out[2];
    assign wire_1688 = lut_tile_5_4_opin_out[3];
    assign wire_1689 = lut_tile_5_4_opin_out[4];
    assign wire_1690 = lut_tile_5_4_opin_out[5];
    assign wire_1691 = lut_tile_5_4_opin_out[6];
    assign wire_1692 = lut_tile_5_4_opin_out[7];
    assign wire_1693 = lut_tile_5_4_opin_out[8];
    assign wire_1694 = lut_tile_5_4_opin_out[9];
    assign wire_2061 = lut_tile_5_5_opin_out[0];
    assign wire_2062 = lut_tile_5_5_opin_out[1];
    assign wire_2063 = lut_tile_5_5_opin_out[2];
    assign wire_2064 = lut_tile_5_5_opin_out[3];
    assign wire_2065 = lut_tile_5_5_opin_out[4];
    assign wire_2066 = lut_tile_5_5_opin_out[5];
    assign wire_2067 = lut_tile_5_5_opin_out[6];
    assign wire_2068 = lut_tile_5_5_opin_out[7];
    assign wire_2069 = lut_tile_5_5_opin_out[8];
    assign wire_2070 = lut_tile_5_5_opin_out[9];
    // LUT TILE CHANXY 
    assign lut_tile_1_1_chanxy_in = {wire_2519, wire_2518, wire_4799, wire_2879, wire_2839, wire_2838, wire_2785, wire_2784, wire_2731, wire_2730, wire_2684, wire_715, wire_341, wire_2517, wire_2516, wire_2539, wire_2434, wire_2559, wire_2514, wire_2513, wire_2512, wire_4797, wire_2841, wire_2836, wire_2835, wire_2834, wire_2783, wire_2782, wire_2729, wire_2728, wire_715, wire_341, wire_2433, wire_2432, wire_2511, wire_2510, wire_2509, wire_2508, wire_2557, wire_2506, wire_4795, wire_2843, wire_2833, wire_2832, wire_2828, wire_2779, wire_2778, wire_2727, wire_2726, wire_715, wire_341, wire_2431, wire_2430, wire_2429, wire_2428, wire_2505, wire_2504, wire_2537, wire_2426, wire_4793, wire_2845, wire_2831, wire_2830, wire_2820, wire_2777, wire_2776, wire_2723, wire_2722, wire_715, wire_341, wire_2425, wire_2424, wire_2503, wire_2502, wire_2423, wire_2422, wire_2421, wire_2420, wire_4791, wire_2847, wire_2827, wire_2826, wire_2812, wire_2775, wire_2774, wire_2721, wire_2720, wire_715, wire_337, wire_2501, wire_2500, wire_2535, wire_2418, wire_2417, wire_2416, wire_2415, wire_2414, wire_4789, wire_2849, wire_2825, wire_2824, wire_2804, wire_2771, wire_2770, wire_2719, wire_2718, wire_715, wire_337, wire_2555, wire_2498, wire_2497, wire_2496, wire_2413, wire_2412, wire_2495, wire_2494, wire_4787, wire_2851, wire_2823, wire_2822, wire_2796, wire_2769, wire_2768, wire_2715, wire_2714, wire_715, wire_337, wire_2493, wire_2492, wire_2533, wire_2410, wire_2553, wire_2490, wire_2489, wire_2488, wire_4785, wire_2853, wire_2819, wire_2818, wire_2788, wire_2767, wire_2766, wire_2713, wire_2712, wire_715, wire_337, wire_2409, wire_2408, wire_2487, wire_2486, wire_2485, wire_2484, wire_2551, wire_2482, wire_4783, wire_2855, wire_2817, wire_2816, wire_2780, wire_2763, wire_2762, wire_2711, wire_2710, wire_711, wire_337, wire_2407, wire_2406, wire_2405, wire_2404, wire_2481, wire_2480, wire_2531, wire_2402, wire_4781, wire_2857, wire_2815, wire_2814, wire_2772, wire_2761, wire_2760, wire_2707, wire_2706, wire_711, wire_337, wire_2401, wire_2400, wire_2479, wire_2478, wire_2399, wire_2398, wire_2397, wire_2396, wire_715, wire_4779, wire_2859, wire_2811, wire_2810, wire_2764, wire_2759, wire_2758, wire_2705, wire_2704, wire_711, wire_337, wire_2477, wire_2476, wire_715, wire_2529, wire_2394, wire_715, wire_2393, wire_2392, wire_715, wire_2391, wire_2390, wire_715, wire_4777, wire_2861, wire_2809, wire_2808, wire_2756, wire_2755, wire_2754, wire_2703, wire_2702, wire_711, wire_337, wire_2549, wire_2474, wire_715, wire_2473, wire_2472, wire_715, wire_2389, wire_2388, wire_715, wire_2471, wire_2470, wire_711, wire_4775, wire_2863, wire_2807, wire_2806, wire_2753, wire_2752, wire_2748, wire_2699, wire_2698, wire_711, wire_333, wire_2469, wire_2468, wire_711, wire_2527, wire_2386, wire_711, wire_2547, wire_2466, wire_711, wire_2465, wire_2464, wire_711, wire_4773, wire_2865, wire_2803, wire_2802, wire_2751, wire_2750, wire_2740, wire_2697, wire_2696, wire_711, wire_333, wire_2385, wire_2384, wire_711, wire_2463, wire_2462, wire_711, wire_2461, wire_2460, wire_711, wire_2545, wire_2458, wire_341, wire_4771, wire_2867, wire_2801, wire_2800, wire_2747, wire_2746, wire_2732, wire_2695, wire_2694, wire_711, wire_333, wire_2383, wire_2382, wire_341, wire_2381, wire_2380, wire_341, wire_2457, wire_2456, wire_341, wire_2525, wire_2378, wire_341, wire_4769, wire_2869, wire_2799, wire_2798, wire_2745, wire_2744, wire_2724, wire_2691, wire_2690, wire_711, wire_333, wire_2377, wire_2376, wire_341, wire_2455, wire_2454, wire_341, wire_2375, wire_2374, wire_341, wire_2373, wire_2372, wire_337, wire_4767, wire_2871, wire_2795, wire_2794, wire_2743, wire_2742, wire_2716, wire_2689, wire_2688, wire_341, wire_333, wire_2453, wire_2452, wire_337, wire_2523, wire_2370, wire_337, wire_2369, wire_2368, wire_337, wire_2367, wire_2366, wire_337, wire_4765, wire_2873, wire_2793, wire_2792, wire_2739, wire_2738, wire_2708, wire_2687, wire_2686, wire_341, wire_333, wire_2543, wire_2450, wire_337, wire_2449, wire_2448, wire_337, wire_2365, wire_2364, wire_337, wire_2447, wire_2446, wire_333, wire_4763, wire_2875, wire_2791, wire_2790, wire_2737, wire_2736, wire_2700, wire_2683, wire_2682, wire_341, wire_333, wire_2445, wire_2444, wire_333, wire_2521, wire_2362, wire_333, wire_2541, wire_2442, wire_333, wire_2441, wire_2440, wire_333, wire_4761, wire_2877, wire_2787, wire_2786, wire_2735, wire_2734, wire_2692, wire_2681, wire_2680, wire_341, wire_333, wire_2361, wire_2360, wire_333, wire_2439, wire_2438, wire_333, wire_2437, wire_2436, wire_333, wire_4439, wire_4438, wire_4763, wire_4759, wire_4758, wire_4748, wire_4705, wire_4704, wire_4651, wire_4650, wire_2879, wire_398, wire_390, wire_4437, wire_4436, wire_4459, wire_4354, wire_4479, wire_4434, wire_4433, wire_4432, wire_4765, wire_4755, wire_4754, wire_4740, wire_4703, wire_4702, wire_4649, wire_4648, wire_2877, wire_398, wire_390, wire_4353, wire_4352, wire_4431, wire_4430, wire_4429, wire_4428, wire_4477, wire_4426, wire_4767, wire_4753, wire_4752, wire_4732, wire_4699, wire_4698, wire_4647, wire_4646, wire_2875, wire_398, wire_390, wire_4351, wire_4350, wire_4349, wire_4348, wire_4425, wire_4424, wire_4457, wire_4346, wire_4769, wire_4751, wire_4750, wire_4724, wire_4697, wire_4696, wire_4643, wire_4642, wire_2873, wire_398, wire_390, wire_4345, wire_4344, wire_4423, wire_4422, wire_4343, wire_4342, wire_4341, wire_4340, wire_4771, wire_4747, wire_4746, wire_4716, wire_4695, wire_4694, wire_4641, wire_4640, wire_2871, wire_398, wire_340, wire_4421, wire_4420, wire_4455, wire_4338, wire_4337, wire_4336, wire_4335, wire_4334, wire_4773, wire_4745, wire_4744, wire_4708, wire_4691, wire_4690, wire_4639, wire_4638, wire_2869, wire_398, wire_340, wire_4475, wire_4418, wire_4417, wire_4416, wire_4333, wire_4332, wire_4415, wire_4414, wire_4775, wire_4743, wire_4742, wire_4700, wire_4689, wire_4688, wire_4635, wire_4634, wire_2867, wire_398, wire_340, wire_4413, wire_4412, wire_4453, wire_4330, wire_4473, wire_4410, wire_4409, wire_4408, wire_4777, wire_4739, wire_4738, wire_4692, wire_4687, wire_4686, wire_4633, wire_4632, wire_2865, wire_398, wire_340, wire_4329, wire_4328, wire_4407, wire_4406, wire_4405, wire_4404, wire_4471, wire_4402, wire_4779, wire_4737, wire_4736, wire_4684, wire_4683, wire_4682, wire_4631, wire_4630, wire_2863, wire_394, wire_340, wire_4327, wire_4326, wire_4325, wire_4324, wire_4401, wire_4400, wire_4451, wire_4322, wire_4781, wire_4735, wire_4734, wire_4681, wire_4680, wire_4676, wire_4627, wire_4626, wire_2861, wire_394, wire_340, wire_4321, wire_4320, wire_4399, wire_4398, wire_4319, wire_4318, wire_4317, wire_4316, wire_398, wire_4783, wire_4731, wire_4730, wire_4679, wire_4678, wire_4668, wire_4625, wire_4624, wire_2859, wire_394, wire_340, wire_4397, wire_4396, wire_398, wire_4449, wire_4314, wire_398, wire_4313, wire_4312, wire_398, wire_4311, wire_4310, wire_398, wire_4785, wire_4729, wire_4728, wire_4675, wire_4674, wire_4660, wire_4623, wire_4622, wire_2857, wire_394, wire_340, wire_4469, wire_4394, wire_398, wire_4393, wire_4392, wire_398, wire_4309, wire_4308, wire_398, wire_4391, wire_4390, wire_394, wire_4787, wire_4727, wire_4726, wire_4673, wire_4672, wire_4652, wire_4619, wire_4618, wire_2855, wire_394, wire_336, wire_4389, wire_4388, wire_394, wire_4447, wire_4306, wire_394, wire_4467, wire_4386, wire_394, wire_4385, wire_4384, wire_394, wire_4789, wire_4723, wire_4722, wire_4671, wire_4670, wire_4644, wire_4617, wire_4616, wire_2853, wire_394, wire_336, wire_4305, wire_4304, wire_394, wire_4383, wire_4382, wire_394, wire_4381, wire_4380, wire_394, wire_4465, wire_4378, wire_390, wire_4791, wire_4721, wire_4720, wire_4667, wire_4666, wire_4636, wire_4615, wire_4614, wire_2851, wire_394, wire_336, wire_4303, wire_4302, wire_390, wire_4301, wire_4300, wire_390, wire_4377, wire_4376, wire_390, wire_4445, wire_4298, wire_390, wire_4793, wire_4719, wire_4718, wire_4665, wire_4664, wire_4628, wire_4611, wire_4610, wire_2849, wire_394, wire_336, wire_4297, wire_4296, wire_390, wire_4375, wire_4374, wire_390, wire_4295, wire_4294, wire_390, wire_4293, wire_4292, wire_340, wire_4795, wire_4715, wire_4714, wire_4663, wire_4662, wire_4620, wire_4609, wire_4608, wire_2847, wire_390, wire_336, wire_4373, wire_4372, wire_340, wire_4443, wire_4290, wire_340, wire_4289, wire_4288, wire_340, wire_4287, wire_4286, wire_340, wire_4797, wire_4713, wire_4712, wire_4659, wire_4658, wire_4612, wire_4607, wire_4606, wire_2845, wire_390, wire_336, wire_4463, wire_4370, wire_340, wire_4369, wire_4368, wire_340, wire_4285, wire_4284, wire_340, wire_4367, wire_4366, wire_336, wire_4799, wire_4711, wire_4710, wire_4657, wire_4656, wire_4604, wire_4603, wire_4602, wire_2843, wire_390, wire_336, wire_4365, wire_4364, wire_336, wire_4441, wire_4282, wire_336, wire_4461, wire_4362, wire_336, wire_4361, wire_4360, wire_336, wire_4761, wire_4756, wire_4707, wire_4706, wire_4655, wire_4654, wire_4601, wire_4600, wire_2841, wire_390, wire_336, wire_4281, wire_4280, wire_336, wire_4359, wire_4358, wire_336, wire_4357, wire_4356, wire_336};
    // CHNAXY TOTAL: 840
    assign wire_2680 = lut_tile_1_1_chanxy_out[0];
    assign wire_2682 = lut_tile_1_1_chanxy_out[1];
    assign wire_2684 = lut_tile_1_1_chanxy_out[2];
    assign wire_2685 = lut_tile_1_1_chanxy_out[3];
    assign wire_2686 = lut_tile_1_1_chanxy_out[4];
    assign wire_2688 = lut_tile_1_1_chanxy_out[5];
    assign wire_2690 = lut_tile_1_1_chanxy_out[6];
    assign wire_2692 = lut_tile_1_1_chanxy_out[7];
    assign wire_2693 = lut_tile_1_1_chanxy_out[8];
    assign wire_2694 = lut_tile_1_1_chanxy_out[9];
    assign wire_2696 = lut_tile_1_1_chanxy_out[10];
    assign wire_2698 = lut_tile_1_1_chanxy_out[11];
    assign wire_2700 = lut_tile_1_1_chanxy_out[12];
    assign wire_2701 = lut_tile_1_1_chanxy_out[13];
    assign wire_2702 = lut_tile_1_1_chanxy_out[14];
    assign wire_2704 = lut_tile_1_1_chanxy_out[15];
    assign wire_2706 = lut_tile_1_1_chanxy_out[16];
    assign wire_2708 = lut_tile_1_1_chanxy_out[17];
    assign wire_2709 = lut_tile_1_1_chanxy_out[18];
    assign wire_2710 = lut_tile_1_1_chanxy_out[19];
    assign wire_2712 = lut_tile_1_1_chanxy_out[20];
    assign wire_2714 = lut_tile_1_1_chanxy_out[21];
    assign wire_2716 = lut_tile_1_1_chanxy_out[22];
    assign wire_2717 = lut_tile_1_1_chanxy_out[23];
    assign wire_2718 = lut_tile_1_1_chanxy_out[24];
    assign wire_2720 = lut_tile_1_1_chanxy_out[25];
    assign wire_2722 = lut_tile_1_1_chanxy_out[26];
    assign wire_2724 = lut_tile_1_1_chanxy_out[27];
    assign wire_2725 = lut_tile_1_1_chanxy_out[28];
    assign wire_2726 = lut_tile_1_1_chanxy_out[29];
    assign wire_2728 = lut_tile_1_1_chanxy_out[30];
    assign wire_2730 = lut_tile_1_1_chanxy_out[31];
    assign wire_2732 = lut_tile_1_1_chanxy_out[32];
    assign wire_2733 = lut_tile_1_1_chanxy_out[33];
    assign wire_2734 = lut_tile_1_1_chanxy_out[34];
    assign wire_2736 = lut_tile_1_1_chanxy_out[35];
    assign wire_2738 = lut_tile_1_1_chanxy_out[36];
    assign wire_2740 = lut_tile_1_1_chanxy_out[37];
    assign wire_2741 = lut_tile_1_1_chanxy_out[38];
    assign wire_2742 = lut_tile_1_1_chanxy_out[39];
    assign wire_2744 = lut_tile_1_1_chanxy_out[40];
    assign wire_2746 = lut_tile_1_1_chanxy_out[41];
    assign wire_2748 = lut_tile_1_1_chanxy_out[42];
    assign wire_2749 = lut_tile_1_1_chanxy_out[43];
    assign wire_2750 = lut_tile_1_1_chanxy_out[44];
    assign wire_2752 = lut_tile_1_1_chanxy_out[45];
    assign wire_2754 = lut_tile_1_1_chanxy_out[46];
    assign wire_2756 = lut_tile_1_1_chanxy_out[47];
    assign wire_2757 = lut_tile_1_1_chanxy_out[48];
    assign wire_2758 = lut_tile_1_1_chanxy_out[49];
    assign wire_2760 = lut_tile_1_1_chanxy_out[50];
    assign wire_2762 = lut_tile_1_1_chanxy_out[51];
    assign wire_2764 = lut_tile_1_1_chanxy_out[52];
    assign wire_2765 = lut_tile_1_1_chanxy_out[53];
    assign wire_2766 = lut_tile_1_1_chanxy_out[54];
    assign wire_2768 = lut_tile_1_1_chanxy_out[55];
    assign wire_2770 = lut_tile_1_1_chanxy_out[56];
    assign wire_2772 = lut_tile_1_1_chanxy_out[57];
    assign wire_2773 = lut_tile_1_1_chanxy_out[58];
    assign wire_2774 = lut_tile_1_1_chanxy_out[59];
    assign wire_2776 = lut_tile_1_1_chanxy_out[60];
    assign wire_2778 = lut_tile_1_1_chanxy_out[61];
    assign wire_2780 = lut_tile_1_1_chanxy_out[62];
    assign wire_2781 = lut_tile_1_1_chanxy_out[63];
    assign wire_2782 = lut_tile_1_1_chanxy_out[64];
    assign wire_2784 = lut_tile_1_1_chanxy_out[65];
    assign wire_2786 = lut_tile_1_1_chanxy_out[66];
    assign wire_2788 = lut_tile_1_1_chanxy_out[67];
    assign wire_2789 = lut_tile_1_1_chanxy_out[68];
    assign wire_2790 = lut_tile_1_1_chanxy_out[69];
    assign wire_2792 = lut_tile_1_1_chanxy_out[70];
    assign wire_2794 = lut_tile_1_1_chanxy_out[71];
    assign wire_2796 = lut_tile_1_1_chanxy_out[72];
    assign wire_2797 = lut_tile_1_1_chanxy_out[73];
    assign wire_2798 = lut_tile_1_1_chanxy_out[74];
    assign wire_2800 = lut_tile_1_1_chanxy_out[75];
    assign wire_2802 = lut_tile_1_1_chanxy_out[76];
    assign wire_2804 = lut_tile_1_1_chanxy_out[77];
    assign wire_2805 = lut_tile_1_1_chanxy_out[78];
    assign wire_2806 = lut_tile_1_1_chanxy_out[79];
    assign wire_2808 = lut_tile_1_1_chanxy_out[80];
    assign wire_2810 = lut_tile_1_1_chanxy_out[81];
    assign wire_2812 = lut_tile_1_1_chanxy_out[82];
    assign wire_2813 = lut_tile_1_1_chanxy_out[83];
    assign wire_2814 = lut_tile_1_1_chanxy_out[84];
    assign wire_2816 = lut_tile_1_1_chanxy_out[85];
    assign wire_2818 = lut_tile_1_1_chanxy_out[86];
    assign wire_2820 = lut_tile_1_1_chanxy_out[87];
    assign wire_2821 = lut_tile_1_1_chanxy_out[88];
    assign wire_2822 = lut_tile_1_1_chanxy_out[89];
    assign wire_2824 = lut_tile_1_1_chanxy_out[90];
    assign wire_2826 = lut_tile_1_1_chanxy_out[91];
    assign wire_2828 = lut_tile_1_1_chanxy_out[92];
    assign wire_2829 = lut_tile_1_1_chanxy_out[93];
    assign wire_2830 = lut_tile_1_1_chanxy_out[94];
    assign wire_2832 = lut_tile_1_1_chanxy_out[95];
    assign wire_2834 = lut_tile_1_1_chanxy_out[96];
    assign wire_2836 = lut_tile_1_1_chanxy_out[97];
    assign wire_2837 = lut_tile_1_1_chanxy_out[98];
    assign wire_2838 = lut_tile_1_1_chanxy_out[99];
    assign wire_4600 = lut_tile_1_1_chanxy_out[100];
    assign wire_4602 = lut_tile_1_1_chanxy_out[101];
    assign wire_4604 = lut_tile_1_1_chanxy_out[102];
    assign wire_4605 = lut_tile_1_1_chanxy_out[103];
    assign wire_4606 = lut_tile_1_1_chanxy_out[104];
    assign wire_4608 = lut_tile_1_1_chanxy_out[105];
    assign wire_4610 = lut_tile_1_1_chanxy_out[106];
    assign wire_4612 = lut_tile_1_1_chanxy_out[107];
    assign wire_4613 = lut_tile_1_1_chanxy_out[108];
    assign wire_4614 = lut_tile_1_1_chanxy_out[109];
    assign wire_4616 = lut_tile_1_1_chanxy_out[110];
    assign wire_4618 = lut_tile_1_1_chanxy_out[111];
    assign wire_4620 = lut_tile_1_1_chanxy_out[112];
    assign wire_4621 = lut_tile_1_1_chanxy_out[113];
    assign wire_4622 = lut_tile_1_1_chanxy_out[114];
    assign wire_4624 = lut_tile_1_1_chanxy_out[115];
    assign wire_4626 = lut_tile_1_1_chanxy_out[116];
    assign wire_4628 = lut_tile_1_1_chanxy_out[117];
    assign wire_4629 = lut_tile_1_1_chanxy_out[118];
    assign wire_4630 = lut_tile_1_1_chanxy_out[119];
    assign wire_4632 = lut_tile_1_1_chanxy_out[120];
    assign wire_4634 = lut_tile_1_1_chanxy_out[121];
    assign wire_4636 = lut_tile_1_1_chanxy_out[122];
    assign wire_4637 = lut_tile_1_1_chanxy_out[123];
    assign wire_4638 = lut_tile_1_1_chanxy_out[124];
    assign wire_4640 = lut_tile_1_1_chanxy_out[125];
    assign wire_4642 = lut_tile_1_1_chanxy_out[126];
    assign wire_4644 = lut_tile_1_1_chanxy_out[127];
    assign wire_4645 = lut_tile_1_1_chanxy_out[128];
    assign wire_4646 = lut_tile_1_1_chanxy_out[129];
    assign wire_4648 = lut_tile_1_1_chanxy_out[130];
    assign wire_4650 = lut_tile_1_1_chanxy_out[131];
    assign wire_4652 = lut_tile_1_1_chanxy_out[132];
    assign wire_4653 = lut_tile_1_1_chanxy_out[133];
    assign wire_4654 = lut_tile_1_1_chanxy_out[134];
    assign wire_4656 = lut_tile_1_1_chanxy_out[135];
    assign wire_4658 = lut_tile_1_1_chanxy_out[136];
    assign wire_4660 = lut_tile_1_1_chanxy_out[137];
    assign wire_4661 = lut_tile_1_1_chanxy_out[138];
    assign wire_4662 = lut_tile_1_1_chanxy_out[139];
    assign wire_4664 = lut_tile_1_1_chanxy_out[140];
    assign wire_4666 = lut_tile_1_1_chanxy_out[141];
    assign wire_4668 = lut_tile_1_1_chanxy_out[142];
    assign wire_4669 = lut_tile_1_1_chanxy_out[143];
    assign wire_4670 = lut_tile_1_1_chanxy_out[144];
    assign wire_4672 = lut_tile_1_1_chanxy_out[145];
    assign wire_4674 = lut_tile_1_1_chanxy_out[146];
    assign wire_4676 = lut_tile_1_1_chanxy_out[147];
    assign wire_4677 = lut_tile_1_1_chanxy_out[148];
    assign wire_4678 = lut_tile_1_1_chanxy_out[149];
    assign wire_4680 = lut_tile_1_1_chanxy_out[150];
    assign wire_4682 = lut_tile_1_1_chanxy_out[151];
    assign wire_4684 = lut_tile_1_1_chanxy_out[152];
    assign wire_4685 = lut_tile_1_1_chanxy_out[153];
    assign wire_4686 = lut_tile_1_1_chanxy_out[154];
    assign wire_4688 = lut_tile_1_1_chanxy_out[155];
    assign wire_4690 = lut_tile_1_1_chanxy_out[156];
    assign wire_4692 = lut_tile_1_1_chanxy_out[157];
    assign wire_4693 = lut_tile_1_1_chanxy_out[158];
    assign wire_4694 = lut_tile_1_1_chanxy_out[159];
    assign wire_4696 = lut_tile_1_1_chanxy_out[160];
    assign wire_4698 = lut_tile_1_1_chanxy_out[161];
    assign wire_4700 = lut_tile_1_1_chanxy_out[162];
    assign wire_4701 = lut_tile_1_1_chanxy_out[163];
    assign wire_4702 = lut_tile_1_1_chanxy_out[164];
    assign wire_4704 = lut_tile_1_1_chanxy_out[165];
    assign wire_4706 = lut_tile_1_1_chanxy_out[166];
    assign wire_4708 = lut_tile_1_1_chanxy_out[167];
    assign wire_4709 = lut_tile_1_1_chanxy_out[168];
    assign wire_4710 = lut_tile_1_1_chanxy_out[169];
    assign wire_4712 = lut_tile_1_1_chanxy_out[170];
    assign wire_4714 = lut_tile_1_1_chanxy_out[171];
    assign wire_4716 = lut_tile_1_1_chanxy_out[172];
    assign wire_4717 = lut_tile_1_1_chanxy_out[173];
    assign wire_4718 = lut_tile_1_1_chanxy_out[174];
    assign wire_4720 = lut_tile_1_1_chanxy_out[175];
    assign wire_4722 = lut_tile_1_1_chanxy_out[176];
    assign wire_4724 = lut_tile_1_1_chanxy_out[177];
    assign wire_4725 = lut_tile_1_1_chanxy_out[178];
    assign wire_4726 = lut_tile_1_1_chanxy_out[179];
    assign wire_4728 = lut_tile_1_1_chanxy_out[180];
    assign wire_4730 = lut_tile_1_1_chanxy_out[181];
    assign wire_4732 = lut_tile_1_1_chanxy_out[182];
    assign wire_4733 = lut_tile_1_1_chanxy_out[183];
    assign wire_4734 = lut_tile_1_1_chanxy_out[184];
    assign wire_4736 = lut_tile_1_1_chanxy_out[185];
    assign wire_4738 = lut_tile_1_1_chanxy_out[186];
    assign wire_4740 = lut_tile_1_1_chanxy_out[187];
    assign wire_4741 = lut_tile_1_1_chanxy_out[188];
    assign wire_4742 = lut_tile_1_1_chanxy_out[189];
    assign wire_4744 = lut_tile_1_1_chanxy_out[190];
    assign wire_4746 = lut_tile_1_1_chanxy_out[191];
    assign wire_4748 = lut_tile_1_1_chanxy_out[192];
    assign wire_4749 = lut_tile_1_1_chanxy_out[193];
    assign wire_4750 = lut_tile_1_1_chanxy_out[194];
    assign wire_4752 = lut_tile_1_1_chanxy_out[195];
    assign wire_4754 = lut_tile_1_1_chanxy_out[196];
    assign wire_4756 = lut_tile_1_1_chanxy_out[197];
    assign wire_4757 = lut_tile_1_1_chanxy_out[198];
    assign wire_4758 = lut_tile_1_1_chanxy_out[199];
   // CHANXY OUT
    assign lut_tile_1_2_chanxy_in = {wire_5119, wire_2919, wire_2879, wire_2878, wire_2785, wire_2784, wire_2731, wire_2730, wire_2686, wire_1091, wire_717, wire_2519, wire_2518, wire_2599, wire_2516, wire_2539, wire_2538, wire_2559, wire_2558, wire_5117, wire_2881, wire_2865, wire_2864, wire_2838, wire_2835, wire_2834, wire_2729, wire_2728, wire_1091, wire_717, wire_2513, wire_2512, wire_2433, wire_2432, wire_2511, wire_2510, wire_2597, wire_2508, wire_5115, wire_2883, wire_2851, wire_2850, wire_2833, wire_2832, wire_2830, wire_2779, wire_2778, wire_1091, wire_717, wire_2557, wire_2556, wire_2431, wire_2430, wire_2577, wire_2428, wire_2505, wire_2504, wire_5113, wire_2885, wire_2877, wire_2876, wire_2822, wire_2777, wire_2776, wire_2723, wire_2722, wire_1091, wire_717, wire_2537, wire_2536, wire_2425, wire_2424, wire_2503, wire_2502, wire_2423, wire_2422, wire_5111, wire_2887, wire_2863, wire_2862, wire_2827, wire_2826, wire_2814, wire_2721, wire_2720, wire_1091, wire_713, wire_2575, wire_2420, wire_2595, wire_2500, wire_2535, wire_2534, wire_2417, wire_2416, wire_5109, wire_2889, wire_2849, wire_2848, wire_2825, wire_2824, wire_2806, wire_2771, wire_2770, wire_1091, wire_713, wire_2415, wire_2414, wire_2555, wire_2554, wire_2497, wire_2496, wire_2573, wire_2412, wire_5107, wire_2891, wire_2875, wire_2874, wire_2798, wire_2769, wire_2768, wire_2715, wire_2714, wire_1091, wire_713, wire_2495, wire_2494, wire_2593, wire_2492, wire_2533, wire_2532, wire_2553, wire_2552, wire_5105, wire_2893, wire_2861, wire_2860, wire_2819, wire_2818, wire_2790, wire_2713, wire_2712, wire_1091, wire_713, wire_2489, wire_2488, wire_2409, wire_2408, wire_2487, wire_2486, wire_2591, wire_2484, wire_5103, wire_2895, wire_2847, wire_2846, wire_2817, wire_2816, wire_2782, wire_2763, wire_2762, wire_1087, wire_713, wire_2551, wire_2550, wire_2407, wire_2406, wire_2571, wire_2404, wire_2481, wire_2480, wire_5101, wire_2897, wire_2873, wire_2872, wire_2774, wire_2761, wire_2760, wire_2707, wire_2706, wire_1087, wire_713, wire_2531, wire_2530, wire_2401, wire_2400, wire_2479, wire_2478, wire_2399, wire_2398, wire_5099, wire_2899, wire_2859, wire_2858, wire_2811, wire_2810, wire_2766, wire_2705, wire_2704, wire_1087, wire_713, wire_2569, wire_2396, wire_1091, wire_2589, wire_2476, wire_1091, wire_2529, wire_2528, wire_1091, wire_2393, wire_2392, wire_1091, wire_5097, wire_2901, wire_2845, wire_2844, wire_2809, wire_2808, wire_2758, wire_2755, wire_2754, wire_1087, wire_713, wire_2391, wire_2390, wire_1091, wire_2549, wire_2548, wire_1091, wire_2473, wire_2472, wire_1091, wire_2567, wire_2388, wire_1091, wire_5095, wire_2903, wire_2871, wire_2870, wire_2753, wire_2752, wire_2750, wire_2699, wire_2698, wire_1087, wire_709, wire_2471, wire_2470, wire_1087, wire_2587, wire_2468, wire_1087, wire_2527, wire_2526, wire_1087, wire_2547, wire_2546, wire_1087, wire_5093, wire_2905, wire_2857, wire_2856, wire_2803, wire_2802, wire_2742, wire_2697, wire_2696, wire_1087, wire_709, wire_2465, wire_2464, wire_1087, wire_2385, wire_2384, wire_1087, wire_2463, wire_2462, wire_1087, wire_2585, wire_2460, wire_1087, wire_5091, wire_2907, wire_2843, wire_2842, wire_2801, wire_2800, wire_2747, wire_2746, wire_2734, wire_1087, wire_709, wire_2545, wire_2544, wire_717, wire_2383, wire_2382, wire_717, wire_2565, wire_2380, wire_717, wire_2457, wire_2456, wire_717, wire_5089, wire_2909, wire_2869, wire_2868, wire_2745, wire_2744, wire_2726, wire_2691, wire_2690, wire_1087, wire_709, wire_2525, wire_2524, wire_717, wire_2377, wire_2376, wire_717, wire_2455, wire_2454, wire_717, wire_2375, wire_2374, wire_717, wire_5087, wire_2911, wire_2855, wire_2854, wire_2795, wire_2794, wire_2718, wire_2689, wire_2688, wire_717, wire_709, wire_2563, wire_2372, wire_713, wire_2583, wire_2452, wire_713, wire_2523, wire_2522, wire_713, wire_2369, wire_2368, wire_713, wire_5085, wire_2913, wire_2841, wire_2840, wire_2793, wire_2792, wire_2739, wire_2738, wire_2710, wire_717, wire_709, wire_2367, wire_2366, wire_713, wire_2543, wire_2542, wire_713, wire_2449, wire_2448, wire_713, wire_2561, wire_2364, wire_713, wire_5083, wire_2915, wire_2867, wire_2866, wire_2737, wire_2736, wire_2702, wire_2683, wire_2682, wire_717, wire_709, wire_2447, wire_2446, wire_709, wire_2581, wire_2444, wire_709, wire_2521, wire_2520, wire_709, wire_2541, wire_2540, wire_709, wire_5081, wire_2917, wire_2853, wire_2852, wire_2787, wire_2786, wire_2694, wire_2681, wire_2680, wire_717, wire_709, wire_2441, wire_2440, wire_709, wire_2361, wire_2360, wire_709, wire_2439, wire_2438, wire_709, wire_2579, wire_2436, wire_709, wire_4797, wire_4759, wire_4758, wire_4756, wire_4705, wire_4704, wire_4651, wire_4650, wire_2836, wire_774, wire_766, wire_4795, wire_4755, wire_4754, wire_4703, wire_4702, wire_4649, wire_4648, wire_4604, wire_2828, wire_774, wire_766, wire_4793, wire_4753, wire_4752, wire_4699, wire_4698, wire_4647, wire_4646, wire_4612, wire_2820, wire_774, wire_766, wire_4791, wire_4751, wire_4750, wire_4697, wire_4696, wire_4643, wire_4642, wire_4620, wire_2812, wire_774, wire_766, wire_4789, wire_4747, wire_4746, wire_4695, wire_4694, wire_4641, wire_4640, wire_4628, wire_2804, wire_774, wire_716, wire_4787, wire_4745, wire_4744, wire_4691, wire_4690, wire_4639, wire_4638, wire_4636, wire_2796, wire_774, wire_716, wire_4785, wire_4743, wire_4742, wire_4689, wire_4688, wire_4644, wire_4635, wire_4634, wire_2788, wire_774, wire_716, wire_4783, wire_4739, wire_4738, wire_4687, wire_4686, wire_4652, wire_4633, wire_4632, wire_2780, wire_774, wire_716, wire_4781, wire_4737, wire_4736, wire_4683, wire_4682, wire_4660, wire_4631, wire_4630, wire_2772, wire_770, wire_716, wire_4779, wire_4735, wire_4734, wire_4681, wire_4680, wire_4668, wire_4627, wire_4626, wire_2764, wire_770, wire_716, wire_4777, wire_4731, wire_4730, wire_4679, wire_4678, wire_4676, wire_4625, wire_4624, wire_2756, wire_770, wire_716, wire_4775, wire_4729, wire_4728, wire_4684, wire_4675, wire_4674, wire_4623, wire_4622, wire_2748, wire_770, wire_716, wire_4773, wire_4727, wire_4726, wire_4692, wire_4673, wire_4672, wire_4619, wire_4618, wire_2740, wire_770, wire_712, wire_4771, wire_4723, wire_4722, wire_4700, wire_4671, wire_4670, wire_4617, wire_4616, wire_2732, wire_770, wire_712, wire_4769, wire_4721, wire_4720, wire_4708, wire_4667, wire_4666, wire_4615, wire_4614, wire_2724, wire_770, wire_712, wire_4767, wire_4719, wire_4718, wire_4716, wire_4665, wire_4664, wire_4611, wire_4610, wire_2716, wire_770, wire_712, wire_4765, wire_4724, wire_4715, wire_4714, wire_4663, wire_4662, wire_4609, wire_4608, wire_2708, wire_766, wire_712, wire_4763, wire_4732, wire_4713, wire_4712, wire_4659, wire_4658, wire_4607, wire_4606, wire_2700, wire_766, wire_712, wire_4761, wire_4740, wire_4711, wire_4710, wire_4657, wire_4656, wire_4603, wire_4602, wire_2692, wire_766, wire_712, wire_4799, wire_4748, wire_4707, wire_4706, wire_4655, wire_4654, wire_4601, wire_4600, wire_2684, wire_766, wire_712, wire_5083, wire_5077, wire_5076, wire_5070, wire_5025, wire_5024, wire_4971, wire_4970, wire_2919, wire_774, wire_766, wire_5085, wire_5075, wire_5074, wire_5062, wire_5021, wire_5020, wire_4969, wire_4968, wire_2917, wire_774, wire_766, wire_5087, wire_5073, wire_5072, wire_5054, wire_5019, wire_5018, wire_4965, wire_4964, wire_2915, wire_774, wire_766, wire_5089, wire_5069, wire_5068, wire_5046, wire_5017, wire_5016, wire_4963, wire_4962, wire_2913, wire_774, wire_766, wire_5091, wire_5067, wire_5066, wire_5038, wire_5013, wire_5012, wire_4961, wire_4960, wire_2911, wire_774, wire_716, wire_5093, wire_5065, wire_5064, wire_5030, wire_5011, wire_5010, wire_4957, wire_4956, wire_2909, wire_774, wire_716, wire_5095, wire_5061, wire_5060, wire_5022, wire_5009, wire_5008, wire_4955, wire_4954, wire_2907, wire_774, wire_716, wire_5097, wire_5059, wire_5058, wire_5014, wire_5005, wire_5004, wire_4953, wire_4952, wire_2905, wire_774, wire_716, wire_5099, wire_5057, wire_5056, wire_5006, wire_5003, wire_5002, wire_4949, wire_4948, wire_2903, wire_770, wire_716, wire_5101, wire_5053, wire_5052, wire_5001, wire_5000, wire_4998, wire_4947, wire_4946, wire_2901, wire_770, wire_716, wire_5103, wire_5051, wire_5050, wire_4997, wire_4996, wire_4990, wire_4945, wire_4944, wire_2899, wire_770, wire_716, wire_5105, wire_5049, wire_5048, wire_4995, wire_4994, wire_4982, wire_4941, wire_4940, wire_2897, wire_770, wire_716, wire_5107, wire_5045, wire_5044, wire_4993, wire_4992, wire_4974, wire_4939, wire_4938, wire_2895, wire_770, wire_712, wire_5109, wire_5043, wire_5042, wire_4989, wire_4988, wire_4966, wire_4937, wire_4936, wire_2893, wire_770, wire_712, wire_5111, wire_5041, wire_5040, wire_4987, wire_4986, wire_4958, wire_4933, wire_4932, wire_2891, wire_770, wire_712, wire_5113, wire_5037, wire_5036, wire_4985, wire_4984, wire_4950, wire_4931, wire_4930, wire_2889, wire_770, wire_712, wire_5115, wire_5035, wire_5034, wire_4981, wire_4980, wire_4942, wire_4929, wire_4928, wire_2887, wire_766, wire_712, wire_5117, wire_5033, wire_5032, wire_4979, wire_4978, wire_4934, wire_4925, wire_4924, wire_2885, wire_766, wire_712, wire_5119, wire_5029, wire_5028, wire_4977, wire_4976, wire_4926, wire_4923, wire_4922, wire_2883, wire_766, wire_712, wire_5081, wire_5078, wire_5027, wire_5026, wire_4973, wire_4972, wire_4921, wire_4920, wire_2881, wire_766, wire_712};
    // CHNAXY TOTAL: 860
    assign wire_2687 = lut_tile_1_2_chanxy_out[0];
    assign wire_2695 = lut_tile_1_2_chanxy_out[1];
    assign wire_2703 = lut_tile_1_2_chanxy_out[2];
    assign wire_2711 = lut_tile_1_2_chanxy_out[3];
    assign wire_2719 = lut_tile_1_2_chanxy_out[4];
    assign wire_2727 = lut_tile_1_2_chanxy_out[5];
    assign wire_2735 = lut_tile_1_2_chanxy_out[6];
    assign wire_2743 = lut_tile_1_2_chanxy_out[7];
    assign wire_2751 = lut_tile_1_2_chanxy_out[8];
    assign wire_2759 = lut_tile_1_2_chanxy_out[9];
    assign wire_2767 = lut_tile_1_2_chanxy_out[10];
    assign wire_2775 = lut_tile_1_2_chanxy_out[11];
    assign wire_2783 = lut_tile_1_2_chanxy_out[12];
    assign wire_2791 = lut_tile_1_2_chanxy_out[13];
    assign wire_2799 = lut_tile_1_2_chanxy_out[14];
    assign wire_2807 = lut_tile_1_2_chanxy_out[15];
    assign wire_2815 = lut_tile_1_2_chanxy_out[16];
    assign wire_2823 = lut_tile_1_2_chanxy_out[17];
    assign wire_2831 = lut_tile_1_2_chanxy_out[18];
    assign wire_2839 = lut_tile_1_2_chanxy_out[19];
    assign wire_2840 = lut_tile_1_2_chanxy_out[20];
    assign wire_2842 = lut_tile_1_2_chanxy_out[21];
    assign wire_2844 = lut_tile_1_2_chanxy_out[22];
    assign wire_2846 = lut_tile_1_2_chanxy_out[23];
    assign wire_2848 = lut_tile_1_2_chanxy_out[24];
    assign wire_2850 = lut_tile_1_2_chanxy_out[25];
    assign wire_2852 = lut_tile_1_2_chanxy_out[26];
    assign wire_2854 = lut_tile_1_2_chanxy_out[27];
    assign wire_2856 = lut_tile_1_2_chanxy_out[28];
    assign wire_2858 = lut_tile_1_2_chanxy_out[29];
    assign wire_2860 = lut_tile_1_2_chanxy_out[30];
    assign wire_2862 = lut_tile_1_2_chanxy_out[31];
    assign wire_2864 = lut_tile_1_2_chanxy_out[32];
    assign wire_2866 = lut_tile_1_2_chanxy_out[33];
    assign wire_2868 = lut_tile_1_2_chanxy_out[34];
    assign wire_2870 = lut_tile_1_2_chanxy_out[35];
    assign wire_2872 = lut_tile_1_2_chanxy_out[36];
    assign wire_2874 = lut_tile_1_2_chanxy_out[37];
    assign wire_2876 = lut_tile_1_2_chanxy_out[38];
    assign wire_2878 = lut_tile_1_2_chanxy_out[39];
    assign wire_4920 = lut_tile_1_2_chanxy_out[40];
    assign wire_4922 = lut_tile_1_2_chanxy_out[41];
    assign wire_4924 = lut_tile_1_2_chanxy_out[42];
    assign wire_4926 = lut_tile_1_2_chanxy_out[43];
    assign wire_4927 = lut_tile_1_2_chanxy_out[44];
    assign wire_4928 = lut_tile_1_2_chanxy_out[45];
    assign wire_4930 = lut_tile_1_2_chanxy_out[46];
    assign wire_4932 = lut_tile_1_2_chanxy_out[47];
    assign wire_4934 = lut_tile_1_2_chanxy_out[48];
    assign wire_4935 = lut_tile_1_2_chanxy_out[49];
    assign wire_4936 = lut_tile_1_2_chanxy_out[50];
    assign wire_4938 = lut_tile_1_2_chanxy_out[51];
    assign wire_4940 = lut_tile_1_2_chanxy_out[52];
    assign wire_4942 = lut_tile_1_2_chanxy_out[53];
    assign wire_4943 = lut_tile_1_2_chanxy_out[54];
    assign wire_4944 = lut_tile_1_2_chanxy_out[55];
    assign wire_4946 = lut_tile_1_2_chanxy_out[56];
    assign wire_4948 = lut_tile_1_2_chanxy_out[57];
    assign wire_4950 = lut_tile_1_2_chanxy_out[58];
    assign wire_4951 = lut_tile_1_2_chanxy_out[59];
    assign wire_4952 = lut_tile_1_2_chanxy_out[60];
    assign wire_4954 = lut_tile_1_2_chanxy_out[61];
    assign wire_4956 = lut_tile_1_2_chanxy_out[62];
    assign wire_4958 = lut_tile_1_2_chanxy_out[63];
    assign wire_4959 = lut_tile_1_2_chanxy_out[64];
    assign wire_4960 = lut_tile_1_2_chanxy_out[65];
    assign wire_4962 = lut_tile_1_2_chanxy_out[66];
    assign wire_4964 = lut_tile_1_2_chanxy_out[67];
    assign wire_4966 = lut_tile_1_2_chanxy_out[68];
    assign wire_4967 = lut_tile_1_2_chanxy_out[69];
    assign wire_4968 = lut_tile_1_2_chanxy_out[70];
    assign wire_4970 = lut_tile_1_2_chanxy_out[71];
    assign wire_4972 = lut_tile_1_2_chanxy_out[72];
    assign wire_4974 = lut_tile_1_2_chanxy_out[73];
    assign wire_4975 = lut_tile_1_2_chanxy_out[74];
    assign wire_4976 = lut_tile_1_2_chanxy_out[75];
    assign wire_4978 = lut_tile_1_2_chanxy_out[76];
    assign wire_4980 = lut_tile_1_2_chanxy_out[77];
    assign wire_4982 = lut_tile_1_2_chanxy_out[78];
    assign wire_4983 = lut_tile_1_2_chanxy_out[79];
    assign wire_4984 = lut_tile_1_2_chanxy_out[80];
    assign wire_4986 = lut_tile_1_2_chanxy_out[81];
    assign wire_4988 = lut_tile_1_2_chanxy_out[82];
    assign wire_4990 = lut_tile_1_2_chanxy_out[83];
    assign wire_4991 = lut_tile_1_2_chanxy_out[84];
    assign wire_4992 = lut_tile_1_2_chanxy_out[85];
    assign wire_4994 = lut_tile_1_2_chanxy_out[86];
    assign wire_4996 = lut_tile_1_2_chanxy_out[87];
    assign wire_4998 = lut_tile_1_2_chanxy_out[88];
    assign wire_4999 = lut_tile_1_2_chanxy_out[89];
    assign wire_5000 = lut_tile_1_2_chanxy_out[90];
    assign wire_5002 = lut_tile_1_2_chanxy_out[91];
    assign wire_5004 = lut_tile_1_2_chanxy_out[92];
    assign wire_5006 = lut_tile_1_2_chanxy_out[93];
    assign wire_5007 = lut_tile_1_2_chanxy_out[94];
    assign wire_5008 = lut_tile_1_2_chanxy_out[95];
    assign wire_5010 = lut_tile_1_2_chanxy_out[96];
    assign wire_5012 = lut_tile_1_2_chanxy_out[97];
    assign wire_5014 = lut_tile_1_2_chanxy_out[98];
    assign wire_5015 = lut_tile_1_2_chanxy_out[99];
    assign wire_5016 = lut_tile_1_2_chanxy_out[100];
    assign wire_5018 = lut_tile_1_2_chanxy_out[101];
    assign wire_5020 = lut_tile_1_2_chanxy_out[102];
    assign wire_5022 = lut_tile_1_2_chanxy_out[103];
    assign wire_5023 = lut_tile_1_2_chanxy_out[104];
    assign wire_5024 = lut_tile_1_2_chanxy_out[105];
    assign wire_5026 = lut_tile_1_2_chanxy_out[106];
    assign wire_5028 = lut_tile_1_2_chanxy_out[107];
    assign wire_5030 = lut_tile_1_2_chanxy_out[108];
    assign wire_5031 = lut_tile_1_2_chanxy_out[109];
    assign wire_5032 = lut_tile_1_2_chanxy_out[110];
    assign wire_5034 = lut_tile_1_2_chanxy_out[111];
    assign wire_5036 = lut_tile_1_2_chanxy_out[112];
    assign wire_5038 = lut_tile_1_2_chanxy_out[113];
    assign wire_5039 = lut_tile_1_2_chanxy_out[114];
    assign wire_5040 = lut_tile_1_2_chanxy_out[115];
    assign wire_5042 = lut_tile_1_2_chanxy_out[116];
    assign wire_5044 = lut_tile_1_2_chanxy_out[117];
    assign wire_5046 = lut_tile_1_2_chanxy_out[118];
    assign wire_5047 = lut_tile_1_2_chanxy_out[119];
    assign wire_5048 = lut_tile_1_2_chanxy_out[120];
    assign wire_5050 = lut_tile_1_2_chanxy_out[121];
    assign wire_5052 = lut_tile_1_2_chanxy_out[122];
    assign wire_5054 = lut_tile_1_2_chanxy_out[123];
    assign wire_5055 = lut_tile_1_2_chanxy_out[124];
    assign wire_5056 = lut_tile_1_2_chanxy_out[125];
    assign wire_5058 = lut_tile_1_2_chanxy_out[126];
    assign wire_5060 = lut_tile_1_2_chanxy_out[127];
    assign wire_5062 = lut_tile_1_2_chanxy_out[128];
    assign wire_5063 = lut_tile_1_2_chanxy_out[129];
    assign wire_5064 = lut_tile_1_2_chanxy_out[130];
    assign wire_5066 = lut_tile_1_2_chanxy_out[131];
    assign wire_5068 = lut_tile_1_2_chanxy_out[132];
    assign wire_5070 = lut_tile_1_2_chanxy_out[133];
    assign wire_5071 = lut_tile_1_2_chanxy_out[134];
    assign wire_5072 = lut_tile_1_2_chanxy_out[135];
    assign wire_5074 = lut_tile_1_2_chanxy_out[136];
    assign wire_5076 = lut_tile_1_2_chanxy_out[137];
    assign wire_5078 = lut_tile_1_2_chanxy_out[138];
    assign wire_5079 = lut_tile_1_2_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_1_3_chanxy_in = {wire_2639, wire_2518, wire_2599, wire_2598, wire_2539, wire_2538, wire_5439, wire_2959, wire_2919, wire_2918, wire_2853, wire_2852, wire_2787, wire_2786, wire_2680, wire_1467, wire_1093, wire_2559, wire_2558, wire_2513, wire_2512, wire_2433, wire_2432, wire_2637, wire_2510, wire_5437, wire_2921, wire_2905, wire_2904, wire_2879, wire_2878, wire_2832, wire_2731, wire_2730, wire_1467, wire_1093, wire_2597, wire_2596, wire_2557, wire_2556, wire_2617, wire_2430, wire_2577, wire_2576, wire_5435, wire_2923, wire_2891, wire_2890, wire_2865, wire_2864, wire_2835, wire_2834, wire_2824, wire_1467, wire_1093, wire_2505, wire_2504, wire_2537, wire_2536, wire_2425, wire_2424, wire_2635, wire_2502, wire_5433, wire_2925, wire_2917, wire_2916, wire_2851, wire_2850, wire_2816, wire_2779, wire_2778, wire_1467, wire_1093, wire_2615, wire_2422, wire_2575, wire_2574, wire_2595, wire_2594, wire_2535, wire_2534, wire_5431, wire_2927, wire_2903, wire_2902, wire_2877, wire_2876, wire_2808, wire_2723, wire_2722, wire_1467, wire_1089, wire_2417, wire_2416, wire_2613, wire_2414, wire_2555, wire_2554, wire_2497, wire_2496, wire_5429, wire_2929, wire_2889, wire_2888, wire_2863, wire_2862, wire_2827, wire_2826, wire_2800, wire_1467, wire_1089, wire_2573, wire_2572, wire_2633, wire_2494, wire_2593, wire_2592, wire_2533, wire_2532, wire_5427, wire_2931, wire_2915, wire_2914, wire_2849, wire_2848, wire_2792, wire_2771, wire_2770, wire_1467, wire_1089, wire_2553, wire_2552, wire_2489, wire_2488, wire_2409, wire_2408, wire_2631, wire_2486, wire_5425, wire_2933, wire_2901, wire_2900, wire_2875, wire_2874, wire_2784, wire_2715, wire_2714, wire_1467, wire_1089, wire_2591, wire_2590, wire_2551, wire_2550, wire_2611, wire_2406, wire_2571, wire_2570, wire_5423, wire_2935, wire_2887, wire_2886, wire_2861, wire_2860, wire_2819, wire_2818, wire_2776, wire_1463, wire_1089, wire_2481, wire_2480, wire_2531, wire_2530, wire_2401, wire_2400, wire_2629, wire_2478, wire_5421, wire_2937, wire_2913, wire_2912, wire_2847, wire_2846, wire_2768, wire_2763, wire_2762, wire_1463, wire_1089, wire_2609, wire_2398, wire_2569, wire_2568, wire_1467, wire_2589, wire_2588, wire_1467, wire_2529, wire_2528, wire_1467, wire_5419, wire_2939, wire_2899, wire_2898, wire_2873, wire_2872, wire_2760, wire_2707, wire_2706, wire_1463, wire_1089, wire_2393, wire_2392, wire_1467, wire_2607, wire_2390, wire_1467, wire_2549, wire_2548, wire_1467, wire_2473, wire_2472, wire_1467, wire_5417, wire_2941, wire_2885, wire_2884, wire_2859, wire_2858, wire_2811, wire_2810, wire_2752, wire_1463, wire_1089, wire_2567, wire_2566, wire_1467, wire_2627, wire_2470, wire_1463, wire_2587, wire_2586, wire_1463, wire_2527, wire_2526, wire_1463, wire_5415, wire_2943, wire_2911, wire_2910, wire_2845, wire_2844, wire_2755, wire_2754, wire_2744, wire_1463, wire_1085, wire_2547, wire_2546, wire_1463, wire_2465, wire_2464, wire_1463, wire_2385, wire_2384, wire_1463, wire_2625, wire_2462, wire_1463, wire_5413, wire_2945, wire_2897, wire_2896, wire_2871, wire_2870, wire_2736, wire_2699, wire_2698, wire_1463, wire_1085, wire_2585, wire_2584, wire_1463, wire_2545, wire_2544, wire_1093, wire_2605, wire_2382, wire_1093, wire_2565, wire_2564, wire_1093, wire_5411, wire_2947, wire_2883, wire_2882, wire_2857, wire_2856, wire_2803, wire_2802, wire_2728, wire_1463, wire_1085, wire_2457, wire_2456, wire_1093, wire_2525, wire_2524, wire_1093, wire_2377, wire_2376, wire_1093, wire_2623, wire_2454, wire_1093, wire_5409, wire_2949, wire_2909, wire_2908, wire_2843, wire_2842, wire_2747, wire_2746, wire_2720, wire_1463, wire_1085, wire_2603, wire_2374, wire_1093, wire_2563, wire_2562, wire_1089, wire_2583, wire_2582, wire_1089, wire_2523, wire_2522, wire_1089, wire_5407, wire_2951, wire_2895, wire_2894, wire_2869, wire_2868, wire_2712, wire_2691, wire_2690, wire_1093, wire_1085, wire_2369, wire_2368, wire_1089, wire_2601, wire_2366, wire_1089, wire_2543, wire_2542, wire_1089, wire_2449, wire_2448, wire_1089, wire_5405, wire_2953, wire_2881, wire_2880, wire_2855, wire_2854, wire_2795, wire_2794, wire_2704, wire_1093, wire_1085, wire_2561, wire_2560, wire_1089, wire_2621, wire_2446, wire_1085, wire_2581, wire_2580, wire_1085, wire_2521, wire_2520, wire_1085, wire_5403, wire_2955, wire_2907, wire_2906, wire_2841, wire_2840, wire_2739, wire_2738, wire_2696, wire_1093, wire_1085, wire_2541, wire_2540, wire_1085, wire_2441, wire_2440, wire_1085, wire_2361, wire_2360, wire_1085, wire_2619, wire_2438, wire_1085, wire_5401, wire_2957, wire_2893, wire_2892, wire_2867, wire_2866, wire_2688, wire_2683, wire_2682, wire_1093, wire_1085, wire_2579, wire_2578, wire_1085, wire_5117, wire_5078, wire_5077, wire_5076, wire_5025, wire_5024, wire_4971, wire_4970, wire_2838, wire_1150, wire_1142, wire_5115, wire_5075, wire_5074, wire_5021, wire_5020, wire_4969, wire_4968, wire_4926, wire_2830, wire_1150, wire_1142, wire_5113, wire_5073, wire_5072, wire_5019, wire_5018, wire_4965, wire_4964, wire_4934, wire_2822, wire_1150, wire_1142, wire_5111, wire_5069, wire_5068, wire_5017, wire_5016, wire_4963, wire_4962, wire_4942, wire_2814, wire_1150, wire_1142, wire_5109, wire_5067, wire_5066, wire_5013, wire_5012, wire_4961, wire_4960, wire_4950, wire_2806, wire_1150, wire_1092, wire_5107, wire_5065, wire_5064, wire_5011, wire_5010, wire_4958, wire_4957, wire_4956, wire_2798, wire_1150, wire_1092, wire_5105, wire_5061, wire_5060, wire_5009, wire_5008, wire_4966, wire_4955, wire_4954, wire_2790, wire_1150, wire_1092, wire_5103, wire_5059, wire_5058, wire_5005, wire_5004, wire_4974, wire_4953, wire_4952, wire_2782, wire_1150, wire_1092, wire_5101, wire_5057, wire_5056, wire_5003, wire_5002, wire_4982, wire_4949, wire_4948, wire_2774, wire_1146, wire_1092, wire_5099, wire_5053, wire_5052, wire_5001, wire_5000, wire_4990, wire_4947, wire_4946, wire_2766, wire_1146, wire_1092, wire_5097, wire_5051, wire_5050, wire_4998, wire_4997, wire_4996, wire_4945, wire_4944, wire_2758, wire_1146, wire_1092, wire_5095, wire_5049, wire_5048, wire_5006, wire_4995, wire_4994, wire_4941, wire_4940, wire_2750, wire_1146, wire_1092, wire_5093, wire_5045, wire_5044, wire_5014, wire_4993, wire_4992, wire_4939, wire_4938, wire_2742, wire_1146, wire_1088, wire_5091, wire_5043, wire_5042, wire_5022, wire_4989, wire_4988, wire_4937, wire_4936, wire_2734, wire_1146, wire_1088, wire_5089, wire_5041, wire_5040, wire_5030, wire_4987, wire_4986, wire_4933, wire_4932, wire_2726, wire_1146, wire_1088, wire_5087, wire_5038, wire_5037, wire_5036, wire_4985, wire_4984, wire_4931, wire_4930, wire_2718, wire_1146, wire_1088, wire_5085, wire_5046, wire_5035, wire_5034, wire_4981, wire_4980, wire_4929, wire_4928, wire_2710, wire_1142, wire_1088, wire_5083, wire_5054, wire_5033, wire_5032, wire_4979, wire_4978, wire_4925, wire_4924, wire_2702, wire_1142, wire_1088, wire_5081, wire_5062, wire_5029, wire_5028, wire_4977, wire_4976, wire_4923, wire_4922, wire_2694, wire_1142, wire_1088, wire_5119, wire_5070, wire_5027, wire_5026, wire_4973, wire_4972, wire_4921, wire_4920, wire_2686, wire_1142, wire_1088, wire_5403, wire_5399, wire_5398, wire_5384, wire_5347, wire_5346, wire_5293, wire_5292, wire_2959, wire_1150, wire_1142, wire_5405, wire_5397, wire_5396, wire_5376, wire_5343, wire_5342, wire_5291, wire_5290, wire_2957, wire_1150, wire_1142, wire_5407, wire_5395, wire_5394, wire_5368, wire_5341, wire_5340, wire_5287, wire_5286, wire_2955, wire_1150, wire_1142, wire_5409, wire_5391, wire_5390, wire_5360, wire_5339, wire_5338, wire_5285, wire_5284, wire_2953, wire_1150, wire_1142, wire_5411, wire_5389, wire_5388, wire_5352, wire_5335, wire_5334, wire_5283, wire_5282, wire_2951, wire_1150, wire_1092, wire_5413, wire_5387, wire_5386, wire_5344, wire_5333, wire_5332, wire_5279, wire_5278, wire_2949, wire_1150, wire_1092, wire_5415, wire_5383, wire_5382, wire_5336, wire_5331, wire_5330, wire_5277, wire_5276, wire_2947, wire_1150, wire_1092, wire_5417, wire_5381, wire_5380, wire_5328, wire_5327, wire_5326, wire_5275, wire_5274, wire_2945, wire_1150, wire_1092, wire_5419, wire_5379, wire_5378, wire_5325, wire_5324, wire_5320, wire_5271, wire_5270, wire_2943, wire_1146, wire_1092, wire_5421, wire_5375, wire_5374, wire_5323, wire_5322, wire_5312, wire_5269, wire_5268, wire_2941, wire_1146, wire_1092, wire_5423, wire_5373, wire_5372, wire_5319, wire_5318, wire_5304, wire_5267, wire_5266, wire_2939, wire_1146, wire_1092, wire_5425, wire_5371, wire_5370, wire_5317, wire_5316, wire_5296, wire_5263, wire_5262, wire_2937, wire_1146, wire_1092, wire_5427, wire_5367, wire_5366, wire_5315, wire_5314, wire_5288, wire_5261, wire_5260, wire_2935, wire_1146, wire_1088, wire_5429, wire_5365, wire_5364, wire_5311, wire_5310, wire_5280, wire_5259, wire_5258, wire_2933, wire_1146, wire_1088, wire_5431, wire_5363, wire_5362, wire_5309, wire_5308, wire_5272, wire_5255, wire_5254, wire_2931, wire_1146, wire_1088, wire_5433, wire_5359, wire_5358, wire_5307, wire_5306, wire_5264, wire_5253, wire_5252, wire_2929, wire_1146, wire_1088, wire_5435, wire_5357, wire_5356, wire_5303, wire_5302, wire_5256, wire_5251, wire_5250, wire_2927, wire_1142, wire_1088, wire_5437, wire_5355, wire_5354, wire_5301, wire_5300, wire_5248, wire_5247, wire_5246, wire_2925, wire_1142, wire_1088, wire_5439, wire_5351, wire_5350, wire_5299, wire_5298, wire_5245, wire_5244, wire_5240, wire_2923, wire_1142, wire_1088, wire_5401, wire_5392, wire_5349, wire_5348, wire_5295, wire_5294, wire_5243, wire_5242, wire_2921, wire_1142, wire_1088};
    // CHNAXY TOTAL: 860
    assign wire_2681 = lut_tile_1_3_chanxy_out[0];
    assign wire_2689 = lut_tile_1_3_chanxy_out[1];
    assign wire_2697 = lut_tile_1_3_chanxy_out[2];
    assign wire_2705 = lut_tile_1_3_chanxy_out[3];
    assign wire_2713 = lut_tile_1_3_chanxy_out[4];
    assign wire_2721 = lut_tile_1_3_chanxy_out[5];
    assign wire_2729 = lut_tile_1_3_chanxy_out[6];
    assign wire_2737 = lut_tile_1_3_chanxy_out[7];
    assign wire_2745 = lut_tile_1_3_chanxy_out[8];
    assign wire_2753 = lut_tile_1_3_chanxy_out[9];
    assign wire_2761 = lut_tile_1_3_chanxy_out[10];
    assign wire_2769 = lut_tile_1_3_chanxy_out[11];
    assign wire_2777 = lut_tile_1_3_chanxy_out[12];
    assign wire_2785 = lut_tile_1_3_chanxy_out[13];
    assign wire_2793 = lut_tile_1_3_chanxy_out[14];
    assign wire_2801 = lut_tile_1_3_chanxy_out[15];
    assign wire_2809 = lut_tile_1_3_chanxy_out[16];
    assign wire_2817 = lut_tile_1_3_chanxy_out[17];
    assign wire_2825 = lut_tile_1_3_chanxy_out[18];
    assign wire_2833 = lut_tile_1_3_chanxy_out[19];
    assign wire_2880 = lut_tile_1_3_chanxy_out[20];
    assign wire_2882 = lut_tile_1_3_chanxy_out[21];
    assign wire_2884 = lut_tile_1_3_chanxy_out[22];
    assign wire_2886 = lut_tile_1_3_chanxy_out[23];
    assign wire_2888 = lut_tile_1_3_chanxy_out[24];
    assign wire_2890 = lut_tile_1_3_chanxy_out[25];
    assign wire_2892 = lut_tile_1_3_chanxy_out[26];
    assign wire_2894 = lut_tile_1_3_chanxy_out[27];
    assign wire_2896 = lut_tile_1_3_chanxy_out[28];
    assign wire_2898 = lut_tile_1_3_chanxy_out[29];
    assign wire_2900 = lut_tile_1_3_chanxy_out[30];
    assign wire_2902 = lut_tile_1_3_chanxy_out[31];
    assign wire_2904 = lut_tile_1_3_chanxy_out[32];
    assign wire_2906 = lut_tile_1_3_chanxy_out[33];
    assign wire_2908 = lut_tile_1_3_chanxy_out[34];
    assign wire_2910 = lut_tile_1_3_chanxy_out[35];
    assign wire_2912 = lut_tile_1_3_chanxy_out[36];
    assign wire_2914 = lut_tile_1_3_chanxy_out[37];
    assign wire_2916 = lut_tile_1_3_chanxy_out[38];
    assign wire_2918 = lut_tile_1_3_chanxy_out[39];
    assign wire_5240 = lut_tile_1_3_chanxy_out[40];
    assign wire_5241 = lut_tile_1_3_chanxy_out[41];
    assign wire_5242 = lut_tile_1_3_chanxy_out[42];
    assign wire_5244 = lut_tile_1_3_chanxy_out[43];
    assign wire_5246 = lut_tile_1_3_chanxy_out[44];
    assign wire_5248 = lut_tile_1_3_chanxy_out[45];
    assign wire_5249 = lut_tile_1_3_chanxy_out[46];
    assign wire_5250 = lut_tile_1_3_chanxy_out[47];
    assign wire_5252 = lut_tile_1_3_chanxy_out[48];
    assign wire_5254 = lut_tile_1_3_chanxy_out[49];
    assign wire_5256 = lut_tile_1_3_chanxy_out[50];
    assign wire_5257 = lut_tile_1_3_chanxy_out[51];
    assign wire_5258 = lut_tile_1_3_chanxy_out[52];
    assign wire_5260 = lut_tile_1_3_chanxy_out[53];
    assign wire_5262 = lut_tile_1_3_chanxy_out[54];
    assign wire_5264 = lut_tile_1_3_chanxy_out[55];
    assign wire_5265 = lut_tile_1_3_chanxy_out[56];
    assign wire_5266 = lut_tile_1_3_chanxy_out[57];
    assign wire_5268 = lut_tile_1_3_chanxy_out[58];
    assign wire_5270 = lut_tile_1_3_chanxy_out[59];
    assign wire_5272 = lut_tile_1_3_chanxy_out[60];
    assign wire_5273 = lut_tile_1_3_chanxy_out[61];
    assign wire_5274 = lut_tile_1_3_chanxy_out[62];
    assign wire_5276 = lut_tile_1_3_chanxy_out[63];
    assign wire_5278 = lut_tile_1_3_chanxy_out[64];
    assign wire_5280 = lut_tile_1_3_chanxy_out[65];
    assign wire_5281 = lut_tile_1_3_chanxy_out[66];
    assign wire_5282 = lut_tile_1_3_chanxy_out[67];
    assign wire_5284 = lut_tile_1_3_chanxy_out[68];
    assign wire_5286 = lut_tile_1_3_chanxy_out[69];
    assign wire_5288 = lut_tile_1_3_chanxy_out[70];
    assign wire_5289 = lut_tile_1_3_chanxy_out[71];
    assign wire_5290 = lut_tile_1_3_chanxy_out[72];
    assign wire_5292 = lut_tile_1_3_chanxy_out[73];
    assign wire_5294 = lut_tile_1_3_chanxy_out[74];
    assign wire_5296 = lut_tile_1_3_chanxy_out[75];
    assign wire_5297 = lut_tile_1_3_chanxy_out[76];
    assign wire_5298 = lut_tile_1_3_chanxy_out[77];
    assign wire_5300 = lut_tile_1_3_chanxy_out[78];
    assign wire_5302 = lut_tile_1_3_chanxy_out[79];
    assign wire_5304 = lut_tile_1_3_chanxy_out[80];
    assign wire_5305 = lut_tile_1_3_chanxy_out[81];
    assign wire_5306 = lut_tile_1_3_chanxy_out[82];
    assign wire_5308 = lut_tile_1_3_chanxy_out[83];
    assign wire_5310 = lut_tile_1_3_chanxy_out[84];
    assign wire_5312 = lut_tile_1_3_chanxy_out[85];
    assign wire_5313 = lut_tile_1_3_chanxy_out[86];
    assign wire_5314 = lut_tile_1_3_chanxy_out[87];
    assign wire_5316 = lut_tile_1_3_chanxy_out[88];
    assign wire_5318 = lut_tile_1_3_chanxy_out[89];
    assign wire_5320 = lut_tile_1_3_chanxy_out[90];
    assign wire_5321 = lut_tile_1_3_chanxy_out[91];
    assign wire_5322 = lut_tile_1_3_chanxy_out[92];
    assign wire_5324 = lut_tile_1_3_chanxy_out[93];
    assign wire_5326 = lut_tile_1_3_chanxy_out[94];
    assign wire_5328 = lut_tile_1_3_chanxy_out[95];
    assign wire_5329 = lut_tile_1_3_chanxy_out[96];
    assign wire_5330 = lut_tile_1_3_chanxy_out[97];
    assign wire_5332 = lut_tile_1_3_chanxy_out[98];
    assign wire_5334 = lut_tile_1_3_chanxy_out[99];
    assign wire_5336 = lut_tile_1_3_chanxy_out[100];
    assign wire_5337 = lut_tile_1_3_chanxy_out[101];
    assign wire_5338 = lut_tile_1_3_chanxy_out[102];
    assign wire_5340 = lut_tile_1_3_chanxy_out[103];
    assign wire_5342 = lut_tile_1_3_chanxy_out[104];
    assign wire_5344 = lut_tile_1_3_chanxy_out[105];
    assign wire_5345 = lut_tile_1_3_chanxy_out[106];
    assign wire_5346 = lut_tile_1_3_chanxy_out[107];
    assign wire_5348 = lut_tile_1_3_chanxy_out[108];
    assign wire_5350 = lut_tile_1_3_chanxy_out[109];
    assign wire_5352 = lut_tile_1_3_chanxy_out[110];
    assign wire_5353 = lut_tile_1_3_chanxy_out[111];
    assign wire_5354 = lut_tile_1_3_chanxy_out[112];
    assign wire_5356 = lut_tile_1_3_chanxy_out[113];
    assign wire_5358 = lut_tile_1_3_chanxy_out[114];
    assign wire_5360 = lut_tile_1_3_chanxy_out[115];
    assign wire_5361 = lut_tile_1_3_chanxy_out[116];
    assign wire_5362 = lut_tile_1_3_chanxy_out[117];
    assign wire_5364 = lut_tile_1_3_chanxy_out[118];
    assign wire_5366 = lut_tile_1_3_chanxy_out[119];
    assign wire_5368 = lut_tile_1_3_chanxy_out[120];
    assign wire_5369 = lut_tile_1_3_chanxy_out[121];
    assign wire_5370 = lut_tile_1_3_chanxy_out[122];
    assign wire_5372 = lut_tile_1_3_chanxy_out[123];
    assign wire_5374 = lut_tile_1_3_chanxy_out[124];
    assign wire_5376 = lut_tile_1_3_chanxy_out[125];
    assign wire_5377 = lut_tile_1_3_chanxy_out[126];
    assign wire_5378 = lut_tile_1_3_chanxy_out[127];
    assign wire_5380 = lut_tile_1_3_chanxy_out[128];
    assign wire_5382 = lut_tile_1_3_chanxy_out[129];
    assign wire_5384 = lut_tile_1_3_chanxy_out[130];
    assign wire_5385 = lut_tile_1_3_chanxy_out[131];
    assign wire_5386 = lut_tile_1_3_chanxy_out[132];
    assign wire_5388 = lut_tile_1_3_chanxy_out[133];
    assign wire_5390 = lut_tile_1_3_chanxy_out[134];
    assign wire_5392 = lut_tile_1_3_chanxy_out[135];
    assign wire_5393 = lut_tile_1_3_chanxy_out[136];
    assign wire_5394 = lut_tile_1_3_chanxy_out[137];
    assign wire_5396 = lut_tile_1_3_chanxy_out[138];
    assign wire_5398 = lut_tile_1_3_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_1_4_chanxy_in = {wire_2639, wire_2638, wire_2599, wire_2598, wire_5759, wire_2999, wire_2947, wire_2946, wire_2919, wire_2918, wire_2853, wire_2852, wire_2682, wire_1843, wire_1469, wire_2539, wire_2538, wire_2559, wire_2558, wire_2679, wire_2512, wire_2659, wire_2432, wire_5757, wire_2961, wire_2933, wire_2932, wire_2905, wire_2904, wire_2879, wire_2878, wire_2834, wire_1843, wire_1469, wire_2637, wire_2636, wire_2597, wire_2596, wire_2557, wire_2556, wire_2617, wire_2616, wire_5755, wire_2963, wire_2959, wire_2958, wire_2891, wire_2890, wire_2865, wire_2864, wire_2826, wire_1843, wire_1469, wire_2577, wire_2576, wire_2677, wire_2504, wire_2537, wire_2536, wire_2657, wire_2424, wire_5753, wire_2965, wire_2945, wire_2944, wire_2917, wire_2916, wire_2851, wire_2850, wire_2818, wire_1843, wire_1469, wire_2635, wire_2634, wire_2615, wire_2614, wire_2575, wire_2574, wire_2595, wire_2594, wire_5751, wire_2967, wire_2931, wire_2930, wire_2903, wire_2902, wire_2877, wire_2876, wire_2810, wire_1843, wire_1465, wire_2535, wire_2534, wire_2655, wire_2416, wire_2613, wire_2612, wire_2555, wire_2554, wire_5749, wire_2969, wire_2957, wire_2956, wire_2889, wire_2888, wire_2863, wire_2862, wire_2802, wire_1843, wire_1465, wire_2675, wire_2496, wire_2573, wire_2572, wire_2633, wire_2632, wire_2593, wire_2592, wire_5747, wire_2971, wire_2943, wire_2942, wire_2915, wire_2914, wire_2849, wire_2848, wire_2794, wire_1843, wire_1465, wire_2533, wire_2532, wire_2553, wire_2552, wire_2673, wire_2488, wire_2653, wire_2408, wire_5745, wire_2973, wire_2929, wire_2928, wire_2901, wire_2900, wire_2875, wire_2874, wire_2786, wire_1843, wire_1465, wire_2631, wire_2630, wire_2591, wire_2590, wire_2551, wire_2550, wire_2611, wire_2610, wire_5743, wire_2975, wire_2955, wire_2954, wire_2887, wire_2886, wire_2861, wire_2860, wire_2778, wire_1839, wire_1465, wire_2571, wire_2570, wire_2671, wire_2480, wire_2531, wire_2530, wire_2651, wire_2400, wire_5741, wire_2977, wire_2941, wire_2940, wire_2913, wire_2912, wire_2847, wire_2846, wire_2770, wire_1839, wire_1465, wire_2629, wire_2628, wire_2609, wire_2608, wire_2569, wire_2568, wire_1843, wire_2589, wire_2588, wire_1843, wire_5739, wire_2979, wire_2927, wire_2926, wire_2899, wire_2898, wire_2873, wire_2872, wire_2762, wire_1839, wire_1465, wire_2529, wire_2528, wire_1843, wire_2649, wire_2392, wire_1843, wire_2607, wire_2606, wire_1843, wire_2549, wire_2548, wire_1843, wire_5737, wire_2981, wire_2953, wire_2952, wire_2885, wire_2884, wire_2859, wire_2858, wire_2754, wire_1839, wire_1465, wire_2669, wire_2472, wire_1843, wire_2567, wire_2566, wire_1843, wire_2627, wire_2626, wire_1839, wire_2587, wire_2586, wire_1839, wire_5735, wire_2983, wire_2939, wire_2938, wire_2911, wire_2910, wire_2845, wire_2844, wire_2746, wire_1839, wire_1461, wire_2527, wire_2526, wire_1839, wire_2547, wire_2546, wire_1839, wire_2667, wire_2464, wire_1839, wire_2647, wire_2384, wire_1839, wire_5733, wire_2985, wire_2925, wire_2924, wire_2897, wire_2896, wire_2871, wire_2870, wire_2738, wire_1839, wire_1461, wire_2625, wire_2624, wire_1839, wire_2585, wire_2584, wire_1839, wire_2545, wire_2544, wire_1469, wire_2605, wire_2604, wire_1469, wire_5731, wire_2987, wire_2951, wire_2950, wire_2883, wire_2882, wire_2857, wire_2856, wire_2730, wire_1839, wire_1461, wire_2565, wire_2564, wire_1469, wire_2665, wire_2456, wire_1469, wire_2525, wire_2524, wire_1469, wire_2645, wire_2376, wire_1469, wire_5729, wire_2989, wire_2937, wire_2936, wire_2909, wire_2908, wire_2843, wire_2842, wire_2722, wire_1839, wire_1461, wire_2623, wire_2622, wire_1469, wire_2603, wire_2602, wire_1469, wire_2563, wire_2562, wire_1465, wire_2583, wire_2582, wire_1465, wire_5727, wire_2991, wire_2923, wire_2922, wire_2895, wire_2894, wire_2869, wire_2868, wire_2714, wire_1469, wire_1461, wire_2523, wire_2522, wire_1465, wire_2643, wire_2368, wire_1465, wire_2601, wire_2600, wire_1465, wire_2543, wire_2542, wire_1465, wire_5725, wire_2993, wire_2949, wire_2948, wire_2881, wire_2880, wire_2855, wire_2854, wire_2706, wire_1469, wire_1461, wire_2663, wire_2448, wire_1465, wire_2561, wire_2560, wire_1465, wire_2621, wire_2620, wire_1461, wire_2581, wire_2580, wire_1461, wire_5723, wire_2995, wire_2935, wire_2934, wire_2907, wire_2906, wire_2841, wire_2840, wire_2698, wire_1469, wire_1461, wire_2521, wire_2520, wire_1461, wire_2541, wire_2540, wire_1461, wire_2661, wire_2440, wire_1461, wire_2641, wire_2360, wire_1461, wire_5721, wire_2997, wire_2921, wire_2920, wire_2893, wire_2892, wire_2867, wire_2866, wire_2690, wire_1469, wire_1461, wire_2619, wire_2618, wire_1461, wire_2579, wire_2578, wire_1461, wire_5437, wire_5399, wire_5398, wire_5392, wire_5347, wire_5346, wire_5293, wire_5292, wire_2832, wire_1526, wire_1518, wire_5435, wire_5397, wire_5396, wire_5343, wire_5342, wire_5291, wire_5290, wire_5240, wire_2824, wire_1526, wire_1518, wire_5433, wire_5395, wire_5394, wire_5341, wire_5340, wire_5287, wire_5286, wire_5248, wire_2816, wire_1526, wire_1518, wire_5431, wire_5391, wire_5390, wire_5339, wire_5338, wire_5285, wire_5284, wire_5256, wire_2808, wire_1526, wire_1518, wire_5429, wire_5389, wire_5388, wire_5335, wire_5334, wire_5283, wire_5282, wire_5264, wire_2800, wire_1526, wire_1468, wire_5427, wire_5387, wire_5386, wire_5333, wire_5332, wire_5279, wire_5278, wire_5272, wire_2792, wire_1526, wire_1468, wire_5425, wire_5383, wire_5382, wire_5331, wire_5330, wire_5280, wire_5277, wire_5276, wire_2784, wire_1526, wire_1468, wire_5423, wire_5381, wire_5380, wire_5327, wire_5326, wire_5288, wire_5275, wire_5274, wire_2776, wire_1526, wire_1468, wire_5421, wire_5379, wire_5378, wire_5325, wire_5324, wire_5296, wire_5271, wire_5270, wire_2768, wire_1522, wire_1468, wire_5419, wire_5375, wire_5374, wire_5323, wire_5322, wire_5304, wire_5269, wire_5268, wire_2760, wire_1522, wire_1468, wire_5417, wire_5373, wire_5372, wire_5319, wire_5318, wire_5312, wire_5267, wire_5266, wire_2752, wire_1522, wire_1468, wire_5415, wire_5371, wire_5370, wire_5320, wire_5317, wire_5316, wire_5263, wire_5262, wire_2744, wire_1522, wire_1468, wire_5413, wire_5367, wire_5366, wire_5328, wire_5315, wire_5314, wire_5261, wire_5260, wire_2736, wire_1522, wire_1464, wire_5411, wire_5365, wire_5364, wire_5336, wire_5311, wire_5310, wire_5259, wire_5258, wire_2728, wire_1522, wire_1464, wire_5409, wire_5363, wire_5362, wire_5344, wire_5309, wire_5308, wire_5255, wire_5254, wire_2720, wire_1522, wire_1464, wire_5407, wire_5359, wire_5358, wire_5352, wire_5307, wire_5306, wire_5253, wire_5252, wire_2712, wire_1522, wire_1464, wire_5405, wire_5360, wire_5357, wire_5356, wire_5303, wire_5302, wire_5251, wire_5250, wire_2704, wire_1518, wire_1464, wire_5403, wire_5368, wire_5355, wire_5354, wire_5301, wire_5300, wire_5247, wire_5246, wire_2696, wire_1518, wire_1464, wire_5401, wire_5376, wire_5351, wire_5350, wire_5299, wire_5298, wire_5245, wire_5244, wire_2688, wire_1518, wire_1464, wire_5439, wire_5384, wire_5349, wire_5348, wire_5295, wire_5294, wire_5243, wire_5242, wire_2680, wire_1518, wire_1464, wire_5723, wire_5719, wire_5718, wire_5706, wire_5665, wire_5664, wire_5613, wire_5612, wire_2999, wire_1526, wire_1518, wire_5725, wire_5717, wire_5716, wire_5698, wire_5663, wire_5662, wire_5609, wire_5608, wire_2997, wire_1526, wire_1518, wire_5727, wire_5713, wire_5712, wire_5690, wire_5661, wire_5660, wire_5607, wire_5606, wire_2995, wire_1526, wire_1518, wire_5729, wire_5711, wire_5710, wire_5682, wire_5657, wire_5656, wire_5605, wire_5604, wire_2993, wire_1526, wire_1518, wire_5731, wire_5709, wire_5708, wire_5674, wire_5655, wire_5654, wire_5601, wire_5600, wire_2991, wire_1526, wire_1468, wire_5733, wire_5705, wire_5704, wire_5666, wire_5653, wire_5652, wire_5599, wire_5598, wire_2989, wire_1526, wire_1468, wire_5735, wire_5703, wire_5702, wire_5658, wire_5649, wire_5648, wire_5597, wire_5596, wire_2987, wire_1526, wire_1468, wire_5737, wire_5701, wire_5700, wire_5650, wire_5647, wire_5646, wire_5593, wire_5592, wire_2985, wire_1526, wire_1468, wire_5739, wire_5697, wire_5696, wire_5645, wire_5644, wire_5642, wire_5591, wire_5590, wire_2983, wire_1522, wire_1468, wire_5741, wire_5695, wire_5694, wire_5641, wire_5640, wire_5634, wire_5589, wire_5588, wire_2981, wire_1522, wire_1468, wire_5743, wire_5693, wire_5692, wire_5639, wire_5638, wire_5626, wire_5585, wire_5584, wire_2979, wire_1522, wire_1468, wire_5745, wire_5689, wire_5688, wire_5637, wire_5636, wire_5618, wire_5583, wire_5582, wire_2977, wire_1522, wire_1468, wire_5747, wire_5687, wire_5686, wire_5633, wire_5632, wire_5610, wire_5581, wire_5580, wire_2975, wire_1522, wire_1464, wire_5749, wire_5685, wire_5684, wire_5631, wire_5630, wire_5602, wire_5577, wire_5576, wire_2973, wire_1522, wire_1464, wire_5751, wire_5681, wire_5680, wire_5629, wire_5628, wire_5594, wire_5575, wire_5574, wire_2971, wire_1522, wire_1464, wire_5753, wire_5679, wire_5678, wire_5625, wire_5624, wire_5586, wire_5573, wire_5572, wire_2969, wire_1522, wire_1464, wire_5755, wire_5677, wire_5676, wire_5623, wire_5622, wire_5578, wire_5569, wire_5568, wire_2967, wire_1518, wire_1464, wire_5757, wire_5673, wire_5672, wire_5621, wire_5620, wire_5570, wire_5567, wire_5566, wire_2965, wire_1518, wire_1464, wire_5759, wire_5671, wire_5670, wire_5617, wire_5616, wire_5565, wire_5564, wire_5562, wire_2963, wire_1518, wire_1464, wire_5721, wire_5714, wire_5669, wire_5668, wire_5615, wire_5614, wire_5561, wire_5560, wire_2961, wire_1518, wire_1464};
    // CHNAXY TOTAL: 860
    assign wire_2683 = lut_tile_1_4_chanxy_out[0];
    assign wire_2691 = lut_tile_1_4_chanxy_out[1];
    assign wire_2699 = lut_tile_1_4_chanxy_out[2];
    assign wire_2707 = lut_tile_1_4_chanxy_out[3];
    assign wire_2715 = lut_tile_1_4_chanxy_out[4];
    assign wire_2723 = lut_tile_1_4_chanxy_out[5];
    assign wire_2731 = lut_tile_1_4_chanxy_out[6];
    assign wire_2739 = lut_tile_1_4_chanxy_out[7];
    assign wire_2747 = lut_tile_1_4_chanxy_out[8];
    assign wire_2755 = lut_tile_1_4_chanxy_out[9];
    assign wire_2763 = lut_tile_1_4_chanxy_out[10];
    assign wire_2771 = lut_tile_1_4_chanxy_out[11];
    assign wire_2779 = lut_tile_1_4_chanxy_out[12];
    assign wire_2787 = lut_tile_1_4_chanxy_out[13];
    assign wire_2795 = lut_tile_1_4_chanxy_out[14];
    assign wire_2803 = lut_tile_1_4_chanxy_out[15];
    assign wire_2811 = lut_tile_1_4_chanxy_out[16];
    assign wire_2819 = lut_tile_1_4_chanxy_out[17];
    assign wire_2827 = lut_tile_1_4_chanxy_out[18];
    assign wire_2835 = lut_tile_1_4_chanxy_out[19];
    assign wire_2920 = lut_tile_1_4_chanxy_out[20];
    assign wire_2922 = lut_tile_1_4_chanxy_out[21];
    assign wire_2924 = lut_tile_1_4_chanxy_out[22];
    assign wire_2926 = lut_tile_1_4_chanxy_out[23];
    assign wire_2928 = lut_tile_1_4_chanxy_out[24];
    assign wire_2930 = lut_tile_1_4_chanxy_out[25];
    assign wire_2932 = lut_tile_1_4_chanxy_out[26];
    assign wire_2934 = lut_tile_1_4_chanxy_out[27];
    assign wire_2936 = lut_tile_1_4_chanxy_out[28];
    assign wire_2938 = lut_tile_1_4_chanxy_out[29];
    assign wire_2940 = lut_tile_1_4_chanxy_out[30];
    assign wire_2942 = lut_tile_1_4_chanxy_out[31];
    assign wire_2944 = lut_tile_1_4_chanxy_out[32];
    assign wire_2946 = lut_tile_1_4_chanxy_out[33];
    assign wire_2948 = lut_tile_1_4_chanxy_out[34];
    assign wire_2950 = lut_tile_1_4_chanxy_out[35];
    assign wire_2952 = lut_tile_1_4_chanxy_out[36];
    assign wire_2954 = lut_tile_1_4_chanxy_out[37];
    assign wire_2956 = lut_tile_1_4_chanxy_out[38];
    assign wire_2958 = lut_tile_1_4_chanxy_out[39];
    assign wire_5560 = lut_tile_1_4_chanxy_out[40];
    assign wire_5562 = lut_tile_1_4_chanxy_out[41];
    assign wire_5563 = lut_tile_1_4_chanxy_out[42];
    assign wire_5564 = lut_tile_1_4_chanxy_out[43];
    assign wire_5566 = lut_tile_1_4_chanxy_out[44];
    assign wire_5568 = lut_tile_1_4_chanxy_out[45];
    assign wire_5570 = lut_tile_1_4_chanxy_out[46];
    assign wire_5571 = lut_tile_1_4_chanxy_out[47];
    assign wire_5572 = lut_tile_1_4_chanxy_out[48];
    assign wire_5574 = lut_tile_1_4_chanxy_out[49];
    assign wire_5576 = lut_tile_1_4_chanxy_out[50];
    assign wire_5578 = lut_tile_1_4_chanxy_out[51];
    assign wire_5579 = lut_tile_1_4_chanxy_out[52];
    assign wire_5580 = lut_tile_1_4_chanxy_out[53];
    assign wire_5582 = lut_tile_1_4_chanxy_out[54];
    assign wire_5584 = lut_tile_1_4_chanxy_out[55];
    assign wire_5586 = lut_tile_1_4_chanxy_out[56];
    assign wire_5587 = lut_tile_1_4_chanxy_out[57];
    assign wire_5588 = lut_tile_1_4_chanxy_out[58];
    assign wire_5590 = lut_tile_1_4_chanxy_out[59];
    assign wire_5592 = lut_tile_1_4_chanxy_out[60];
    assign wire_5594 = lut_tile_1_4_chanxy_out[61];
    assign wire_5595 = lut_tile_1_4_chanxy_out[62];
    assign wire_5596 = lut_tile_1_4_chanxy_out[63];
    assign wire_5598 = lut_tile_1_4_chanxy_out[64];
    assign wire_5600 = lut_tile_1_4_chanxy_out[65];
    assign wire_5602 = lut_tile_1_4_chanxy_out[66];
    assign wire_5603 = lut_tile_1_4_chanxy_out[67];
    assign wire_5604 = lut_tile_1_4_chanxy_out[68];
    assign wire_5606 = lut_tile_1_4_chanxy_out[69];
    assign wire_5608 = lut_tile_1_4_chanxy_out[70];
    assign wire_5610 = lut_tile_1_4_chanxy_out[71];
    assign wire_5611 = lut_tile_1_4_chanxy_out[72];
    assign wire_5612 = lut_tile_1_4_chanxy_out[73];
    assign wire_5614 = lut_tile_1_4_chanxy_out[74];
    assign wire_5616 = lut_tile_1_4_chanxy_out[75];
    assign wire_5618 = lut_tile_1_4_chanxy_out[76];
    assign wire_5619 = lut_tile_1_4_chanxy_out[77];
    assign wire_5620 = lut_tile_1_4_chanxy_out[78];
    assign wire_5622 = lut_tile_1_4_chanxy_out[79];
    assign wire_5624 = lut_tile_1_4_chanxy_out[80];
    assign wire_5626 = lut_tile_1_4_chanxy_out[81];
    assign wire_5627 = lut_tile_1_4_chanxy_out[82];
    assign wire_5628 = lut_tile_1_4_chanxy_out[83];
    assign wire_5630 = lut_tile_1_4_chanxy_out[84];
    assign wire_5632 = lut_tile_1_4_chanxy_out[85];
    assign wire_5634 = lut_tile_1_4_chanxy_out[86];
    assign wire_5635 = lut_tile_1_4_chanxy_out[87];
    assign wire_5636 = lut_tile_1_4_chanxy_out[88];
    assign wire_5638 = lut_tile_1_4_chanxy_out[89];
    assign wire_5640 = lut_tile_1_4_chanxy_out[90];
    assign wire_5642 = lut_tile_1_4_chanxy_out[91];
    assign wire_5643 = lut_tile_1_4_chanxy_out[92];
    assign wire_5644 = lut_tile_1_4_chanxy_out[93];
    assign wire_5646 = lut_tile_1_4_chanxy_out[94];
    assign wire_5648 = lut_tile_1_4_chanxy_out[95];
    assign wire_5650 = lut_tile_1_4_chanxy_out[96];
    assign wire_5651 = lut_tile_1_4_chanxy_out[97];
    assign wire_5652 = lut_tile_1_4_chanxy_out[98];
    assign wire_5654 = lut_tile_1_4_chanxy_out[99];
    assign wire_5656 = lut_tile_1_4_chanxy_out[100];
    assign wire_5658 = lut_tile_1_4_chanxy_out[101];
    assign wire_5659 = lut_tile_1_4_chanxy_out[102];
    assign wire_5660 = lut_tile_1_4_chanxy_out[103];
    assign wire_5662 = lut_tile_1_4_chanxy_out[104];
    assign wire_5664 = lut_tile_1_4_chanxy_out[105];
    assign wire_5666 = lut_tile_1_4_chanxy_out[106];
    assign wire_5667 = lut_tile_1_4_chanxy_out[107];
    assign wire_5668 = lut_tile_1_4_chanxy_out[108];
    assign wire_5670 = lut_tile_1_4_chanxy_out[109];
    assign wire_5672 = lut_tile_1_4_chanxy_out[110];
    assign wire_5674 = lut_tile_1_4_chanxy_out[111];
    assign wire_5675 = lut_tile_1_4_chanxy_out[112];
    assign wire_5676 = lut_tile_1_4_chanxy_out[113];
    assign wire_5678 = lut_tile_1_4_chanxy_out[114];
    assign wire_5680 = lut_tile_1_4_chanxy_out[115];
    assign wire_5682 = lut_tile_1_4_chanxy_out[116];
    assign wire_5683 = lut_tile_1_4_chanxy_out[117];
    assign wire_5684 = lut_tile_1_4_chanxy_out[118];
    assign wire_5686 = lut_tile_1_4_chanxy_out[119];
    assign wire_5688 = lut_tile_1_4_chanxy_out[120];
    assign wire_5690 = lut_tile_1_4_chanxy_out[121];
    assign wire_5691 = lut_tile_1_4_chanxy_out[122];
    assign wire_5692 = lut_tile_1_4_chanxy_out[123];
    assign wire_5694 = lut_tile_1_4_chanxy_out[124];
    assign wire_5696 = lut_tile_1_4_chanxy_out[125];
    assign wire_5698 = lut_tile_1_4_chanxy_out[126];
    assign wire_5699 = lut_tile_1_4_chanxy_out[127];
    assign wire_5700 = lut_tile_1_4_chanxy_out[128];
    assign wire_5702 = lut_tile_1_4_chanxy_out[129];
    assign wire_5704 = lut_tile_1_4_chanxy_out[130];
    assign wire_5706 = lut_tile_1_4_chanxy_out[131];
    assign wire_5707 = lut_tile_1_4_chanxy_out[132];
    assign wire_5708 = lut_tile_1_4_chanxy_out[133];
    assign wire_5710 = lut_tile_1_4_chanxy_out[134];
    assign wire_5712 = lut_tile_1_4_chanxy_out[135];
    assign wire_5714 = lut_tile_1_4_chanxy_out[136];
    assign wire_5715 = lut_tile_1_4_chanxy_out[137];
    assign wire_5716 = lut_tile_1_4_chanxy_out[138];
    assign wire_5718 = lut_tile_1_4_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_1_5_chanxy_in = {wire_2520, wire_2163, wire_6079, wire_2918, wire_2908, wire_2898, wire_2888, wire_2163, wire_2157, wire_2148, wire_1845, wire_2560, wire_2163, wire_2600, wire_2163, wire_2642, wire_2163, wire_2522, wire_2163, wire_6077, wire_2878, wire_2868, wire_2858, wire_2848, wire_2163, wire_2157, wire_2148, wire_1845, wire_2562, wire_2163, wire_2602, wire_2163, wire_2644, wire_2163, wire_2524, wire_2160, wire_6075, wire_2998, wire_2988, wire_2978, wire_2968, wire_2163, wire_2157, wire_2148, wire_1845, wire_2564, wire_2160, wire_2604, wire_2160, wire_2646, wire_2160, wire_2526, wire_2160, wire_6073, wire_2958, wire_2948, wire_2938, wire_2928, wire_2163, wire_2157, wire_2148, wire_1845, wire_2566, wire_2160, wire_2606, wire_2160, wire_2648, wire_2160, wire_2528, wire_2157, wire_6071, wire_2916, wire_2906, wire_2896, wire_2886, wire_2163, wire_2154, wire_2148, wire_1841, wire_2568, wire_2157, wire_2608, wire_2157, wire_2650, wire_2157, wire_2530, wire_2157, wire_6069, wire_2876, wire_2866, wire_2856, wire_2846, wire_2163, wire_2154, wire_2148, wire_1841, wire_2570, wire_2157, wire_2610, wire_2157, wire_2652, wire_2157, wire_2532, wire_2154, wire_6067, wire_2996, wire_2986, wire_2976, wire_2966, wire_2163, wire_2154, wire_2148, wire_1841, wire_2572, wire_2154, wire_2612, wire_2154, wire_2654, wire_2154, wire_2534, wire_2154, wire_6065, wire_2956, wire_2946, wire_2936, wire_2926, wire_2163, wire_2154, wire_2148, wire_1841, wire_2574, wire_2154, wire_2614, wire_2154, wire_2656, wire_2154, wire_2536, wire_2151, wire_6063, wire_2914, wire_2904, wire_2894, wire_2884, wire_2160, wire_2154, wire_2145, wire_1841, wire_2576, wire_2151, wire_2616, wire_2151, wire_2658, wire_2151, wire_2538, wire_2151, wire_6061, wire_2874, wire_2864, wire_2854, wire_2844, wire_2160, wire_2154, wire_2145, wire_1841, wire_2578, wire_2151, wire_2618, wire_2151, wire_2660, wire_2151, wire_2540, wire_2148, wire_6059, wire_2994, wire_2984, wire_2974, wire_2964, wire_2160, wire_2154, wire_2145, wire_1841, wire_2580, wire_2148, wire_2620, wire_2148, wire_2662, wire_2148, wire_2542, wire_2148, wire_6057, wire_2954, wire_2944, wire_2934, wire_2924, wire_2160, wire_2154, wire_2145, wire_1841, wire_2582, wire_2148, wire_2622, wire_2148, wire_2664, wire_2148, wire_2544, wire_2145, wire_6055, wire_2912, wire_2902, wire_2892, wire_2882, wire_2166, wire_2160, wire_2151, wire_2145, wire_1837, wire_2584, wire_2145, wire_2624, wire_2145, wire_2666, wire_2145, wire_2546, wire_2145, wire_6053, wire_2872, wire_2862, wire_2852, wire_2842, wire_2166, wire_2160, wire_2151, wire_2145, wire_1837, wire_2586, wire_2145, wire_2626, wire_2145, wire_2668, wire_2145, wire_2548, wire_1845, wire_6051, wire_2992, wire_2982, wire_2972, wire_2962, wire_2166, wire_2160, wire_2151, wire_2145, wire_1837, wire_2588, wire_1845, wire_2628, wire_1845, wire_2670, wire_1845, wire_2550, wire_1845, wire_6049, wire_2952, wire_2942, wire_2932, wire_2922, wire_2166, wire_2160, wire_2151, wire_2145, wire_1837, wire_2590, wire_1845, wire_2630, wire_1845, wire_2672, wire_1845, wire_2552, wire_1841, wire_6047, wire_2910, wire_2900, wire_2890, wire_2880, wire_2166, wire_2157, wire_2151, wire_1845, wire_1837, wire_2592, wire_1841, wire_2632, wire_1841, wire_2674, wire_1841, wire_2554, wire_1841, wire_6045, wire_2870, wire_2860, wire_2850, wire_2840, wire_2166, wire_2157, wire_2151, wire_1845, wire_1837, wire_2594, wire_1841, wire_2634, wire_1841, wire_2676, wire_1841, wire_2556, wire_2166, wire_1837, wire_6043, wire_2990, wire_2980, wire_2970, wire_2960, wire_2166, wire_2157, wire_2151, wire_1845, wire_1837, wire_2596, wire_2166, wire_1837, wire_2636, wire_2166, wire_1837, wire_2678, wire_2166, wire_1837, wire_2558, wire_2166, wire_1837, wire_6041, wire_2950, wire_2940, wire_2930, wire_2920, wire_2166, wire_2157, wire_2151, wire_1845, wire_1837, wire_2598, wire_2166, wire_1837, wire_2638, wire_2166, wire_1837, wire_2640, wire_2166, wire_1837, wire_6079, wire_6036, wire_5757, wire_5719, wire_5718, wire_5714, wire_5665, wire_5664, wire_5613, wire_5612, wire_2834, wire_1902, wire_1894, wire_6031, wire_6030, wire_5755, wire_5717, wire_5716, wire_5663, wire_5662, wire_5609, wire_5608, wire_5562, wire_2826, wire_1902, wire_1894, wire_6077, wire_6028, wire_5753, wire_5713, wire_5712, wire_5661, wire_5660, wire_5607, wire_5606, wire_5570, wire_2818, wire_1902, wire_1894, wire_5943, wire_5942, wire_5751, wire_5711, wire_5710, wire_5657, wire_5656, wire_5605, wire_5604, wire_5578, wire_2810, wire_1902, wire_1894, wire_5937, wire_5936, wire_5749, wire_5709, wire_5708, wire_5655, wire_5654, wire_5601, wire_5600, wire_5586, wire_2802, wire_1902, wire_1844, wire_5935, wire_5934, wire_5747, wire_5705, wire_5704, wire_5653, wire_5652, wire_5599, wire_5598, wire_5594, wire_2794, wire_1902, wire_1844, wire_6073, wire_6012, wire_5745, wire_5703, wire_5702, wire_5649, wire_5648, wire_5602, wire_5597, wire_5596, wire_2786, wire_1902, wire_1844, wire_6007, wire_6006, wire_5743, wire_5701, wire_5700, wire_5647, wire_5646, wire_5610, wire_5593, wire_5592, wire_2778, wire_1902, wire_1844, wire_6071, wire_6004, wire_5741, wire_5697, wire_5696, wire_5645, wire_5644, wire_5618, wire_5591, wire_5590, wire_2770, wire_1898, wire_1844, wire_5919, wire_5918, wire_5739, wire_5695, wire_5694, wire_5641, wire_5640, wire_5626, wire_5589, wire_5588, wire_2762, wire_1898, wire_1844, wire_5913, wire_5912, wire_1902, wire_5737, wire_5693, wire_5692, wire_5639, wire_5638, wire_5634, wire_5585, wire_5584, wire_2754, wire_1898, wire_1844, wire_5911, wire_5910, wire_1902, wire_5735, wire_5689, wire_5688, wire_5642, wire_5637, wire_5636, wire_5583, wire_5582, wire_2746, wire_1898, wire_1844, wire_6067, wire_5988, wire_1898, wire_5733, wire_5687, wire_5686, wire_5650, wire_5633, wire_5632, wire_5581, wire_5580, wire_2738, wire_1898, wire_1840, wire_5983, wire_5982, wire_1898, wire_5731, wire_5685, wire_5684, wire_5658, wire_5631, wire_5630, wire_5577, wire_5576, wire_2730, wire_1898, wire_1840, wire_6065, wire_5980, wire_1894, wire_5729, wire_5681, wire_5680, wire_5666, wire_5629, wire_5628, wire_5575, wire_5574, wire_2722, wire_1898, wire_1840, wire_5895, wire_5894, wire_1894, wire_5727, wire_5679, wire_5678, wire_5674, wire_5625, wire_5624, wire_5573, wire_5572, wire_2714, wire_1898, wire_1840, wire_5889, wire_5888, wire_1844, wire_5725, wire_5682, wire_5677, wire_5676, wire_5623, wire_5622, wire_5569, wire_5568, wire_2706, wire_1894, wire_1840, wire_5887, wire_5886, wire_1844, wire_5723, wire_5690, wire_5673, wire_5672, wire_5621, wire_5620, wire_5567, wire_5566, wire_2698, wire_1894, wire_1840, wire_6061, wire_5964, wire_1840, wire_5721, wire_5698, wire_5671, wire_5670, wire_5617, wire_5616, wire_5565, wire_5564, wire_2690, wire_1894, wire_1840, wire_5959, wire_5958, wire_1840, wire_5759, wire_5706, wire_5669, wire_5668, wire_5615, wire_5614, wire_5561, wire_5560, wire_2682, wire_1894, wire_1840, wire_6035, wire_6034, wire_5953, wire_5952, wire_5947, wire_5946, wire_6055, wire_5940, wire_6023, wire_6022, wire_6017, wire_6016, wire_6011, wire_6010, wire_5929, wire_5928, wire_5923, wire_5922, wire_6049, wire_5916, wire_5999, wire_5998, wire_1902, wire_5993, wire_5992, wire_1902, wire_5987, wire_5986, wire_1898, wire_5905, wire_5904, wire_1898, wire_5899, wire_5898, wire_1894, wire_6043, wire_5892, wire_1894, wire_5975, wire_5974, wire_1844, wire_5969, wire_5968, wire_1844, wire_5963, wire_5962, wire_1840, wire_5881, wire_5880, wire_1840, wire_6039, wire_6038, wire_5955, wire_5954, wire_5951, wire_5950, wire_5945, wire_5944, wire_6025, wire_6024, wire_6075, wire_6020, wire_6015, wire_6014, wire_5931, wire_5930, wire_5927, wire_5926, wire_5921, wire_5920, wire_6001, wire_6000, wire_1902, wire_6069, wire_5996, wire_1902, wire_5991, wire_5990, wire_1898, wire_5907, wire_5906, wire_1898, wire_5903, wire_5902, wire_1894, wire_5897, wire_5896, wire_1894, wire_5977, wire_5976, wire_1844, wire_6063, wire_5972, wire_1844, wire_5967, wire_5966, wire_1840, wire_5883, wire_5882, wire_1840, wire_6059, wire_5956, wire_6033, wire_6032, wire_6057, wire_5948, wire_6027, wire_6026, wire_5939, wire_5938, wire_6019, wire_6018, wire_6053, wire_5932, wire_6009, wire_6008, wire_6051, wire_5924, wire_6003, wire_6002, wire_5915, wire_5914, wire_1902, wire_5995, wire_5994, wire_1902, wire_6047, wire_5908, wire_1898, wire_5985, wire_5984, wire_1898, wire_6045, wire_5900, wire_1894, wire_5979, wire_5978, wire_1894, wire_5891, wire_5890, wire_1844, wire_5971, wire_5970, wire_1844, wire_6041, wire_5884, wire_1840, wire_5961, wire_5960, wire_1840};
    // CHNAXY TOTAL: 776
    assign wire_2841 = lut_tile_1_5_chanxy_out[0];
    assign wire_2843 = lut_tile_1_5_chanxy_out[1];
    assign wire_2845 = lut_tile_1_5_chanxy_out[2];
    assign wire_2847 = lut_tile_1_5_chanxy_out[3];
    assign wire_2849 = lut_tile_1_5_chanxy_out[4];
    assign wire_2851 = lut_tile_1_5_chanxy_out[5];
    assign wire_2853 = lut_tile_1_5_chanxy_out[6];
    assign wire_2855 = lut_tile_1_5_chanxy_out[7];
    assign wire_2857 = lut_tile_1_5_chanxy_out[8];
    assign wire_2859 = lut_tile_1_5_chanxy_out[9];
    assign wire_2861 = lut_tile_1_5_chanxy_out[10];
    assign wire_2863 = lut_tile_1_5_chanxy_out[11];
    assign wire_2865 = lut_tile_1_5_chanxy_out[12];
    assign wire_2867 = lut_tile_1_5_chanxy_out[13];
    assign wire_2869 = lut_tile_1_5_chanxy_out[14];
    assign wire_2871 = lut_tile_1_5_chanxy_out[15];
    assign wire_2873 = lut_tile_1_5_chanxy_out[16];
    assign wire_2875 = lut_tile_1_5_chanxy_out[17];
    assign wire_2877 = lut_tile_1_5_chanxy_out[18];
    assign wire_2879 = lut_tile_1_5_chanxy_out[19];
    assign wire_2881 = lut_tile_1_5_chanxy_out[20];
    assign wire_2883 = lut_tile_1_5_chanxy_out[21];
    assign wire_2885 = lut_tile_1_5_chanxy_out[22];
    assign wire_2887 = lut_tile_1_5_chanxy_out[23];
    assign wire_2889 = lut_tile_1_5_chanxy_out[24];
    assign wire_2891 = lut_tile_1_5_chanxy_out[25];
    assign wire_2893 = lut_tile_1_5_chanxy_out[26];
    assign wire_2895 = lut_tile_1_5_chanxy_out[27];
    assign wire_2897 = lut_tile_1_5_chanxy_out[28];
    assign wire_2899 = lut_tile_1_5_chanxy_out[29];
    assign wire_2901 = lut_tile_1_5_chanxy_out[30];
    assign wire_2903 = lut_tile_1_5_chanxy_out[31];
    assign wire_2905 = lut_tile_1_5_chanxy_out[32];
    assign wire_2907 = lut_tile_1_5_chanxy_out[33];
    assign wire_2909 = lut_tile_1_5_chanxy_out[34];
    assign wire_2911 = lut_tile_1_5_chanxy_out[35];
    assign wire_2913 = lut_tile_1_5_chanxy_out[36];
    assign wire_2915 = lut_tile_1_5_chanxy_out[37];
    assign wire_2917 = lut_tile_1_5_chanxy_out[38];
    assign wire_2919 = lut_tile_1_5_chanxy_out[39];
    assign wire_2921 = lut_tile_1_5_chanxy_out[40];
    assign wire_2923 = lut_tile_1_5_chanxy_out[41];
    assign wire_2925 = lut_tile_1_5_chanxy_out[42];
    assign wire_2927 = lut_tile_1_5_chanxy_out[43];
    assign wire_2929 = lut_tile_1_5_chanxy_out[44];
    assign wire_2931 = lut_tile_1_5_chanxy_out[45];
    assign wire_2933 = lut_tile_1_5_chanxy_out[46];
    assign wire_2935 = lut_tile_1_5_chanxy_out[47];
    assign wire_2937 = lut_tile_1_5_chanxy_out[48];
    assign wire_2939 = lut_tile_1_5_chanxy_out[49];
    assign wire_2941 = lut_tile_1_5_chanxy_out[50];
    assign wire_2943 = lut_tile_1_5_chanxy_out[51];
    assign wire_2945 = lut_tile_1_5_chanxy_out[52];
    assign wire_2947 = lut_tile_1_5_chanxy_out[53];
    assign wire_2949 = lut_tile_1_5_chanxy_out[54];
    assign wire_2951 = lut_tile_1_5_chanxy_out[55];
    assign wire_2953 = lut_tile_1_5_chanxy_out[56];
    assign wire_2955 = lut_tile_1_5_chanxy_out[57];
    assign wire_2957 = lut_tile_1_5_chanxy_out[58];
    assign wire_2959 = lut_tile_1_5_chanxy_out[59];
    assign wire_2960 = lut_tile_1_5_chanxy_out[60];
    assign wire_2961 = lut_tile_1_5_chanxy_out[61];
    assign wire_2962 = lut_tile_1_5_chanxy_out[62];
    assign wire_2963 = lut_tile_1_5_chanxy_out[63];
    assign wire_2964 = lut_tile_1_5_chanxy_out[64];
    assign wire_2965 = lut_tile_1_5_chanxy_out[65];
    assign wire_2966 = lut_tile_1_5_chanxy_out[66];
    assign wire_2967 = lut_tile_1_5_chanxy_out[67];
    assign wire_2968 = lut_tile_1_5_chanxy_out[68];
    assign wire_2969 = lut_tile_1_5_chanxy_out[69];
    assign wire_2970 = lut_tile_1_5_chanxy_out[70];
    assign wire_2971 = lut_tile_1_5_chanxy_out[71];
    assign wire_2972 = lut_tile_1_5_chanxy_out[72];
    assign wire_2973 = lut_tile_1_5_chanxy_out[73];
    assign wire_2974 = lut_tile_1_5_chanxy_out[74];
    assign wire_2975 = lut_tile_1_5_chanxy_out[75];
    assign wire_2976 = lut_tile_1_5_chanxy_out[76];
    assign wire_2977 = lut_tile_1_5_chanxy_out[77];
    assign wire_2978 = lut_tile_1_5_chanxy_out[78];
    assign wire_2979 = lut_tile_1_5_chanxy_out[79];
    assign wire_2980 = lut_tile_1_5_chanxy_out[80];
    assign wire_2981 = lut_tile_1_5_chanxy_out[81];
    assign wire_2982 = lut_tile_1_5_chanxy_out[82];
    assign wire_2983 = lut_tile_1_5_chanxy_out[83];
    assign wire_2984 = lut_tile_1_5_chanxy_out[84];
    assign wire_2985 = lut_tile_1_5_chanxy_out[85];
    assign wire_2986 = lut_tile_1_5_chanxy_out[86];
    assign wire_2987 = lut_tile_1_5_chanxy_out[87];
    assign wire_2988 = lut_tile_1_5_chanxy_out[88];
    assign wire_2989 = lut_tile_1_5_chanxy_out[89];
    assign wire_2990 = lut_tile_1_5_chanxy_out[90];
    assign wire_2991 = lut_tile_1_5_chanxy_out[91];
    assign wire_2992 = lut_tile_1_5_chanxy_out[92];
    assign wire_2993 = lut_tile_1_5_chanxy_out[93];
    assign wire_2994 = lut_tile_1_5_chanxy_out[94];
    assign wire_2995 = lut_tile_1_5_chanxy_out[95];
    assign wire_2996 = lut_tile_1_5_chanxy_out[96];
    assign wire_2997 = lut_tile_1_5_chanxy_out[97];
    assign wire_2998 = lut_tile_1_5_chanxy_out[98];
    assign wire_2999 = lut_tile_1_5_chanxy_out[99];
    assign wire_5880 = lut_tile_1_5_chanxy_out[100];
    assign wire_5882 = lut_tile_1_5_chanxy_out[101];
    assign wire_5884 = lut_tile_1_5_chanxy_out[102];
    assign wire_5885 = lut_tile_1_5_chanxy_out[103];
    assign wire_5886 = lut_tile_1_5_chanxy_out[104];
    assign wire_5888 = lut_tile_1_5_chanxy_out[105];
    assign wire_5890 = lut_tile_1_5_chanxy_out[106];
    assign wire_5892 = lut_tile_1_5_chanxy_out[107];
    assign wire_5893 = lut_tile_1_5_chanxy_out[108];
    assign wire_5894 = lut_tile_1_5_chanxy_out[109];
    assign wire_5896 = lut_tile_1_5_chanxy_out[110];
    assign wire_5898 = lut_tile_1_5_chanxy_out[111];
    assign wire_5900 = lut_tile_1_5_chanxy_out[112];
    assign wire_5901 = lut_tile_1_5_chanxy_out[113];
    assign wire_5902 = lut_tile_1_5_chanxy_out[114];
    assign wire_5904 = lut_tile_1_5_chanxy_out[115];
    assign wire_5906 = lut_tile_1_5_chanxy_out[116];
    assign wire_5908 = lut_tile_1_5_chanxy_out[117];
    assign wire_5909 = lut_tile_1_5_chanxy_out[118];
    assign wire_5910 = lut_tile_1_5_chanxy_out[119];
    assign wire_5912 = lut_tile_1_5_chanxy_out[120];
    assign wire_5914 = lut_tile_1_5_chanxy_out[121];
    assign wire_5916 = lut_tile_1_5_chanxy_out[122];
    assign wire_5917 = lut_tile_1_5_chanxy_out[123];
    assign wire_5918 = lut_tile_1_5_chanxy_out[124];
    assign wire_5920 = lut_tile_1_5_chanxy_out[125];
    assign wire_5922 = lut_tile_1_5_chanxy_out[126];
    assign wire_5924 = lut_tile_1_5_chanxy_out[127];
    assign wire_5925 = lut_tile_1_5_chanxy_out[128];
    assign wire_5926 = lut_tile_1_5_chanxy_out[129];
    assign wire_5928 = lut_tile_1_5_chanxy_out[130];
    assign wire_5930 = lut_tile_1_5_chanxy_out[131];
    assign wire_5932 = lut_tile_1_5_chanxy_out[132];
    assign wire_5933 = lut_tile_1_5_chanxy_out[133];
    assign wire_5934 = lut_tile_1_5_chanxy_out[134];
    assign wire_5936 = lut_tile_1_5_chanxy_out[135];
    assign wire_5938 = lut_tile_1_5_chanxy_out[136];
    assign wire_5940 = lut_tile_1_5_chanxy_out[137];
    assign wire_5941 = lut_tile_1_5_chanxy_out[138];
    assign wire_5942 = lut_tile_1_5_chanxy_out[139];
    assign wire_5944 = lut_tile_1_5_chanxy_out[140];
    assign wire_5946 = lut_tile_1_5_chanxy_out[141];
    assign wire_5948 = lut_tile_1_5_chanxy_out[142];
    assign wire_5949 = lut_tile_1_5_chanxy_out[143];
    assign wire_5950 = lut_tile_1_5_chanxy_out[144];
    assign wire_5952 = lut_tile_1_5_chanxy_out[145];
    assign wire_5954 = lut_tile_1_5_chanxy_out[146];
    assign wire_5956 = lut_tile_1_5_chanxy_out[147];
    assign wire_5957 = lut_tile_1_5_chanxy_out[148];
    assign wire_5958 = lut_tile_1_5_chanxy_out[149];
    assign wire_5960 = lut_tile_1_5_chanxy_out[150];
    assign wire_5962 = lut_tile_1_5_chanxy_out[151];
    assign wire_5964 = lut_tile_1_5_chanxy_out[152];
    assign wire_5965 = lut_tile_1_5_chanxy_out[153];
    assign wire_5966 = lut_tile_1_5_chanxy_out[154];
    assign wire_5968 = lut_tile_1_5_chanxy_out[155];
    assign wire_5970 = lut_tile_1_5_chanxy_out[156];
    assign wire_5972 = lut_tile_1_5_chanxy_out[157];
    assign wire_5973 = lut_tile_1_5_chanxy_out[158];
    assign wire_5974 = lut_tile_1_5_chanxy_out[159];
    assign wire_5976 = lut_tile_1_5_chanxy_out[160];
    assign wire_5978 = lut_tile_1_5_chanxy_out[161];
    assign wire_5980 = lut_tile_1_5_chanxy_out[162];
    assign wire_5981 = lut_tile_1_5_chanxy_out[163];
    assign wire_5982 = lut_tile_1_5_chanxy_out[164];
    assign wire_5984 = lut_tile_1_5_chanxy_out[165];
    assign wire_5986 = lut_tile_1_5_chanxy_out[166];
    assign wire_5988 = lut_tile_1_5_chanxy_out[167];
    assign wire_5989 = lut_tile_1_5_chanxy_out[168];
    assign wire_5990 = lut_tile_1_5_chanxy_out[169];
    assign wire_5992 = lut_tile_1_5_chanxy_out[170];
    assign wire_5994 = lut_tile_1_5_chanxy_out[171];
    assign wire_5996 = lut_tile_1_5_chanxy_out[172];
    assign wire_5997 = lut_tile_1_5_chanxy_out[173];
    assign wire_5998 = lut_tile_1_5_chanxy_out[174];
    assign wire_6000 = lut_tile_1_5_chanxy_out[175];
    assign wire_6002 = lut_tile_1_5_chanxy_out[176];
    assign wire_6004 = lut_tile_1_5_chanxy_out[177];
    assign wire_6005 = lut_tile_1_5_chanxy_out[178];
    assign wire_6006 = lut_tile_1_5_chanxy_out[179];
    assign wire_6008 = lut_tile_1_5_chanxy_out[180];
    assign wire_6010 = lut_tile_1_5_chanxy_out[181];
    assign wire_6012 = lut_tile_1_5_chanxy_out[182];
    assign wire_6013 = lut_tile_1_5_chanxy_out[183];
    assign wire_6014 = lut_tile_1_5_chanxy_out[184];
    assign wire_6016 = lut_tile_1_5_chanxy_out[185];
    assign wire_6018 = lut_tile_1_5_chanxy_out[186];
    assign wire_6020 = lut_tile_1_5_chanxy_out[187];
    assign wire_6021 = lut_tile_1_5_chanxy_out[188];
    assign wire_6022 = lut_tile_1_5_chanxy_out[189];
    assign wire_6024 = lut_tile_1_5_chanxy_out[190];
    assign wire_6026 = lut_tile_1_5_chanxy_out[191];
    assign wire_6028 = lut_tile_1_5_chanxy_out[192];
    assign wire_6029 = lut_tile_1_5_chanxy_out[193];
    assign wire_6030 = lut_tile_1_5_chanxy_out[194];
    assign wire_6032 = lut_tile_1_5_chanxy_out[195];
    assign wire_6034 = lut_tile_1_5_chanxy_out[196];
    assign wire_6036 = lut_tile_1_5_chanxy_out[197];
    assign wire_6037 = lut_tile_1_5_chanxy_out[198];
    assign wire_6038 = lut_tile_1_5_chanxy_out[199];
   // CHANXY OUT
    assign lut_tile_2_1_chanxy_in = {wire_4756, wire_2841, wire_2839, wire_2838, wire_2785, wire_2784, wire_2731, wire_2730, wire_2692, wire_771, wire_397, wire_4748, wire_2879, wire_2835, wire_2834, wire_2783, wire_2782, wire_2729, wire_2728, wire_2700, wire_771, wire_397, wire_4740, wire_2877, wire_2833, wire_2832, wire_2779, wire_2778, wire_2727, wire_2726, wire_2708, wire_771, wire_397, wire_4732, wire_2875, wire_2831, wire_2830, wire_2777, wire_2776, wire_2723, wire_2722, wire_2716, wire_771, wire_397, wire_4724, wire_2873, wire_2827, wire_2826, wire_2775, wire_2774, wire_2724, wire_2721, wire_2720, wire_771, wire_393, wire_4716, wire_2871, wire_2825, wire_2824, wire_2771, wire_2770, wire_2732, wire_2719, wire_2718, wire_771, wire_393, wire_4708, wire_2869, wire_2823, wire_2822, wire_2769, wire_2768, wire_2740, wire_2715, wire_2714, wire_771, wire_393, wire_4700, wire_2867, wire_2819, wire_2818, wire_2767, wire_2766, wire_2748, wire_2713, wire_2712, wire_771, wire_393, wire_4692, wire_2865, wire_2817, wire_2816, wire_2763, wire_2762, wire_2756, wire_2711, wire_2710, wire_767, wire_393, wire_4684, wire_2863, wire_2815, wire_2814, wire_2764, wire_2761, wire_2760, wire_2707, wire_2706, wire_767, wire_393, wire_4676, wire_2861, wire_2811, wire_2810, wire_2772, wire_2759, wire_2758, wire_2705, wire_2704, wire_767, wire_393, wire_4668, wire_2859, wire_2809, wire_2808, wire_2780, wire_2755, wire_2754, wire_2703, wire_2702, wire_767, wire_393, wire_4660, wire_2857, wire_2807, wire_2806, wire_2788, wire_2753, wire_2752, wire_2699, wire_2698, wire_767, wire_389, wire_4652, wire_2855, wire_2803, wire_2802, wire_2796, wire_2751, wire_2750, wire_2697, wire_2696, wire_767, wire_389, wire_4644, wire_2853, wire_2804, wire_2801, wire_2800, wire_2747, wire_2746, wire_2695, wire_2694, wire_767, wire_389, wire_4636, wire_2851, wire_2812, wire_2799, wire_2798, wire_2745, wire_2744, wire_2691, wire_2690, wire_767, wire_389, wire_4628, wire_2849, wire_2820, wire_2795, wire_2794, wire_2743, wire_2742, wire_2689, wire_2688, wire_397, wire_389, wire_4620, wire_2847, wire_2828, wire_2793, wire_2792, wire_2739, wire_2738, wire_2687, wire_2686, wire_397, wire_389, wire_4612, wire_2845, wire_2836, wire_2791, wire_2790, wire_2737, wire_2736, wire_2683, wire_2682, wire_397, wire_389, wire_4604, wire_2843, wire_2787, wire_2786, wire_2735, wire_2734, wire_2684, wire_2681, wire_2680, wire_397, wire_389, wire_4839, wire_3199, wire_3157, wire_3156, wire_3105, wire_3104, wire_3051, wire_3050, wire_3006, wire_771, wire_397, wire_4837, wire_3161, wire_3158, wire_3155, wire_3154, wire_3101, wire_3100, wire_3049, wire_3048, wire_771, wire_397, wire_4835, wire_3163, wire_3153, wire_3152, wire_3150, wire_3099, wire_3098, wire_3045, wire_3044, wire_771, wire_397, wire_4833, wire_3165, wire_3149, wire_3148, wire_3142, wire_3097, wire_3096, wire_3043, wire_3042, wire_771, wire_397, wire_4831, wire_3167, wire_3147, wire_3146, wire_3134, wire_3093, wire_3092, wire_3041, wire_3040, wire_771, wire_393, wire_4829, wire_3169, wire_3145, wire_3144, wire_3126, wire_3091, wire_3090, wire_3037, wire_3036, wire_771, wire_393, wire_4827, wire_3171, wire_3141, wire_3140, wire_3118, wire_3089, wire_3088, wire_3035, wire_3034, wire_771, wire_393, wire_4825, wire_3173, wire_3139, wire_3138, wire_3110, wire_3085, wire_3084, wire_3033, wire_3032, wire_771, wire_393, wire_4823, wire_3175, wire_3137, wire_3136, wire_3102, wire_3083, wire_3082, wire_3029, wire_3028, wire_767, wire_393, wire_4821, wire_3177, wire_3133, wire_3132, wire_3094, wire_3081, wire_3080, wire_3027, wire_3026, wire_767, wire_393, wire_4819, wire_3179, wire_3131, wire_3130, wire_3086, wire_3077, wire_3076, wire_3025, wire_3024, wire_767, wire_393, wire_4817, wire_3181, wire_3129, wire_3128, wire_3078, wire_3075, wire_3074, wire_3021, wire_3020, wire_767, wire_393, wire_4815, wire_3183, wire_3125, wire_3124, wire_3073, wire_3072, wire_3070, wire_3019, wire_3018, wire_767, wire_389, wire_4813, wire_3185, wire_3123, wire_3122, wire_3069, wire_3068, wire_3062, wire_3017, wire_3016, wire_767, wire_389, wire_4811, wire_3187, wire_3121, wire_3120, wire_3067, wire_3066, wire_3054, wire_3013, wire_3012, wire_767, wire_389, wire_4809, wire_3189, wire_3117, wire_3116, wire_3065, wire_3064, wire_3046, wire_3011, wire_3010, wire_767, wire_389, wire_4807, wire_3191, wire_3115, wire_3114, wire_3061, wire_3060, wire_3038, wire_3009, wire_3008, wire_397, wire_389, wire_4805, wire_3193, wire_3113, wire_3112, wire_3059, wire_3058, wire_3030, wire_3005, wire_3004, wire_397, wire_389, wire_4803, wire_3195, wire_3109, wire_3108, wire_3057, wire_3056, wire_3022, wire_3003, wire_3002, wire_397, wire_389, wire_4801, wire_3197, wire_3107, wire_3106, wire_3053, wire_3052, wire_3014, wire_3001, wire_3000, wire_397, wire_389, wire_4803, wire_4799, wire_4798, wire_4750, wire_4705, wire_4704, wire_4651, wire_4650, wire_3199, wire_454, wire_446, wire_4439, wire_4438, wire_4519, wire_4436, wire_4459, wire_4458, wire_4479, wire_4478, wire_4805, wire_4785, wire_4784, wire_4755, wire_4754, wire_4742, wire_4649, wire_4648, wire_3197, wire_454, wire_446, wire_4433, wire_4432, wire_4353, wire_4352, wire_4431, wire_4430, wire_4517, wire_4428, wire_4807, wire_4771, wire_4770, wire_4753, wire_4752, wire_4734, wire_4699, wire_4698, wire_3195, wire_454, wire_446, wire_4477, wire_4476, wire_4351, wire_4350, wire_4497, wire_4348, wire_4425, wire_4424, wire_4809, wire_4797, wire_4796, wire_4726, wire_4697, wire_4696, wire_4643, wire_4642, wire_3193, wire_454, wire_446, wire_4457, wire_4456, wire_4345, wire_4344, wire_4423, wire_4422, wire_4343, wire_4342, wire_4811, wire_4783, wire_4782, wire_4747, wire_4746, wire_4718, wire_4641, wire_4640, wire_3191, wire_454, wire_396, wire_4495, wire_4340, wire_4515, wire_4420, wire_4455, wire_4454, wire_4337, wire_4336, wire_4813, wire_4769, wire_4768, wire_4745, wire_4744, wire_4710, wire_4691, wire_4690, wire_3189, wire_454, wire_396, wire_4335, wire_4334, wire_4475, wire_4474, wire_4417, wire_4416, wire_4493, wire_4332, wire_4815, wire_4795, wire_4794, wire_4702, wire_4689, wire_4688, wire_4635, wire_4634, wire_3187, wire_454, wire_396, wire_4415, wire_4414, wire_4513, wire_4412, wire_4453, wire_4452, wire_4473, wire_4472, wire_4817, wire_4781, wire_4780, wire_4739, wire_4738, wire_4694, wire_4633, wire_4632, wire_3185, wire_454, wire_396, wire_4409, wire_4408, wire_4329, wire_4328, wire_4407, wire_4406, wire_4511, wire_4404, wire_4819, wire_4767, wire_4766, wire_4737, wire_4736, wire_4686, wire_4683, wire_4682, wire_3183, wire_450, wire_396, wire_4471, wire_4470, wire_4327, wire_4326, wire_4491, wire_4324, wire_4401, wire_4400, wire_4821, wire_4793, wire_4792, wire_4681, wire_4680, wire_4678, wire_4627, wire_4626, wire_3181, wire_450, wire_396, wire_4451, wire_4450, wire_4321, wire_4320, wire_4399, wire_4398, wire_4319, wire_4318, wire_4823, wire_4779, wire_4778, wire_4731, wire_4730, wire_4670, wire_4625, wire_4624, wire_3179, wire_450, wire_396, wire_4489, wire_4316, wire_454, wire_4509, wire_4396, wire_454, wire_4449, wire_4448, wire_454, wire_4313, wire_4312, wire_454, wire_4825, wire_4765, wire_4764, wire_4729, wire_4728, wire_4675, wire_4674, wire_4662, wire_3177, wire_450, wire_396, wire_4311, wire_4310, wire_454, wire_4469, wire_4468, wire_454, wire_4393, wire_4392, wire_454, wire_4487, wire_4308, wire_454, wire_4827, wire_4791, wire_4790, wire_4673, wire_4672, wire_4654, wire_4619, wire_4618, wire_3175, wire_450, wire_392, wire_4391, wire_4390, wire_450, wire_4507, wire_4388, wire_450, wire_4447, wire_4446, wire_450, wire_4467, wire_4466, wire_450, wire_4829, wire_4777, wire_4776, wire_4723, wire_4722, wire_4646, wire_4617, wire_4616, wire_3173, wire_450, wire_392, wire_4385, wire_4384, wire_450, wire_4305, wire_4304, wire_450, wire_4383, wire_4382, wire_450, wire_4505, wire_4380, wire_450, wire_4831, wire_4763, wire_4762, wire_4721, wire_4720, wire_4667, wire_4666, wire_4638, wire_3171, wire_450, wire_392, wire_4465, wire_4464, wire_446, wire_4303, wire_4302, wire_446, wire_4485, wire_4300, wire_446, wire_4377, wire_4376, wire_446, wire_4833, wire_4789, wire_4788, wire_4665, wire_4664, wire_4630, wire_4611, wire_4610, wire_3169, wire_450, wire_392, wire_4445, wire_4444, wire_446, wire_4297, wire_4296, wire_446, wire_4375, wire_4374, wire_446, wire_4295, wire_4294, wire_446, wire_4835, wire_4775, wire_4774, wire_4715, wire_4714, wire_4622, wire_4609, wire_4608, wire_3167, wire_446, wire_392, wire_4483, wire_4292, wire_396, wire_4503, wire_4372, wire_396, wire_4443, wire_4442, wire_396, wire_4289, wire_4288, wire_396, wire_4837, wire_4761, wire_4760, wire_4713, wire_4712, wire_4659, wire_4658, wire_4614, wire_3165, wire_446, wire_392, wire_4287, wire_4286, wire_396, wire_4463, wire_4462, wire_396, wire_4369, wire_4368, wire_396, wire_4481, wire_4284, wire_396, wire_4839, wire_4787, wire_4786, wire_4657, wire_4656, wire_4606, wire_4603, wire_4602, wire_3163, wire_446, wire_392, wire_4367, wire_4366, wire_392, wire_4501, wire_4364, wire_392, wire_4441, wire_4440, wire_392, wire_4461, wire_4460, wire_392, wire_4801, wire_4773, wire_4772, wire_4758, wire_4707, wire_4706, wire_4601, wire_4600, wire_3161, wire_446, wire_392, wire_4361, wire_4360, wire_392, wire_4281, wire_4280, wire_392, wire_4359, wire_4358, wire_392, wire_4499, wire_4356, wire_392};
    // CHNAXY TOTAL: 860
    assign wire_3000 = lut_tile_2_1_chanxy_out[0];
    assign wire_3002 = lut_tile_2_1_chanxy_out[1];
    assign wire_3004 = lut_tile_2_1_chanxy_out[2];
    assign wire_3006 = lut_tile_2_1_chanxy_out[3];
    assign wire_3007 = lut_tile_2_1_chanxy_out[4];
    assign wire_3008 = lut_tile_2_1_chanxy_out[5];
    assign wire_3010 = lut_tile_2_1_chanxy_out[6];
    assign wire_3012 = lut_tile_2_1_chanxy_out[7];
    assign wire_3014 = lut_tile_2_1_chanxy_out[8];
    assign wire_3015 = lut_tile_2_1_chanxy_out[9];
    assign wire_3016 = lut_tile_2_1_chanxy_out[10];
    assign wire_3018 = lut_tile_2_1_chanxy_out[11];
    assign wire_3020 = lut_tile_2_1_chanxy_out[12];
    assign wire_3022 = lut_tile_2_1_chanxy_out[13];
    assign wire_3023 = lut_tile_2_1_chanxy_out[14];
    assign wire_3024 = lut_tile_2_1_chanxy_out[15];
    assign wire_3026 = lut_tile_2_1_chanxy_out[16];
    assign wire_3028 = lut_tile_2_1_chanxy_out[17];
    assign wire_3030 = lut_tile_2_1_chanxy_out[18];
    assign wire_3031 = lut_tile_2_1_chanxy_out[19];
    assign wire_3032 = lut_tile_2_1_chanxy_out[20];
    assign wire_3034 = lut_tile_2_1_chanxy_out[21];
    assign wire_3036 = lut_tile_2_1_chanxy_out[22];
    assign wire_3038 = lut_tile_2_1_chanxy_out[23];
    assign wire_3039 = lut_tile_2_1_chanxy_out[24];
    assign wire_3040 = lut_tile_2_1_chanxy_out[25];
    assign wire_3042 = lut_tile_2_1_chanxy_out[26];
    assign wire_3044 = lut_tile_2_1_chanxy_out[27];
    assign wire_3046 = lut_tile_2_1_chanxy_out[28];
    assign wire_3047 = lut_tile_2_1_chanxy_out[29];
    assign wire_3048 = lut_tile_2_1_chanxy_out[30];
    assign wire_3050 = lut_tile_2_1_chanxy_out[31];
    assign wire_3052 = lut_tile_2_1_chanxy_out[32];
    assign wire_3054 = lut_tile_2_1_chanxy_out[33];
    assign wire_3055 = lut_tile_2_1_chanxy_out[34];
    assign wire_3056 = lut_tile_2_1_chanxy_out[35];
    assign wire_3058 = lut_tile_2_1_chanxy_out[36];
    assign wire_3060 = lut_tile_2_1_chanxy_out[37];
    assign wire_3062 = lut_tile_2_1_chanxy_out[38];
    assign wire_3063 = lut_tile_2_1_chanxy_out[39];
    assign wire_3064 = lut_tile_2_1_chanxy_out[40];
    assign wire_3066 = lut_tile_2_1_chanxy_out[41];
    assign wire_3068 = lut_tile_2_1_chanxy_out[42];
    assign wire_3070 = lut_tile_2_1_chanxy_out[43];
    assign wire_3071 = lut_tile_2_1_chanxy_out[44];
    assign wire_3072 = lut_tile_2_1_chanxy_out[45];
    assign wire_3074 = lut_tile_2_1_chanxy_out[46];
    assign wire_3076 = lut_tile_2_1_chanxy_out[47];
    assign wire_3078 = lut_tile_2_1_chanxy_out[48];
    assign wire_3079 = lut_tile_2_1_chanxy_out[49];
    assign wire_3080 = lut_tile_2_1_chanxy_out[50];
    assign wire_3082 = lut_tile_2_1_chanxy_out[51];
    assign wire_3084 = lut_tile_2_1_chanxy_out[52];
    assign wire_3086 = lut_tile_2_1_chanxy_out[53];
    assign wire_3087 = lut_tile_2_1_chanxy_out[54];
    assign wire_3088 = lut_tile_2_1_chanxy_out[55];
    assign wire_3090 = lut_tile_2_1_chanxy_out[56];
    assign wire_3092 = lut_tile_2_1_chanxy_out[57];
    assign wire_3094 = lut_tile_2_1_chanxy_out[58];
    assign wire_3095 = lut_tile_2_1_chanxy_out[59];
    assign wire_3096 = lut_tile_2_1_chanxy_out[60];
    assign wire_3098 = lut_tile_2_1_chanxy_out[61];
    assign wire_3100 = lut_tile_2_1_chanxy_out[62];
    assign wire_3102 = lut_tile_2_1_chanxy_out[63];
    assign wire_3103 = lut_tile_2_1_chanxy_out[64];
    assign wire_3104 = lut_tile_2_1_chanxy_out[65];
    assign wire_3106 = lut_tile_2_1_chanxy_out[66];
    assign wire_3108 = lut_tile_2_1_chanxy_out[67];
    assign wire_3110 = lut_tile_2_1_chanxy_out[68];
    assign wire_3111 = lut_tile_2_1_chanxy_out[69];
    assign wire_3112 = lut_tile_2_1_chanxy_out[70];
    assign wire_3114 = lut_tile_2_1_chanxy_out[71];
    assign wire_3116 = lut_tile_2_1_chanxy_out[72];
    assign wire_3118 = lut_tile_2_1_chanxy_out[73];
    assign wire_3119 = lut_tile_2_1_chanxy_out[74];
    assign wire_3120 = lut_tile_2_1_chanxy_out[75];
    assign wire_3122 = lut_tile_2_1_chanxy_out[76];
    assign wire_3124 = lut_tile_2_1_chanxy_out[77];
    assign wire_3126 = lut_tile_2_1_chanxy_out[78];
    assign wire_3127 = lut_tile_2_1_chanxy_out[79];
    assign wire_3128 = lut_tile_2_1_chanxy_out[80];
    assign wire_3130 = lut_tile_2_1_chanxy_out[81];
    assign wire_3132 = lut_tile_2_1_chanxy_out[82];
    assign wire_3134 = lut_tile_2_1_chanxy_out[83];
    assign wire_3135 = lut_tile_2_1_chanxy_out[84];
    assign wire_3136 = lut_tile_2_1_chanxy_out[85];
    assign wire_3138 = lut_tile_2_1_chanxy_out[86];
    assign wire_3140 = lut_tile_2_1_chanxy_out[87];
    assign wire_3142 = lut_tile_2_1_chanxy_out[88];
    assign wire_3143 = lut_tile_2_1_chanxy_out[89];
    assign wire_3144 = lut_tile_2_1_chanxy_out[90];
    assign wire_3146 = lut_tile_2_1_chanxy_out[91];
    assign wire_3148 = lut_tile_2_1_chanxy_out[92];
    assign wire_3150 = lut_tile_2_1_chanxy_out[93];
    assign wire_3151 = lut_tile_2_1_chanxy_out[94];
    assign wire_3152 = lut_tile_2_1_chanxy_out[95];
    assign wire_3154 = lut_tile_2_1_chanxy_out[96];
    assign wire_3156 = lut_tile_2_1_chanxy_out[97];
    assign wire_3158 = lut_tile_2_1_chanxy_out[98];
    assign wire_3159 = lut_tile_2_1_chanxy_out[99];
    assign wire_4607 = lut_tile_2_1_chanxy_out[100];
    assign wire_4615 = lut_tile_2_1_chanxy_out[101];
    assign wire_4623 = lut_tile_2_1_chanxy_out[102];
    assign wire_4631 = lut_tile_2_1_chanxy_out[103];
    assign wire_4639 = lut_tile_2_1_chanxy_out[104];
    assign wire_4647 = lut_tile_2_1_chanxy_out[105];
    assign wire_4655 = lut_tile_2_1_chanxy_out[106];
    assign wire_4663 = lut_tile_2_1_chanxy_out[107];
    assign wire_4671 = lut_tile_2_1_chanxy_out[108];
    assign wire_4679 = lut_tile_2_1_chanxy_out[109];
    assign wire_4687 = lut_tile_2_1_chanxy_out[110];
    assign wire_4695 = lut_tile_2_1_chanxy_out[111];
    assign wire_4703 = lut_tile_2_1_chanxy_out[112];
    assign wire_4711 = lut_tile_2_1_chanxy_out[113];
    assign wire_4719 = lut_tile_2_1_chanxy_out[114];
    assign wire_4727 = lut_tile_2_1_chanxy_out[115];
    assign wire_4735 = lut_tile_2_1_chanxy_out[116];
    assign wire_4743 = lut_tile_2_1_chanxy_out[117];
    assign wire_4751 = lut_tile_2_1_chanxy_out[118];
    assign wire_4759 = lut_tile_2_1_chanxy_out[119];
    assign wire_4760 = lut_tile_2_1_chanxy_out[120];
    assign wire_4762 = lut_tile_2_1_chanxy_out[121];
    assign wire_4764 = lut_tile_2_1_chanxy_out[122];
    assign wire_4766 = lut_tile_2_1_chanxy_out[123];
    assign wire_4768 = lut_tile_2_1_chanxy_out[124];
    assign wire_4770 = lut_tile_2_1_chanxy_out[125];
    assign wire_4772 = lut_tile_2_1_chanxy_out[126];
    assign wire_4774 = lut_tile_2_1_chanxy_out[127];
    assign wire_4776 = lut_tile_2_1_chanxy_out[128];
    assign wire_4778 = lut_tile_2_1_chanxy_out[129];
    assign wire_4780 = lut_tile_2_1_chanxy_out[130];
    assign wire_4782 = lut_tile_2_1_chanxy_out[131];
    assign wire_4784 = lut_tile_2_1_chanxy_out[132];
    assign wire_4786 = lut_tile_2_1_chanxy_out[133];
    assign wire_4788 = lut_tile_2_1_chanxy_out[134];
    assign wire_4790 = lut_tile_2_1_chanxy_out[135];
    assign wire_4792 = lut_tile_2_1_chanxy_out[136];
    assign wire_4794 = lut_tile_2_1_chanxy_out[137];
    assign wire_4796 = lut_tile_2_1_chanxy_out[138];
    assign wire_4798 = lut_tile_2_1_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_2_2_chanxy_in = {wire_5078, wire_2881, wire_2879, wire_2878, wire_2785, wire_2784, wire_2731, wire_2730, wire_2694, wire_1147, wire_773, wire_5070, wire_2919, wire_2865, wire_2864, wire_2835, wire_2834, wire_2729, wire_2728, wire_2702, wire_1147, wire_773, wire_5062, wire_2917, wire_2851, wire_2850, wire_2833, wire_2832, wire_2779, wire_2778, wire_2710, wire_1147, wire_773, wire_5054, wire_2915, wire_2877, wire_2876, wire_2777, wire_2776, wire_2723, wire_2722, wire_2718, wire_1147, wire_773, wire_5046, wire_2913, wire_2863, wire_2862, wire_2827, wire_2826, wire_2726, wire_2721, wire_2720, wire_1147, wire_769, wire_5038, wire_2911, wire_2849, wire_2848, wire_2825, wire_2824, wire_2771, wire_2770, wire_2734, wire_1147, wire_769, wire_5030, wire_2909, wire_2875, wire_2874, wire_2769, wire_2768, wire_2742, wire_2715, wire_2714, wire_1147, wire_769, wire_5022, wire_2907, wire_2861, wire_2860, wire_2819, wire_2818, wire_2750, wire_2713, wire_2712, wire_1147, wire_769, wire_5014, wire_2905, wire_2847, wire_2846, wire_2817, wire_2816, wire_2763, wire_2762, wire_2758, wire_1143, wire_769, wire_5006, wire_2903, wire_2873, wire_2872, wire_2766, wire_2761, wire_2760, wire_2707, wire_2706, wire_1143, wire_769, wire_4998, wire_2901, wire_2859, wire_2858, wire_2811, wire_2810, wire_2774, wire_2705, wire_2704, wire_1143, wire_769, wire_4990, wire_2899, wire_2845, wire_2844, wire_2809, wire_2808, wire_2782, wire_2755, wire_2754, wire_1143, wire_769, wire_4982, wire_2897, wire_2871, wire_2870, wire_2790, wire_2753, wire_2752, wire_2699, wire_2698, wire_1143, wire_765, wire_4974, wire_2895, wire_2857, wire_2856, wire_2803, wire_2802, wire_2798, wire_2697, wire_2696, wire_1143, wire_765, wire_4966, wire_2893, wire_2843, wire_2842, wire_2806, wire_2801, wire_2800, wire_2747, wire_2746, wire_1143, wire_765, wire_4958, wire_2891, wire_2869, wire_2868, wire_2814, wire_2745, wire_2744, wire_2691, wire_2690, wire_1143, wire_765, wire_4950, wire_2889, wire_2855, wire_2854, wire_2822, wire_2795, wire_2794, wire_2689, wire_2688, wire_773, wire_765, wire_4942, wire_2887, wire_2841, wire_2840, wire_2830, wire_2793, wire_2792, wire_2739, wire_2738, wire_773, wire_765, wire_4934, wire_2885, wire_2867, wire_2866, wire_2838, wire_2737, wire_2736, wire_2683, wire_2682, wire_773, wire_765, wire_4926, wire_2883, wire_2853, wire_2852, wire_2787, wire_2786, wire_2686, wire_2681, wire_2680, wire_773, wire_765, wire_5159, wire_3239, wire_3199, wire_3198, wire_3107, wire_3106, wire_3053, wire_3052, wire_3000, wire_1147, wire_773, wire_5157, wire_3201, wire_3185, wire_3184, wire_3157, wire_3156, wire_3152, wire_3051, wire_3050, wire_1147, wire_773, wire_5155, wire_3203, wire_3171, wire_3170, wire_3155, wire_3154, wire_3144, wire_3101, wire_3100, wire_1147, wire_773, wire_5153, wire_3205, wire_3197, wire_3196, wire_3136, wire_3099, wire_3098, wire_3045, wire_3044, wire_1147, wire_773, wire_5151, wire_3207, wire_3183, wire_3182, wire_3149, wire_3148, wire_3128, wire_3043, wire_3042, wire_1147, wire_769, wire_5149, wire_3209, wire_3169, wire_3168, wire_3147, wire_3146, wire_3120, wire_3093, wire_3092, wire_1147, wire_769, wire_5147, wire_3211, wire_3195, wire_3194, wire_3112, wire_3091, wire_3090, wire_3037, wire_3036, wire_1147, wire_769, wire_5145, wire_3213, wire_3181, wire_3180, wire_3141, wire_3140, wire_3104, wire_3035, wire_3034, wire_1147, wire_769, wire_5143, wire_3215, wire_3167, wire_3166, wire_3139, wire_3138, wire_3096, wire_3085, wire_3084, wire_1143, wire_769, wire_5141, wire_3217, wire_3193, wire_3192, wire_3088, wire_3083, wire_3082, wire_3029, wire_3028, wire_1143, wire_769, wire_5139, wire_3219, wire_3179, wire_3178, wire_3133, wire_3132, wire_3080, wire_3027, wire_3026, wire_1143, wire_769, wire_5137, wire_3221, wire_3165, wire_3164, wire_3131, wire_3130, wire_3077, wire_3076, wire_3072, wire_1143, wire_769, wire_5135, wire_3223, wire_3191, wire_3190, wire_3075, wire_3074, wire_3064, wire_3021, wire_3020, wire_1143, wire_765, wire_5133, wire_3225, wire_3177, wire_3176, wire_3125, wire_3124, wire_3056, wire_3019, wire_3018, wire_1143, wire_765, wire_5131, wire_3227, wire_3163, wire_3162, wire_3123, wire_3122, wire_3069, wire_3068, wire_3048, wire_1143, wire_765, wire_5129, wire_3229, wire_3189, wire_3188, wire_3067, wire_3066, wire_3040, wire_3013, wire_3012, wire_1143, wire_765, wire_5127, wire_3231, wire_3175, wire_3174, wire_3117, wire_3116, wire_3032, wire_3011, wire_3010, wire_773, wire_765, wire_5125, wire_3233, wire_3161, wire_3160, wire_3115, wire_3114, wire_3061, wire_3060, wire_3024, wire_773, wire_765, wire_5123, wire_3235, wire_3187, wire_3186, wire_3059, wire_3058, wire_3016, wire_3005, wire_3004, wire_773, wire_765, wire_5121, wire_3237, wire_3173, wire_3172, wire_3109, wire_3108, wire_3008, wire_3003, wire_3002, wire_773, wire_765, wire_4837, wire_4799, wire_4798, wire_4758, wire_4705, wire_4704, wire_4651, wire_4650, wire_3158, wire_830, wire_822, wire_4835, wire_4785, wire_4784, wire_4755, wire_4754, wire_4649, wire_4648, wire_4606, wire_3150, wire_830, wire_822, wire_4833, wire_4771, wire_4770, wire_4753, wire_4752, wire_4699, wire_4698, wire_4614, wire_3142, wire_830, wire_822, wire_4831, wire_4797, wire_4796, wire_4697, wire_4696, wire_4643, wire_4642, wire_4622, wire_3134, wire_830, wire_822, wire_4829, wire_4783, wire_4782, wire_4747, wire_4746, wire_4641, wire_4640, wire_4630, wire_3126, wire_830, wire_772, wire_4827, wire_4769, wire_4768, wire_4745, wire_4744, wire_4691, wire_4690, wire_4638, wire_3118, wire_830, wire_772, wire_4825, wire_4795, wire_4794, wire_4689, wire_4688, wire_4646, wire_4635, wire_4634, wire_3110, wire_830, wire_772, wire_4823, wire_4781, wire_4780, wire_4739, wire_4738, wire_4654, wire_4633, wire_4632, wire_3102, wire_830, wire_772, wire_4821, wire_4767, wire_4766, wire_4737, wire_4736, wire_4683, wire_4682, wire_4662, wire_3094, wire_826, wire_772, wire_4819, wire_4793, wire_4792, wire_4681, wire_4680, wire_4670, wire_4627, wire_4626, wire_3086, wire_826, wire_772, wire_4817, wire_4779, wire_4778, wire_4731, wire_4730, wire_4678, wire_4625, wire_4624, wire_3078, wire_826, wire_772, wire_4815, wire_4765, wire_4764, wire_4729, wire_4728, wire_4686, wire_4675, wire_4674, wire_3070, wire_826, wire_772, wire_4813, wire_4791, wire_4790, wire_4694, wire_4673, wire_4672, wire_4619, wire_4618, wire_3062, wire_826, wire_768, wire_4811, wire_4777, wire_4776, wire_4723, wire_4722, wire_4702, wire_4617, wire_4616, wire_3054, wire_826, wire_768, wire_4809, wire_4763, wire_4762, wire_4721, wire_4720, wire_4710, wire_4667, wire_4666, wire_3046, wire_826, wire_768, wire_4807, wire_4789, wire_4788, wire_4718, wire_4665, wire_4664, wire_4611, wire_4610, wire_3038, wire_826, wire_768, wire_4805, wire_4775, wire_4774, wire_4726, wire_4715, wire_4714, wire_4609, wire_4608, wire_3030, wire_822, wire_768, wire_4803, wire_4761, wire_4760, wire_4734, wire_4713, wire_4712, wire_4659, wire_4658, wire_3022, wire_822, wire_768, wire_4801, wire_4787, wire_4786, wire_4742, wire_4657, wire_4656, wire_4603, wire_4602, wire_3014, wire_822, wire_768, wire_4839, wire_4773, wire_4772, wire_4750, wire_4707, wire_4706, wire_4601, wire_4600, wire_3006, wire_822, wire_768, wire_5123, wire_5119, wire_5118, wire_5064, wire_5027, wire_5026, wire_4973, wire_4972, wire_3239, wire_830, wire_822, wire_5125, wire_5105, wire_5104, wire_5077, wire_5076, wire_5056, wire_4971, wire_4970, wire_3237, wire_830, wire_822, wire_5127, wire_5091, wire_5090, wire_5075, wire_5074, wire_5048, wire_5021, wire_5020, wire_3235, wire_830, wire_822, wire_5129, wire_5117, wire_5116, wire_5040, wire_5019, wire_5018, wire_4965, wire_4964, wire_3233, wire_830, wire_822, wire_5131, wire_5103, wire_5102, wire_5069, wire_5068, wire_5032, wire_4963, wire_4962, wire_3231, wire_830, wire_772, wire_5133, wire_5089, wire_5088, wire_5067, wire_5066, wire_5024, wire_5013, wire_5012, wire_3229, wire_830, wire_772, wire_5135, wire_5115, wire_5114, wire_5016, wire_5011, wire_5010, wire_4957, wire_4956, wire_3227, wire_830, wire_772, wire_5137, wire_5101, wire_5100, wire_5061, wire_5060, wire_5008, wire_4955, wire_4954, wire_3225, wire_830, wire_772, wire_5139, wire_5087, wire_5086, wire_5059, wire_5058, wire_5005, wire_5004, wire_5000, wire_3223, wire_826, wire_772, wire_5141, wire_5113, wire_5112, wire_5003, wire_5002, wire_4992, wire_4949, wire_4948, wire_3221, wire_826, wire_772, wire_5143, wire_5099, wire_5098, wire_5053, wire_5052, wire_4984, wire_4947, wire_4946, wire_3219, wire_826, wire_772, wire_5145, wire_5085, wire_5084, wire_5051, wire_5050, wire_4997, wire_4996, wire_4976, wire_3217, wire_826, wire_772, wire_5147, wire_5111, wire_5110, wire_4995, wire_4994, wire_4968, wire_4941, wire_4940, wire_3215, wire_826, wire_768, wire_5149, wire_5097, wire_5096, wire_5045, wire_5044, wire_4960, wire_4939, wire_4938, wire_3213, wire_826, wire_768, wire_5151, wire_5083, wire_5082, wire_5043, wire_5042, wire_4989, wire_4988, wire_4952, wire_3211, wire_826, wire_768, wire_5153, wire_5109, wire_5108, wire_4987, wire_4986, wire_4944, wire_4933, wire_4932, wire_3209, wire_826, wire_768, wire_5155, wire_5095, wire_5094, wire_5037, wire_5036, wire_4936, wire_4931, wire_4930, wire_3207, wire_822, wire_768, wire_5157, wire_5081, wire_5080, wire_5035, wire_5034, wire_4981, wire_4980, wire_4928, wire_3205, wire_822, wire_768, wire_5159, wire_5107, wire_5106, wire_4979, wire_4978, wire_4925, wire_4924, wire_4920, wire_3203, wire_822, wire_768, wire_5121, wire_5093, wire_5092, wire_5072, wire_5029, wire_5028, wire_4923, wire_4922, wire_3201, wire_822, wire_768};
    // CHNAXY TOTAL: 880
    assign wire_3001 = lut_tile_2_2_chanxy_out[0];
    assign wire_3009 = lut_tile_2_2_chanxy_out[1];
    assign wire_3017 = lut_tile_2_2_chanxy_out[2];
    assign wire_3025 = lut_tile_2_2_chanxy_out[3];
    assign wire_3033 = lut_tile_2_2_chanxy_out[4];
    assign wire_3041 = lut_tile_2_2_chanxy_out[5];
    assign wire_3049 = lut_tile_2_2_chanxy_out[6];
    assign wire_3057 = lut_tile_2_2_chanxy_out[7];
    assign wire_3065 = lut_tile_2_2_chanxy_out[8];
    assign wire_3073 = lut_tile_2_2_chanxy_out[9];
    assign wire_3081 = lut_tile_2_2_chanxy_out[10];
    assign wire_3089 = lut_tile_2_2_chanxy_out[11];
    assign wire_3097 = lut_tile_2_2_chanxy_out[12];
    assign wire_3105 = lut_tile_2_2_chanxy_out[13];
    assign wire_3113 = lut_tile_2_2_chanxy_out[14];
    assign wire_3121 = lut_tile_2_2_chanxy_out[15];
    assign wire_3129 = lut_tile_2_2_chanxy_out[16];
    assign wire_3137 = lut_tile_2_2_chanxy_out[17];
    assign wire_3145 = lut_tile_2_2_chanxy_out[18];
    assign wire_3153 = lut_tile_2_2_chanxy_out[19];
    assign wire_3160 = lut_tile_2_2_chanxy_out[20];
    assign wire_3162 = lut_tile_2_2_chanxy_out[21];
    assign wire_3164 = lut_tile_2_2_chanxy_out[22];
    assign wire_3166 = lut_tile_2_2_chanxy_out[23];
    assign wire_3168 = lut_tile_2_2_chanxy_out[24];
    assign wire_3170 = lut_tile_2_2_chanxy_out[25];
    assign wire_3172 = lut_tile_2_2_chanxy_out[26];
    assign wire_3174 = lut_tile_2_2_chanxy_out[27];
    assign wire_3176 = lut_tile_2_2_chanxy_out[28];
    assign wire_3178 = lut_tile_2_2_chanxy_out[29];
    assign wire_3180 = lut_tile_2_2_chanxy_out[30];
    assign wire_3182 = lut_tile_2_2_chanxy_out[31];
    assign wire_3184 = lut_tile_2_2_chanxy_out[32];
    assign wire_3186 = lut_tile_2_2_chanxy_out[33];
    assign wire_3188 = lut_tile_2_2_chanxy_out[34];
    assign wire_3190 = lut_tile_2_2_chanxy_out[35];
    assign wire_3192 = lut_tile_2_2_chanxy_out[36];
    assign wire_3194 = lut_tile_2_2_chanxy_out[37];
    assign wire_3196 = lut_tile_2_2_chanxy_out[38];
    assign wire_3198 = lut_tile_2_2_chanxy_out[39];
    assign wire_4921 = lut_tile_2_2_chanxy_out[40];
    assign wire_4929 = lut_tile_2_2_chanxy_out[41];
    assign wire_4937 = lut_tile_2_2_chanxy_out[42];
    assign wire_4945 = lut_tile_2_2_chanxy_out[43];
    assign wire_4953 = lut_tile_2_2_chanxy_out[44];
    assign wire_4961 = lut_tile_2_2_chanxy_out[45];
    assign wire_4969 = lut_tile_2_2_chanxy_out[46];
    assign wire_4977 = lut_tile_2_2_chanxy_out[47];
    assign wire_4985 = lut_tile_2_2_chanxy_out[48];
    assign wire_4993 = lut_tile_2_2_chanxy_out[49];
    assign wire_5001 = lut_tile_2_2_chanxy_out[50];
    assign wire_5009 = lut_tile_2_2_chanxy_out[51];
    assign wire_5017 = lut_tile_2_2_chanxy_out[52];
    assign wire_5025 = lut_tile_2_2_chanxy_out[53];
    assign wire_5033 = lut_tile_2_2_chanxy_out[54];
    assign wire_5041 = lut_tile_2_2_chanxy_out[55];
    assign wire_5049 = lut_tile_2_2_chanxy_out[56];
    assign wire_5057 = lut_tile_2_2_chanxy_out[57];
    assign wire_5065 = lut_tile_2_2_chanxy_out[58];
    assign wire_5073 = lut_tile_2_2_chanxy_out[59];
    assign wire_5080 = lut_tile_2_2_chanxy_out[60];
    assign wire_5082 = lut_tile_2_2_chanxy_out[61];
    assign wire_5084 = lut_tile_2_2_chanxy_out[62];
    assign wire_5086 = lut_tile_2_2_chanxy_out[63];
    assign wire_5088 = lut_tile_2_2_chanxy_out[64];
    assign wire_5090 = lut_tile_2_2_chanxy_out[65];
    assign wire_5092 = lut_tile_2_2_chanxy_out[66];
    assign wire_5094 = lut_tile_2_2_chanxy_out[67];
    assign wire_5096 = lut_tile_2_2_chanxy_out[68];
    assign wire_5098 = lut_tile_2_2_chanxy_out[69];
    assign wire_5100 = lut_tile_2_2_chanxy_out[70];
    assign wire_5102 = lut_tile_2_2_chanxy_out[71];
    assign wire_5104 = lut_tile_2_2_chanxy_out[72];
    assign wire_5106 = lut_tile_2_2_chanxy_out[73];
    assign wire_5108 = lut_tile_2_2_chanxy_out[74];
    assign wire_5110 = lut_tile_2_2_chanxy_out[75];
    assign wire_5112 = lut_tile_2_2_chanxy_out[76];
    assign wire_5114 = lut_tile_2_2_chanxy_out[77];
    assign wire_5116 = lut_tile_2_2_chanxy_out[78];
    assign wire_5118 = lut_tile_2_2_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_2_3_chanxy_in = {wire_5392, wire_2921, wire_2919, wire_2918, wire_2853, wire_2852, wire_2787, wire_2786, wire_2688, wire_1523, wire_1149, wire_5384, wire_2959, wire_2905, wire_2904, wire_2879, wire_2878, wire_2731, wire_2730, wire_2696, wire_1523, wire_1149, wire_5376, wire_2957, wire_2891, wire_2890, wire_2865, wire_2864, wire_2835, wire_2834, wire_2704, wire_1523, wire_1149, wire_5368, wire_2955, wire_2917, wire_2916, wire_2851, wire_2850, wire_2779, wire_2778, wire_2712, wire_1523, wire_1149, wire_5360, wire_2953, wire_2903, wire_2902, wire_2877, wire_2876, wire_2723, wire_2722, wire_2720, wire_1523, wire_1145, wire_5352, wire_2951, wire_2889, wire_2888, wire_2863, wire_2862, wire_2827, wire_2826, wire_2728, wire_1523, wire_1145, wire_5344, wire_2949, wire_2915, wire_2914, wire_2849, wire_2848, wire_2771, wire_2770, wire_2736, wire_1523, wire_1145, wire_5336, wire_2947, wire_2901, wire_2900, wire_2875, wire_2874, wire_2744, wire_2715, wire_2714, wire_1523, wire_1145, wire_5328, wire_2945, wire_2887, wire_2886, wire_2861, wire_2860, wire_2819, wire_2818, wire_2752, wire_1519, wire_1145, wire_5320, wire_2943, wire_2913, wire_2912, wire_2847, wire_2846, wire_2763, wire_2762, wire_2760, wire_1519, wire_1145, wire_5312, wire_2941, wire_2899, wire_2898, wire_2873, wire_2872, wire_2768, wire_2707, wire_2706, wire_1519, wire_1145, wire_5304, wire_2939, wire_2885, wire_2884, wire_2859, wire_2858, wire_2811, wire_2810, wire_2776, wire_1519, wire_1145, wire_5296, wire_2937, wire_2911, wire_2910, wire_2845, wire_2844, wire_2784, wire_2755, wire_2754, wire_1519, wire_1141, wire_5288, wire_2935, wire_2897, wire_2896, wire_2871, wire_2870, wire_2792, wire_2699, wire_2698, wire_1519, wire_1141, wire_5280, wire_2933, wire_2883, wire_2882, wire_2857, wire_2856, wire_2803, wire_2802, wire_2800, wire_1519, wire_1141, wire_5272, wire_2931, wire_2909, wire_2908, wire_2843, wire_2842, wire_2808, wire_2747, wire_2746, wire_1519, wire_1141, wire_5264, wire_2929, wire_2895, wire_2894, wire_2869, wire_2868, wire_2816, wire_2691, wire_2690, wire_1149, wire_1141, wire_5256, wire_2927, wire_2881, wire_2880, wire_2855, wire_2854, wire_2824, wire_2795, wire_2794, wire_1149, wire_1141, wire_5248, wire_2925, wire_2907, wire_2906, wire_2841, wire_2840, wire_2832, wire_2739, wire_2738, wire_1149, wire_1141, wire_5240, wire_2923, wire_2893, wire_2892, wire_2867, wire_2866, wire_2683, wire_2682, wire_2680, wire_1149, wire_1141, wire_5479, wire_3279, wire_3227, wire_3226, wire_3199, wire_3198, wire_3053, wire_3052, wire_3002, wire_1523, wire_1149, wire_5477, wire_3241, wire_3213, wire_3212, wire_3185, wire_3184, wire_3157, wire_3156, wire_3154, wire_1523, wire_1149, wire_5475, wire_3243, wire_3239, wire_3238, wire_3171, wire_3170, wire_3146, wire_3101, wire_3100, wire_1523, wire_1149, wire_5473, wire_3245, wire_3225, wire_3224, wire_3197, wire_3196, wire_3138, wire_3045, wire_3044, wire_1523, wire_1149, wire_5471, wire_3247, wire_3211, wire_3210, wire_3183, wire_3182, wire_3149, wire_3148, wire_3130, wire_1523, wire_1145, wire_5469, wire_3249, wire_3237, wire_3236, wire_3169, wire_3168, wire_3122, wire_3093, wire_3092, wire_1523, wire_1145, wire_5467, wire_3251, wire_3223, wire_3222, wire_3195, wire_3194, wire_3114, wire_3037, wire_3036, wire_1523, wire_1145, wire_5465, wire_3253, wire_3209, wire_3208, wire_3181, wire_3180, wire_3141, wire_3140, wire_3106, wire_1523, wire_1145, wire_5463, wire_3255, wire_3235, wire_3234, wire_3167, wire_3166, wire_3098, wire_3085, wire_3084, wire_1519, wire_1145, wire_5461, wire_3257, wire_3221, wire_3220, wire_3193, wire_3192, wire_3090, wire_3029, wire_3028, wire_1519, wire_1145, wire_5459, wire_3259, wire_3207, wire_3206, wire_3179, wire_3178, wire_3133, wire_3132, wire_3082, wire_1519, wire_1145, wire_5457, wire_3261, wire_3233, wire_3232, wire_3165, wire_3164, wire_3077, wire_3076, wire_3074, wire_1519, wire_1145, wire_5455, wire_3263, wire_3219, wire_3218, wire_3191, wire_3190, wire_3066, wire_3021, wire_3020, wire_1519, wire_1141, wire_5453, wire_3265, wire_3205, wire_3204, wire_3177, wire_3176, wire_3125, wire_3124, wire_3058, wire_1519, wire_1141, wire_5451, wire_3267, wire_3231, wire_3230, wire_3163, wire_3162, wire_3069, wire_3068, wire_3050, wire_1519, wire_1141, wire_5449, wire_3269, wire_3217, wire_3216, wire_3189, wire_3188, wire_3042, wire_3013, wire_3012, wire_1519, wire_1141, wire_5447, wire_3271, wire_3203, wire_3202, wire_3175, wire_3174, wire_3117, wire_3116, wire_3034, wire_1149, wire_1141, wire_5445, wire_3273, wire_3229, wire_3228, wire_3161, wire_3160, wire_3061, wire_3060, wire_3026, wire_1149, wire_1141, wire_5443, wire_3275, wire_3215, wire_3214, wire_3187, wire_3186, wire_3018, wire_3005, wire_3004, wire_1149, wire_1141, wire_5441, wire_3277, wire_3201, wire_3200, wire_3173, wire_3172, wire_3109, wire_3108, wire_3010, wire_1149, wire_1141, wire_5157, wire_5119, wire_5118, wire_5072, wire_5027, wire_5026, wire_4973, wire_4972, wire_3152, wire_1206, wire_1198, wire_5155, wire_5105, wire_5104, wire_5077, wire_5076, wire_4971, wire_4970, wire_4920, wire_3144, wire_1206, wire_1198, wire_5153, wire_5091, wire_5090, wire_5075, wire_5074, wire_5021, wire_5020, wire_4928, wire_3136, wire_1206, wire_1198, wire_5151, wire_5117, wire_5116, wire_5019, wire_5018, wire_4965, wire_4964, wire_4936, wire_3128, wire_1206, wire_1198, wire_5149, wire_5103, wire_5102, wire_5069, wire_5068, wire_4963, wire_4962, wire_4944, wire_3120, wire_1206, wire_1148, wire_5147, wire_5089, wire_5088, wire_5067, wire_5066, wire_5013, wire_5012, wire_4952, wire_3112, wire_1206, wire_1148, wire_5145, wire_5115, wire_5114, wire_5011, wire_5010, wire_4960, wire_4957, wire_4956, wire_3104, wire_1206, wire_1148, wire_5143, wire_5101, wire_5100, wire_5061, wire_5060, wire_4968, wire_4955, wire_4954, wire_3096, wire_1206, wire_1148, wire_5141, wire_5087, wire_5086, wire_5059, wire_5058, wire_5005, wire_5004, wire_4976, wire_3088, wire_1202, wire_1148, wire_5139, wire_5113, wire_5112, wire_5003, wire_5002, wire_4984, wire_4949, wire_4948, wire_3080, wire_1202, wire_1148, wire_5137, wire_5099, wire_5098, wire_5053, wire_5052, wire_4992, wire_4947, wire_4946, wire_3072, wire_1202, wire_1148, wire_5135, wire_5085, wire_5084, wire_5051, wire_5050, wire_5000, wire_4997, wire_4996, wire_3064, wire_1202, wire_1148, wire_5133, wire_5111, wire_5110, wire_5008, wire_4995, wire_4994, wire_4941, wire_4940, wire_3056, wire_1202, wire_1144, wire_5131, wire_5097, wire_5096, wire_5045, wire_5044, wire_5016, wire_4939, wire_4938, wire_3048, wire_1202, wire_1144, wire_5129, wire_5083, wire_5082, wire_5043, wire_5042, wire_5024, wire_4989, wire_4988, wire_3040, wire_1202, wire_1144, wire_5127, wire_5109, wire_5108, wire_5032, wire_4987, wire_4986, wire_4933, wire_4932, wire_3032, wire_1202, wire_1144, wire_5125, wire_5095, wire_5094, wire_5040, wire_5037, wire_5036, wire_4931, wire_4930, wire_3024, wire_1198, wire_1144, wire_5123, wire_5081, wire_5080, wire_5048, wire_5035, wire_5034, wire_4981, wire_4980, wire_3016, wire_1198, wire_1144, wire_5121, wire_5107, wire_5106, wire_5056, wire_4979, wire_4978, wire_4925, wire_4924, wire_3008, wire_1198, wire_1144, wire_5159, wire_5093, wire_5092, wire_5064, wire_5029, wire_5028, wire_4923, wire_4922, wire_3000, wire_1198, wire_1144, wire_5443, wire_5427, wire_5426, wire_5399, wire_5398, wire_5386, wire_5293, wire_5292, wire_3279, wire_1206, wire_1198, wire_5445, wire_5413, wire_5412, wire_5397, wire_5396, wire_5378, wire_5343, wire_5342, wire_3277, wire_1206, wire_1198, wire_5447, wire_5439, wire_5438, wire_5370, wire_5341, wire_5340, wire_5287, wire_5286, wire_3275, wire_1206, wire_1198, wire_5449, wire_5425, wire_5424, wire_5391, wire_5390, wire_5362, wire_5285, wire_5284, wire_3273, wire_1206, wire_1198, wire_5451, wire_5411, wire_5410, wire_5389, wire_5388, wire_5354, wire_5335, wire_5334, wire_3271, wire_1206, wire_1148, wire_5453, wire_5437, wire_5436, wire_5346, wire_5333, wire_5332, wire_5279, wire_5278, wire_3269, wire_1206, wire_1148, wire_5455, wire_5423, wire_5422, wire_5383, wire_5382, wire_5338, wire_5277, wire_5276, wire_3267, wire_1206, wire_1148, wire_5457, wire_5409, wire_5408, wire_5381, wire_5380, wire_5330, wire_5327, wire_5326, wire_3265, wire_1206, wire_1148, wire_5459, wire_5435, wire_5434, wire_5325, wire_5324, wire_5322, wire_5271, wire_5270, wire_3263, wire_1202, wire_1148, wire_5461, wire_5421, wire_5420, wire_5375, wire_5374, wire_5314, wire_5269, wire_5268, wire_3261, wire_1202, wire_1148, wire_5463, wire_5407, wire_5406, wire_5373, wire_5372, wire_5319, wire_5318, wire_5306, wire_3259, wire_1202, wire_1148, wire_5465, wire_5433, wire_5432, wire_5317, wire_5316, wire_5298, wire_5263, wire_5262, wire_3257, wire_1202, wire_1148, wire_5467, wire_5419, wire_5418, wire_5367, wire_5366, wire_5290, wire_5261, wire_5260, wire_3255, wire_1202, wire_1144, wire_5469, wire_5405, wire_5404, wire_5365, wire_5364, wire_5311, wire_5310, wire_5282, wire_3253, wire_1202, wire_1144, wire_5471, wire_5431, wire_5430, wire_5309, wire_5308, wire_5274, wire_5255, wire_5254, wire_3251, wire_1202, wire_1144, wire_5473, wire_5417, wire_5416, wire_5359, wire_5358, wire_5266, wire_5253, wire_5252, wire_3249, wire_1202, wire_1144, wire_5475, wire_5403, wire_5402, wire_5357, wire_5356, wire_5303, wire_5302, wire_5258, wire_3247, wire_1198, wire_1144, wire_5477, wire_5429, wire_5428, wire_5301, wire_5300, wire_5250, wire_5247, wire_5246, wire_3245, wire_1198, wire_1144, wire_5479, wire_5415, wire_5414, wire_5351, wire_5350, wire_5245, wire_5244, wire_5242, wire_3243, wire_1198, wire_1144, wire_5441, wire_5401, wire_5400, wire_5394, wire_5349, wire_5348, wire_5295, wire_5294, wire_3241, wire_1198, wire_1144};
    // CHNAXY TOTAL: 880
    assign wire_3003 = lut_tile_2_3_chanxy_out[0];
    assign wire_3011 = lut_tile_2_3_chanxy_out[1];
    assign wire_3019 = lut_tile_2_3_chanxy_out[2];
    assign wire_3027 = lut_tile_2_3_chanxy_out[3];
    assign wire_3035 = lut_tile_2_3_chanxy_out[4];
    assign wire_3043 = lut_tile_2_3_chanxy_out[5];
    assign wire_3051 = lut_tile_2_3_chanxy_out[6];
    assign wire_3059 = lut_tile_2_3_chanxy_out[7];
    assign wire_3067 = lut_tile_2_3_chanxy_out[8];
    assign wire_3075 = lut_tile_2_3_chanxy_out[9];
    assign wire_3083 = lut_tile_2_3_chanxy_out[10];
    assign wire_3091 = lut_tile_2_3_chanxy_out[11];
    assign wire_3099 = lut_tile_2_3_chanxy_out[12];
    assign wire_3107 = lut_tile_2_3_chanxy_out[13];
    assign wire_3115 = lut_tile_2_3_chanxy_out[14];
    assign wire_3123 = lut_tile_2_3_chanxy_out[15];
    assign wire_3131 = lut_tile_2_3_chanxy_out[16];
    assign wire_3139 = lut_tile_2_3_chanxy_out[17];
    assign wire_3147 = lut_tile_2_3_chanxy_out[18];
    assign wire_3155 = lut_tile_2_3_chanxy_out[19];
    assign wire_3200 = lut_tile_2_3_chanxy_out[20];
    assign wire_3202 = lut_tile_2_3_chanxy_out[21];
    assign wire_3204 = lut_tile_2_3_chanxy_out[22];
    assign wire_3206 = lut_tile_2_3_chanxy_out[23];
    assign wire_3208 = lut_tile_2_3_chanxy_out[24];
    assign wire_3210 = lut_tile_2_3_chanxy_out[25];
    assign wire_3212 = lut_tile_2_3_chanxy_out[26];
    assign wire_3214 = lut_tile_2_3_chanxy_out[27];
    assign wire_3216 = lut_tile_2_3_chanxy_out[28];
    assign wire_3218 = lut_tile_2_3_chanxy_out[29];
    assign wire_3220 = lut_tile_2_3_chanxy_out[30];
    assign wire_3222 = lut_tile_2_3_chanxy_out[31];
    assign wire_3224 = lut_tile_2_3_chanxy_out[32];
    assign wire_3226 = lut_tile_2_3_chanxy_out[33];
    assign wire_3228 = lut_tile_2_3_chanxy_out[34];
    assign wire_3230 = lut_tile_2_3_chanxy_out[35];
    assign wire_3232 = lut_tile_2_3_chanxy_out[36];
    assign wire_3234 = lut_tile_2_3_chanxy_out[37];
    assign wire_3236 = lut_tile_2_3_chanxy_out[38];
    assign wire_3238 = lut_tile_2_3_chanxy_out[39];
    assign wire_5243 = lut_tile_2_3_chanxy_out[40];
    assign wire_5251 = lut_tile_2_3_chanxy_out[41];
    assign wire_5259 = lut_tile_2_3_chanxy_out[42];
    assign wire_5267 = lut_tile_2_3_chanxy_out[43];
    assign wire_5275 = lut_tile_2_3_chanxy_out[44];
    assign wire_5283 = lut_tile_2_3_chanxy_out[45];
    assign wire_5291 = lut_tile_2_3_chanxy_out[46];
    assign wire_5299 = lut_tile_2_3_chanxy_out[47];
    assign wire_5307 = lut_tile_2_3_chanxy_out[48];
    assign wire_5315 = lut_tile_2_3_chanxy_out[49];
    assign wire_5323 = lut_tile_2_3_chanxy_out[50];
    assign wire_5331 = lut_tile_2_3_chanxy_out[51];
    assign wire_5339 = lut_tile_2_3_chanxy_out[52];
    assign wire_5347 = lut_tile_2_3_chanxy_out[53];
    assign wire_5355 = lut_tile_2_3_chanxy_out[54];
    assign wire_5363 = lut_tile_2_3_chanxy_out[55];
    assign wire_5371 = lut_tile_2_3_chanxy_out[56];
    assign wire_5379 = lut_tile_2_3_chanxy_out[57];
    assign wire_5387 = lut_tile_2_3_chanxy_out[58];
    assign wire_5395 = lut_tile_2_3_chanxy_out[59];
    assign wire_5400 = lut_tile_2_3_chanxy_out[60];
    assign wire_5402 = lut_tile_2_3_chanxy_out[61];
    assign wire_5404 = lut_tile_2_3_chanxy_out[62];
    assign wire_5406 = lut_tile_2_3_chanxy_out[63];
    assign wire_5408 = lut_tile_2_3_chanxy_out[64];
    assign wire_5410 = lut_tile_2_3_chanxy_out[65];
    assign wire_5412 = lut_tile_2_3_chanxy_out[66];
    assign wire_5414 = lut_tile_2_3_chanxy_out[67];
    assign wire_5416 = lut_tile_2_3_chanxy_out[68];
    assign wire_5418 = lut_tile_2_3_chanxy_out[69];
    assign wire_5420 = lut_tile_2_3_chanxy_out[70];
    assign wire_5422 = lut_tile_2_3_chanxy_out[71];
    assign wire_5424 = lut_tile_2_3_chanxy_out[72];
    assign wire_5426 = lut_tile_2_3_chanxy_out[73];
    assign wire_5428 = lut_tile_2_3_chanxy_out[74];
    assign wire_5430 = lut_tile_2_3_chanxy_out[75];
    assign wire_5432 = lut_tile_2_3_chanxy_out[76];
    assign wire_5434 = lut_tile_2_3_chanxy_out[77];
    assign wire_5436 = lut_tile_2_3_chanxy_out[78];
    assign wire_5438 = lut_tile_2_3_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_2_4_chanxy_in = {wire_5714, wire_2961, wire_2947, wire_2946, wire_2919, wire_2918, wire_2853, wire_2852, wire_2690, wire_1899, wire_1525, wire_5706, wire_2999, wire_2933, wire_2932, wire_2905, wire_2904, wire_2879, wire_2878, wire_2698, wire_1899, wire_1525, wire_5698, wire_2997, wire_2959, wire_2958, wire_2891, wire_2890, wire_2865, wire_2864, wire_2706, wire_1899, wire_1525, wire_5690, wire_2995, wire_2945, wire_2944, wire_2917, wire_2916, wire_2851, wire_2850, wire_2714, wire_1899, wire_1525, wire_5682, wire_2993, wire_2931, wire_2930, wire_2903, wire_2902, wire_2877, wire_2876, wire_2722, wire_1899, wire_1521, wire_5674, wire_2991, wire_2957, wire_2956, wire_2889, wire_2888, wire_2863, wire_2862, wire_2730, wire_1899, wire_1521, wire_5666, wire_2989, wire_2943, wire_2942, wire_2915, wire_2914, wire_2849, wire_2848, wire_2738, wire_1899, wire_1521, wire_5658, wire_2987, wire_2929, wire_2928, wire_2901, wire_2900, wire_2875, wire_2874, wire_2746, wire_1899, wire_1521, wire_5650, wire_2985, wire_2955, wire_2954, wire_2887, wire_2886, wire_2861, wire_2860, wire_2754, wire_1895, wire_1521, wire_5642, wire_2983, wire_2941, wire_2940, wire_2913, wire_2912, wire_2847, wire_2846, wire_2762, wire_1895, wire_1521, wire_5634, wire_2981, wire_2927, wire_2926, wire_2899, wire_2898, wire_2873, wire_2872, wire_2770, wire_1895, wire_1521, wire_5626, wire_2979, wire_2953, wire_2952, wire_2885, wire_2884, wire_2859, wire_2858, wire_2778, wire_1895, wire_1521, wire_5618, wire_2977, wire_2939, wire_2938, wire_2911, wire_2910, wire_2845, wire_2844, wire_2786, wire_1895, wire_1517, wire_5610, wire_2975, wire_2925, wire_2924, wire_2897, wire_2896, wire_2871, wire_2870, wire_2794, wire_1895, wire_1517, wire_5602, wire_2973, wire_2951, wire_2950, wire_2883, wire_2882, wire_2857, wire_2856, wire_2802, wire_1895, wire_1517, wire_5594, wire_2971, wire_2937, wire_2936, wire_2909, wire_2908, wire_2843, wire_2842, wire_2810, wire_1895, wire_1517, wire_5586, wire_2969, wire_2923, wire_2922, wire_2895, wire_2894, wire_2869, wire_2868, wire_2818, wire_1525, wire_1517, wire_5578, wire_2967, wire_2949, wire_2948, wire_2881, wire_2880, wire_2855, wire_2854, wire_2826, wire_1525, wire_1517, wire_5570, wire_2965, wire_2935, wire_2934, wire_2907, wire_2906, wire_2841, wire_2840, wire_2834, wire_1525, wire_1517, wire_5562, wire_2963, wire_2921, wire_2920, wire_2893, wire_2892, wire_2867, wire_2866, wire_2682, wire_1525, wire_1517, wire_5799, wire_3319, wire_3253, wire_3252, wire_3227, wire_3226, wire_3199, wire_3198, wire_3004, wire_1899, wire_1525, wire_5797, wire_3281, wire_3279, wire_3278, wire_3213, wire_3212, wire_3185, wire_3184, wire_3156, wire_1899, wire_1525, wire_5795, wire_3283, wire_3265, wire_3264, wire_3239, wire_3238, wire_3171, wire_3170, wire_3148, wire_1899, wire_1525, wire_5793, wire_3285, wire_3251, wire_3250, wire_3225, wire_3224, wire_3197, wire_3196, wire_3140, wire_1899, wire_1525, wire_5791, wire_3287, wire_3277, wire_3276, wire_3211, wire_3210, wire_3183, wire_3182, wire_3132, wire_1899, wire_1521, wire_5789, wire_3289, wire_3263, wire_3262, wire_3237, wire_3236, wire_3169, wire_3168, wire_3124, wire_1899, wire_1521, wire_5787, wire_3291, wire_3249, wire_3248, wire_3223, wire_3222, wire_3195, wire_3194, wire_3116, wire_1899, wire_1521, wire_5785, wire_3293, wire_3275, wire_3274, wire_3209, wire_3208, wire_3181, wire_3180, wire_3108, wire_1899, wire_1521, wire_5783, wire_3295, wire_3261, wire_3260, wire_3235, wire_3234, wire_3167, wire_3166, wire_3100, wire_1895, wire_1521, wire_5781, wire_3297, wire_3247, wire_3246, wire_3221, wire_3220, wire_3193, wire_3192, wire_3092, wire_1895, wire_1521, wire_5779, wire_3299, wire_3273, wire_3272, wire_3207, wire_3206, wire_3179, wire_3178, wire_3084, wire_1895, wire_1521, wire_5777, wire_3301, wire_3259, wire_3258, wire_3233, wire_3232, wire_3165, wire_3164, wire_3076, wire_1895, wire_1521, wire_5775, wire_3303, wire_3245, wire_3244, wire_3219, wire_3218, wire_3191, wire_3190, wire_3068, wire_1895, wire_1517, wire_5773, wire_3305, wire_3271, wire_3270, wire_3205, wire_3204, wire_3177, wire_3176, wire_3060, wire_1895, wire_1517, wire_5771, wire_3307, wire_3257, wire_3256, wire_3231, wire_3230, wire_3163, wire_3162, wire_3052, wire_1895, wire_1517, wire_5769, wire_3309, wire_3243, wire_3242, wire_3217, wire_3216, wire_3189, wire_3188, wire_3044, wire_1895, wire_1517, wire_5767, wire_3311, wire_3269, wire_3268, wire_3203, wire_3202, wire_3175, wire_3174, wire_3036, wire_1525, wire_1517, wire_5765, wire_3313, wire_3255, wire_3254, wire_3229, wire_3228, wire_3161, wire_3160, wire_3028, wire_1525, wire_1517, wire_5763, wire_3315, wire_3241, wire_3240, wire_3215, wire_3214, wire_3187, wire_3186, wire_3020, wire_1525, wire_1517, wire_5761, wire_3317, wire_3267, wire_3266, wire_3201, wire_3200, wire_3173, wire_3172, wire_3012, wire_1525, wire_1517, wire_5477, wire_5427, wire_5426, wire_5399, wire_5398, wire_5394, wire_5293, wire_5292, wire_3154, wire_1582, wire_1574, wire_5475, wire_5413, wire_5412, wire_5397, wire_5396, wire_5343, wire_5342, wire_5242, wire_3146, wire_1582, wire_1574, wire_5473, wire_5439, wire_5438, wire_5341, wire_5340, wire_5287, wire_5286, wire_5250, wire_3138, wire_1582, wire_1574, wire_5471, wire_5425, wire_5424, wire_5391, wire_5390, wire_5285, wire_5284, wire_5258, wire_3130, wire_1582, wire_1574, wire_5469, wire_5411, wire_5410, wire_5389, wire_5388, wire_5335, wire_5334, wire_5266, wire_3122, wire_1582, wire_1524, wire_5467, wire_5437, wire_5436, wire_5333, wire_5332, wire_5279, wire_5278, wire_5274, wire_3114, wire_1582, wire_1524, wire_5465, wire_5423, wire_5422, wire_5383, wire_5382, wire_5282, wire_5277, wire_5276, wire_3106, wire_1582, wire_1524, wire_5463, wire_5409, wire_5408, wire_5381, wire_5380, wire_5327, wire_5326, wire_5290, wire_3098, wire_1582, wire_1524, wire_5461, wire_5435, wire_5434, wire_5325, wire_5324, wire_5298, wire_5271, wire_5270, wire_3090, wire_1578, wire_1524, wire_5459, wire_5421, wire_5420, wire_5375, wire_5374, wire_5306, wire_5269, wire_5268, wire_3082, wire_1578, wire_1524, wire_5457, wire_5407, wire_5406, wire_5373, wire_5372, wire_5319, wire_5318, wire_5314, wire_3074, wire_1578, wire_1524, wire_5455, wire_5433, wire_5432, wire_5322, wire_5317, wire_5316, wire_5263, wire_5262, wire_3066, wire_1578, wire_1524, wire_5453, wire_5419, wire_5418, wire_5367, wire_5366, wire_5330, wire_5261, wire_5260, wire_3058, wire_1578, wire_1520, wire_5451, wire_5405, wire_5404, wire_5365, wire_5364, wire_5338, wire_5311, wire_5310, wire_3050, wire_1578, wire_1520, wire_5449, wire_5431, wire_5430, wire_5346, wire_5309, wire_5308, wire_5255, wire_5254, wire_3042, wire_1578, wire_1520, wire_5447, wire_5417, wire_5416, wire_5359, wire_5358, wire_5354, wire_5253, wire_5252, wire_3034, wire_1578, wire_1520, wire_5445, wire_5403, wire_5402, wire_5362, wire_5357, wire_5356, wire_5303, wire_5302, wire_3026, wire_1574, wire_1520, wire_5443, wire_5429, wire_5428, wire_5370, wire_5301, wire_5300, wire_5247, wire_5246, wire_3018, wire_1574, wire_1520, wire_5441, wire_5415, wire_5414, wire_5378, wire_5351, wire_5350, wire_5245, wire_5244, wire_3010, wire_1574, wire_1520, wire_5479, wire_5401, wire_5400, wire_5386, wire_5349, wire_5348, wire_5295, wire_5294, wire_3002, wire_1574, wire_1520, wire_5763, wire_5733, wire_5732, wire_5719, wire_5718, wire_5708, wire_5665, wire_5664, wire_3319, wire_1582, wire_1574, wire_5765, wire_5759, wire_5758, wire_5700, wire_5663, wire_5662, wire_5609, wire_5608, wire_3317, wire_1582, wire_1574, wire_5767, wire_5745, wire_5744, wire_5713, wire_5712, wire_5692, wire_5607, wire_5606, wire_3315, wire_1582, wire_1574, wire_5769, wire_5731, wire_5730, wire_5711, wire_5710, wire_5684, wire_5657, wire_5656, wire_3313, wire_1582, wire_1574, wire_5771, wire_5757, wire_5756, wire_5676, wire_5655, wire_5654, wire_5601, wire_5600, wire_3311, wire_1582, wire_1524, wire_5773, wire_5743, wire_5742, wire_5705, wire_5704, wire_5668, wire_5599, wire_5598, wire_3309, wire_1582, wire_1524, wire_5775, wire_5729, wire_5728, wire_5703, wire_5702, wire_5660, wire_5649, wire_5648, wire_3307, wire_1582, wire_1524, wire_5777, wire_5755, wire_5754, wire_5652, wire_5647, wire_5646, wire_5593, wire_5592, wire_3305, wire_1582, wire_1524, wire_5779, wire_5741, wire_5740, wire_5697, wire_5696, wire_5644, wire_5591, wire_5590, wire_3303, wire_1578, wire_1524, wire_5781, wire_5727, wire_5726, wire_5695, wire_5694, wire_5641, wire_5640, wire_5636, wire_3301, wire_1578, wire_1524, wire_5783, wire_5753, wire_5752, wire_5639, wire_5638, wire_5628, wire_5585, wire_5584, wire_3299, wire_1578, wire_1524, wire_5785, wire_5739, wire_5738, wire_5689, wire_5688, wire_5620, wire_5583, wire_5582, wire_3297, wire_1578, wire_1524, wire_5787, wire_5725, wire_5724, wire_5687, wire_5686, wire_5633, wire_5632, wire_5612, wire_3295, wire_1578, wire_1520, wire_5789, wire_5751, wire_5750, wire_5631, wire_5630, wire_5604, wire_5577, wire_5576, wire_3293, wire_1578, wire_1520, wire_5791, wire_5737, wire_5736, wire_5681, wire_5680, wire_5596, wire_5575, wire_5574, wire_3291, wire_1578, wire_1520, wire_5793, wire_5723, wire_5722, wire_5679, wire_5678, wire_5625, wire_5624, wire_5588, wire_3289, wire_1578, wire_1520, wire_5795, wire_5749, wire_5748, wire_5623, wire_5622, wire_5580, wire_5569, wire_5568, wire_3287, wire_1574, wire_1520, wire_5797, wire_5735, wire_5734, wire_5673, wire_5672, wire_5572, wire_5567, wire_5566, wire_3285, wire_1574, wire_1520, wire_5799, wire_5721, wire_5720, wire_5671, wire_5670, wire_5617, wire_5616, wire_5564, wire_3283, wire_1574, wire_1520, wire_5761, wire_5747, wire_5746, wire_5716, wire_5615, wire_5614, wire_5561, wire_5560, wire_3281, wire_1574, wire_1520};
    // CHNAXY TOTAL: 880
    assign wire_3005 = lut_tile_2_4_chanxy_out[0];
    assign wire_3013 = lut_tile_2_4_chanxy_out[1];
    assign wire_3021 = lut_tile_2_4_chanxy_out[2];
    assign wire_3029 = lut_tile_2_4_chanxy_out[3];
    assign wire_3037 = lut_tile_2_4_chanxy_out[4];
    assign wire_3045 = lut_tile_2_4_chanxy_out[5];
    assign wire_3053 = lut_tile_2_4_chanxy_out[6];
    assign wire_3061 = lut_tile_2_4_chanxy_out[7];
    assign wire_3069 = lut_tile_2_4_chanxy_out[8];
    assign wire_3077 = lut_tile_2_4_chanxy_out[9];
    assign wire_3085 = lut_tile_2_4_chanxy_out[10];
    assign wire_3093 = lut_tile_2_4_chanxy_out[11];
    assign wire_3101 = lut_tile_2_4_chanxy_out[12];
    assign wire_3109 = lut_tile_2_4_chanxy_out[13];
    assign wire_3117 = lut_tile_2_4_chanxy_out[14];
    assign wire_3125 = lut_tile_2_4_chanxy_out[15];
    assign wire_3133 = lut_tile_2_4_chanxy_out[16];
    assign wire_3141 = lut_tile_2_4_chanxy_out[17];
    assign wire_3149 = lut_tile_2_4_chanxy_out[18];
    assign wire_3157 = lut_tile_2_4_chanxy_out[19];
    assign wire_3240 = lut_tile_2_4_chanxy_out[20];
    assign wire_3242 = lut_tile_2_4_chanxy_out[21];
    assign wire_3244 = lut_tile_2_4_chanxy_out[22];
    assign wire_3246 = lut_tile_2_4_chanxy_out[23];
    assign wire_3248 = lut_tile_2_4_chanxy_out[24];
    assign wire_3250 = lut_tile_2_4_chanxy_out[25];
    assign wire_3252 = lut_tile_2_4_chanxy_out[26];
    assign wire_3254 = lut_tile_2_4_chanxy_out[27];
    assign wire_3256 = lut_tile_2_4_chanxy_out[28];
    assign wire_3258 = lut_tile_2_4_chanxy_out[29];
    assign wire_3260 = lut_tile_2_4_chanxy_out[30];
    assign wire_3262 = lut_tile_2_4_chanxy_out[31];
    assign wire_3264 = lut_tile_2_4_chanxy_out[32];
    assign wire_3266 = lut_tile_2_4_chanxy_out[33];
    assign wire_3268 = lut_tile_2_4_chanxy_out[34];
    assign wire_3270 = lut_tile_2_4_chanxy_out[35];
    assign wire_3272 = lut_tile_2_4_chanxy_out[36];
    assign wire_3274 = lut_tile_2_4_chanxy_out[37];
    assign wire_3276 = lut_tile_2_4_chanxy_out[38];
    assign wire_3278 = lut_tile_2_4_chanxy_out[39];
    assign wire_5565 = lut_tile_2_4_chanxy_out[40];
    assign wire_5573 = lut_tile_2_4_chanxy_out[41];
    assign wire_5581 = lut_tile_2_4_chanxy_out[42];
    assign wire_5589 = lut_tile_2_4_chanxy_out[43];
    assign wire_5597 = lut_tile_2_4_chanxy_out[44];
    assign wire_5605 = lut_tile_2_4_chanxy_out[45];
    assign wire_5613 = lut_tile_2_4_chanxy_out[46];
    assign wire_5621 = lut_tile_2_4_chanxy_out[47];
    assign wire_5629 = lut_tile_2_4_chanxy_out[48];
    assign wire_5637 = lut_tile_2_4_chanxy_out[49];
    assign wire_5645 = lut_tile_2_4_chanxy_out[50];
    assign wire_5653 = lut_tile_2_4_chanxy_out[51];
    assign wire_5661 = lut_tile_2_4_chanxy_out[52];
    assign wire_5669 = lut_tile_2_4_chanxy_out[53];
    assign wire_5677 = lut_tile_2_4_chanxy_out[54];
    assign wire_5685 = lut_tile_2_4_chanxy_out[55];
    assign wire_5693 = lut_tile_2_4_chanxy_out[56];
    assign wire_5701 = lut_tile_2_4_chanxy_out[57];
    assign wire_5709 = lut_tile_2_4_chanxy_out[58];
    assign wire_5717 = lut_tile_2_4_chanxy_out[59];
    assign wire_5720 = lut_tile_2_4_chanxy_out[60];
    assign wire_5722 = lut_tile_2_4_chanxy_out[61];
    assign wire_5724 = lut_tile_2_4_chanxy_out[62];
    assign wire_5726 = lut_tile_2_4_chanxy_out[63];
    assign wire_5728 = lut_tile_2_4_chanxy_out[64];
    assign wire_5730 = lut_tile_2_4_chanxy_out[65];
    assign wire_5732 = lut_tile_2_4_chanxy_out[66];
    assign wire_5734 = lut_tile_2_4_chanxy_out[67];
    assign wire_5736 = lut_tile_2_4_chanxy_out[68];
    assign wire_5738 = lut_tile_2_4_chanxy_out[69];
    assign wire_5740 = lut_tile_2_4_chanxy_out[70];
    assign wire_5742 = lut_tile_2_4_chanxy_out[71];
    assign wire_5744 = lut_tile_2_4_chanxy_out[72];
    assign wire_5746 = lut_tile_2_4_chanxy_out[73];
    assign wire_5748 = lut_tile_2_4_chanxy_out[74];
    assign wire_5750 = lut_tile_2_4_chanxy_out[75];
    assign wire_5752 = lut_tile_2_4_chanxy_out[76];
    assign wire_5754 = lut_tile_2_4_chanxy_out[77];
    assign wire_5756 = lut_tile_2_4_chanxy_out[78];
    assign wire_5758 = lut_tile_2_4_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_2_5_chanxy_in = {wire_6036, wire_2918, wire_2908, wire_2898, wire_2888, wire_2211, wire_2205, wire_2196, wire_1901, wire_6028, wire_2878, wire_2868, wire_2858, wire_2848, wire_2211, wire_2205, wire_2196, wire_1901, wire_6020, wire_2998, wire_2988, wire_2978, wire_2968, wire_2211, wire_2205, wire_2196, wire_1901, wire_6012, wire_2958, wire_2948, wire_2938, wire_2928, wire_2211, wire_2205, wire_2196, wire_1901, wire_6004, wire_2916, wire_2906, wire_2896, wire_2886, wire_2211, wire_2202, wire_2196, wire_1897, wire_5996, wire_2876, wire_2866, wire_2856, wire_2846, wire_2211, wire_2202, wire_2196, wire_1897, wire_5988, wire_2996, wire_2986, wire_2976, wire_2966, wire_2211, wire_2202, wire_2196, wire_1897, wire_5980, wire_2956, wire_2946, wire_2936, wire_2926, wire_2211, wire_2202, wire_2196, wire_1897, wire_5972, wire_2914, wire_2904, wire_2894, wire_2884, wire_2208, wire_2202, wire_2193, wire_1897, wire_5964, wire_2874, wire_2864, wire_2854, wire_2844, wire_2208, wire_2202, wire_2193, wire_1897, wire_5956, wire_2994, wire_2984, wire_2974, wire_2964, wire_2208, wire_2202, wire_2193, wire_1897, wire_5948, wire_2954, wire_2944, wire_2934, wire_2924, wire_2208, wire_2202, wire_2193, wire_1897, wire_5940, wire_2912, wire_2902, wire_2892, wire_2882, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_5932, wire_2872, wire_2862, wire_2852, wire_2842, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_5924, wire_2992, wire_2982, wire_2972, wire_2962, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_5916, wire_2952, wire_2942, wire_2932, wire_2922, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_5908, wire_2910, wire_2900, wire_2890, wire_2880, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_5900, wire_2870, wire_2860, wire_2850, wire_2840, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_5892, wire_2990, wire_2980, wire_2970, wire_2960, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_5884, wire_2950, wire_2940, wire_2930, wire_2920, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_6119, wire_3198, wire_3188, wire_3178, wire_3168, wire_2211, wire_2205, wire_2196, wire_1901, wire_6117, wire_3318, wire_3308, wire_3298, wire_3288, wire_2211, wire_2205, wire_2196, wire_1901, wire_6115, wire_3278, wire_3268, wire_3258, wire_3248, wire_2211, wire_2205, wire_2196, wire_1901, wire_6113, wire_3238, wire_3228, wire_3218, wire_3208, wire_2211, wire_2205, wire_2196, wire_1901, wire_6111, wire_3196, wire_3186, wire_3176, wire_3166, wire_2211, wire_2202, wire_2196, wire_1897, wire_6109, wire_3316, wire_3306, wire_3296, wire_3286, wire_2211, wire_2202, wire_2196, wire_1897, wire_6107, wire_3276, wire_3266, wire_3256, wire_3246, wire_2211, wire_2202, wire_2196, wire_1897, wire_6105, wire_3236, wire_3226, wire_3216, wire_3206, wire_2211, wire_2202, wire_2196, wire_1897, wire_6103, wire_3194, wire_3184, wire_3174, wire_3164, wire_2208, wire_2202, wire_2193, wire_1897, wire_6101, wire_3314, wire_3304, wire_3294, wire_3284, wire_2208, wire_2202, wire_2193, wire_1897, wire_6099, wire_3274, wire_3264, wire_3254, wire_3244, wire_2208, wire_2202, wire_2193, wire_1897, wire_6097, wire_3234, wire_3224, wire_3214, wire_3204, wire_2208, wire_2202, wire_2193, wire_1897, wire_6095, wire_3192, wire_3182, wire_3172, wire_3162, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_6093, wire_3312, wire_3302, wire_3292, wire_3282, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_6091, wire_3272, wire_3262, wire_3252, wire_3242, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_6089, wire_3232, wire_3222, wire_3212, wire_3202, wire_2214, wire_2208, wire_2199, wire_2193, wire_1893, wire_6087, wire_3190, wire_3180, wire_3170, wire_3160, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_6085, wire_3310, wire_3300, wire_3290, wire_3280, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_6083, wire_3270, wire_3260, wire_3250, wire_3240, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_6081, wire_3230, wire_3220, wire_3210, wire_3200, wire_2214, wire_2205, wire_2199, wire_1901, wire_1893, wire_6059, wire_6058, wire_5797, wire_5733, wire_5732, wire_5719, wire_5718, wire_5716, wire_5665, wire_5664, wire_3156, wire_1958, wire_1950, wire_6033, wire_6032, wire_5795, wire_5759, wire_5758, wire_5663, wire_5662, wire_5609, wire_5608, wire_5564, wire_3148, wire_1958, wire_1950, wire_6057, wire_6056, wire_5793, wire_5745, wire_5744, wire_5713, wire_5712, wire_5607, wire_5606, wire_5572, wire_3140, wire_1958, wire_1950, wire_6027, wire_6026, wire_5791, wire_5731, wire_5730, wire_5711, wire_5710, wire_5657, wire_5656, wire_5580, wire_3132, wire_1958, wire_1950, wire_5939, wire_5938, wire_5789, wire_5757, wire_5756, wire_5655, wire_5654, wire_5601, wire_5600, wire_5588, wire_3124, wire_1958, wire_1900, wire_6019, wire_6018, wire_5787, wire_5743, wire_5742, wire_5705, wire_5704, wire_5599, wire_5598, wire_5596, wire_3116, wire_1958, wire_1900, wire_6053, wire_6052, wire_5785, wire_5729, wire_5728, wire_5703, wire_5702, wire_5649, wire_5648, wire_5604, wire_3108, wire_1958, wire_1900, wire_6009, wire_6008, wire_5783, wire_5755, wire_5754, wire_5647, wire_5646, wire_5612, wire_5593, wire_5592, wire_3100, wire_1958, wire_1900, wire_6051, wire_6050, wire_5781, wire_5741, wire_5740, wire_5697, wire_5696, wire_5620, wire_5591, wire_5590, wire_3092, wire_1954, wire_1900, wire_6003, wire_6002, wire_5779, wire_5727, wire_5726, wire_5695, wire_5694, wire_5641, wire_5640, wire_5628, wire_3084, wire_1954, wire_1900, wire_5915, wire_5914, wire_1958, wire_5777, wire_5753, wire_5752, wire_5639, wire_5638, wire_5636, wire_5585, wire_5584, wire_3076, wire_1954, wire_1900, wire_5995, wire_5994, wire_1958, wire_5775, wire_5739, wire_5738, wire_5689, wire_5688, wire_5644, wire_5583, wire_5582, wire_3068, wire_1954, wire_1900, wire_6047, wire_6046, wire_1954, wire_5773, wire_5725, wire_5724, wire_5687, wire_5686, wire_5652, wire_5633, wire_5632, wire_3060, wire_1954, wire_1896, wire_5985, wire_5984, wire_1954, wire_5771, wire_5751, wire_5750, wire_5660, wire_5631, wire_5630, wire_5577, wire_5576, wire_3052, wire_1954, wire_1896, wire_6045, wire_6044, wire_1950, wire_5769, wire_5737, wire_5736, wire_5681, wire_5680, wire_5668, wire_5575, wire_5574, wire_3044, wire_1954, wire_1896, wire_5979, wire_5978, wire_1950, wire_5767, wire_5723, wire_5722, wire_5679, wire_5678, wire_5676, wire_5625, wire_5624, wire_3036, wire_1954, wire_1896, wire_5891, wire_5890, wire_1900, wire_5765, wire_5749, wire_5748, wire_5684, wire_5623, wire_5622, wire_5569, wire_5568, wire_3028, wire_1950, wire_1896, wire_5971, wire_5970, wire_1900, wire_5763, wire_5735, wire_5734, wire_5692, wire_5673, wire_5672, wire_5567, wire_5566, wire_3020, wire_1950, wire_1896, wire_6041, wire_6040, wire_1896, wire_5761, wire_5721, wire_5720, wire_5700, wire_5671, wire_5670, wire_5617, wire_5616, wire_3012, wire_1950, wire_1896, wire_5961, wire_5960, wire_1896, wire_5799, wire_5747, wire_5746, wire_5708, wire_5615, wire_5614, wire_5561, wire_5560, wire_3004, wire_1950, wire_1896, wire_6079, wire_6078, wire_6117, wire_6030, wire_6077, wire_6076, wire_6095, wire_5942, wire_5937, wire_5936, wire_6093, wire_5934, wire_6073, wire_6072, wire_6111, wire_6006, wire_6071, wire_6070, wire_6089, wire_5918, wire_5913, wire_5912, wire_1958, wire_6087, wire_5910, wire_1958, wire_6067, wire_6066, wire_1954, wire_6105, wire_5982, wire_1954, wire_6065, wire_6064, wire_1950, wire_6083, wire_5894, wire_1950, wire_5889, wire_5888, wire_1900, wire_6081, wire_5886, wire_1900, wire_6061, wire_6060, wire_1896, wire_6099, wire_5958, wire_1896, wire_6035, wire_6034, wire_5953, wire_5952, wire_5947, wire_5946, wire_6055, wire_6054, wire_6115, wire_6022, wire_6017, wire_6016, wire_6011, wire_6010, wire_5929, wire_5928, wire_5923, wire_5922, wire_6049, wire_6048, wire_6109, wire_5998, wire_1958, wire_5993, wire_5992, wire_1958, wire_5987, wire_5986, wire_1954, wire_5905, wire_5904, wire_1954, wire_5899, wire_5898, wire_1950, wire_6043, wire_6042, wire_1950, wire_6103, wire_5974, wire_1900, wire_5969, wire_5968, wire_1900, wire_5963, wire_5962, wire_1896, wire_5881, wire_5880, wire_1896, wire_6119, wire_6038, wire_5955, wire_5954, wire_6097, wire_5950, wire_5945, wire_5944, wire_6025, wire_6024, wire_6075, wire_6074, wire_6113, wire_6014, wire_5931, wire_5930, wire_6091, wire_5926, wire_5921, wire_5920, wire_6001, wire_6000, wire_1958, wire_6069, wire_6068, wire_1958, wire_6107, wire_5990, wire_1954, wire_5907, wire_5906, wire_1954, wire_6085, wire_5902, wire_1950, wire_5897, wire_5896, wire_1950, wire_5977, wire_5976, wire_1900, wire_6063, wire_6062, wire_1900, wire_6101, wire_5966, wire_1896, wire_5883, wire_5882, wire_1896};
    // CHNAXY TOTAL: 796
    assign wire_3161 = lut_tile_2_5_chanxy_out[0];
    assign wire_3163 = lut_tile_2_5_chanxy_out[1];
    assign wire_3165 = lut_tile_2_5_chanxy_out[2];
    assign wire_3167 = lut_tile_2_5_chanxy_out[3];
    assign wire_3169 = lut_tile_2_5_chanxy_out[4];
    assign wire_3171 = lut_tile_2_5_chanxy_out[5];
    assign wire_3173 = lut_tile_2_5_chanxy_out[6];
    assign wire_3175 = lut_tile_2_5_chanxy_out[7];
    assign wire_3177 = lut_tile_2_5_chanxy_out[8];
    assign wire_3179 = lut_tile_2_5_chanxy_out[9];
    assign wire_3181 = lut_tile_2_5_chanxy_out[10];
    assign wire_3183 = lut_tile_2_5_chanxy_out[11];
    assign wire_3185 = lut_tile_2_5_chanxy_out[12];
    assign wire_3187 = lut_tile_2_5_chanxy_out[13];
    assign wire_3189 = lut_tile_2_5_chanxy_out[14];
    assign wire_3191 = lut_tile_2_5_chanxy_out[15];
    assign wire_3193 = lut_tile_2_5_chanxy_out[16];
    assign wire_3195 = lut_tile_2_5_chanxy_out[17];
    assign wire_3197 = lut_tile_2_5_chanxy_out[18];
    assign wire_3199 = lut_tile_2_5_chanxy_out[19];
    assign wire_3201 = lut_tile_2_5_chanxy_out[20];
    assign wire_3203 = lut_tile_2_5_chanxy_out[21];
    assign wire_3205 = lut_tile_2_5_chanxy_out[22];
    assign wire_3207 = lut_tile_2_5_chanxy_out[23];
    assign wire_3209 = lut_tile_2_5_chanxy_out[24];
    assign wire_3211 = lut_tile_2_5_chanxy_out[25];
    assign wire_3213 = lut_tile_2_5_chanxy_out[26];
    assign wire_3215 = lut_tile_2_5_chanxy_out[27];
    assign wire_3217 = lut_tile_2_5_chanxy_out[28];
    assign wire_3219 = lut_tile_2_5_chanxy_out[29];
    assign wire_3221 = lut_tile_2_5_chanxy_out[30];
    assign wire_3223 = lut_tile_2_5_chanxy_out[31];
    assign wire_3225 = lut_tile_2_5_chanxy_out[32];
    assign wire_3227 = lut_tile_2_5_chanxy_out[33];
    assign wire_3229 = lut_tile_2_5_chanxy_out[34];
    assign wire_3231 = lut_tile_2_5_chanxy_out[35];
    assign wire_3233 = lut_tile_2_5_chanxy_out[36];
    assign wire_3235 = lut_tile_2_5_chanxy_out[37];
    assign wire_3237 = lut_tile_2_5_chanxy_out[38];
    assign wire_3239 = lut_tile_2_5_chanxy_out[39];
    assign wire_3241 = lut_tile_2_5_chanxy_out[40];
    assign wire_3243 = lut_tile_2_5_chanxy_out[41];
    assign wire_3245 = lut_tile_2_5_chanxy_out[42];
    assign wire_3247 = lut_tile_2_5_chanxy_out[43];
    assign wire_3249 = lut_tile_2_5_chanxy_out[44];
    assign wire_3251 = lut_tile_2_5_chanxy_out[45];
    assign wire_3253 = lut_tile_2_5_chanxy_out[46];
    assign wire_3255 = lut_tile_2_5_chanxy_out[47];
    assign wire_3257 = lut_tile_2_5_chanxy_out[48];
    assign wire_3259 = lut_tile_2_5_chanxy_out[49];
    assign wire_3261 = lut_tile_2_5_chanxy_out[50];
    assign wire_3263 = lut_tile_2_5_chanxy_out[51];
    assign wire_3265 = lut_tile_2_5_chanxy_out[52];
    assign wire_3267 = lut_tile_2_5_chanxy_out[53];
    assign wire_3269 = lut_tile_2_5_chanxy_out[54];
    assign wire_3271 = lut_tile_2_5_chanxy_out[55];
    assign wire_3273 = lut_tile_2_5_chanxy_out[56];
    assign wire_3275 = lut_tile_2_5_chanxy_out[57];
    assign wire_3277 = lut_tile_2_5_chanxy_out[58];
    assign wire_3279 = lut_tile_2_5_chanxy_out[59];
    assign wire_3280 = lut_tile_2_5_chanxy_out[60];
    assign wire_3281 = lut_tile_2_5_chanxy_out[61];
    assign wire_3282 = lut_tile_2_5_chanxy_out[62];
    assign wire_3283 = lut_tile_2_5_chanxy_out[63];
    assign wire_3284 = lut_tile_2_5_chanxy_out[64];
    assign wire_3285 = lut_tile_2_5_chanxy_out[65];
    assign wire_3286 = lut_tile_2_5_chanxy_out[66];
    assign wire_3287 = lut_tile_2_5_chanxy_out[67];
    assign wire_3288 = lut_tile_2_5_chanxy_out[68];
    assign wire_3289 = lut_tile_2_5_chanxy_out[69];
    assign wire_3290 = lut_tile_2_5_chanxy_out[70];
    assign wire_3291 = lut_tile_2_5_chanxy_out[71];
    assign wire_3292 = lut_tile_2_5_chanxy_out[72];
    assign wire_3293 = lut_tile_2_5_chanxy_out[73];
    assign wire_3294 = lut_tile_2_5_chanxy_out[74];
    assign wire_3295 = lut_tile_2_5_chanxy_out[75];
    assign wire_3296 = lut_tile_2_5_chanxy_out[76];
    assign wire_3297 = lut_tile_2_5_chanxy_out[77];
    assign wire_3298 = lut_tile_2_5_chanxy_out[78];
    assign wire_3299 = lut_tile_2_5_chanxy_out[79];
    assign wire_3300 = lut_tile_2_5_chanxy_out[80];
    assign wire_3301 = lut_tile_2_5_chanxy_out[81];
    assign wire_3302 = lut_tile_2_5_chanxy_out[82];
    assign wire_3303 = lut_tile_2_5_chanxy_out[83];
    assign wire_3304 = lut_tile_2_5_chanxy_out[84];
    assign wire_3305 = lut_tile_2_5_chanxy_out[85];
    assign wire_3306 = lut_tile_2_5_chanxy_out[86];
    assign wire_3307 = lut_tile_2_5_chanxy_out[87];
    assign wire_3308 = lut_tile_2_5_chanxy_out[88];
    assign wire_3309 = lut_tile_2_5_chanxy_out[89];
    assign wire_3310 = lut_tile_2_5_chanxy_out[90];
    assign wire_3311 = lut_tile_2_5_chanxy_out[91];
    assign wire_3312 = lut_tile_2_5_chanxy_out[92];
    assign wire_3313 = lut_tile_2_5_chanxy_out[93];
    assign wire_3314 = lut_tile_2_5_chanxy_out[94];
    assign wire_3315 = lut_tile_2_5_chanxy_out[95];
    assign wire_3316 = lut_tile_2_5_chanxy_out[96];
    assign wire_3317 = lut_tile_2_5_chanxy_out[97];
    assign wire_3318 = lut_tile_2_5_chanxy_out[98];
    assign wire_3319 = lut_tile_2_5_chanxy_out[99];
    assign wire_5887 = lut_tile_2_5_chanxy_out[100];
    assign wire_5895 = lut_tile_2_5_chanxy_out[101];
    assign wire_5903 = lut_tile_2_5_chanxy_out[102];
    assign wire_5911 = lut_tile_2_5_chanxy_out[103];
    assign wire_5919 = lut_tile_2_5_chanxy_out[104];
    assign wire_5927 = lut_tile_2_5_chanxy_out[105];
    assign wire_5935 = lut_tile_2_5_chanxy_out[106];
    assign wire_5943 = lut_tile_2_5_chanxy_out[107];
    assign wire_5951 = lut_tile_2_5_chanxy_out[108];
    assign wire_5959 = lut_tile_2_5_chanxy_out[109];
    assign wire_5967 = lut_tile_2_5_chanxy_out[110];
    assign wire_5975 = lut_tile_2_5_chanxy_out[111];
    assign wire_5983 = lut_tile_2_5_chanxy_out[112];
    assign wire_5991 = lut_tile_2_5_chanxy_out[113];
    assign wire_5999 = lut_tile_2_5_chanxy_out[114];
    assign wire_6007 = lut_tile_2_5_chanxy_out[115];
    assign wire_6015 = lut_tile_2_5_chanxy_out[116];
    assign wire_6023 = lut_tile_2_5_chanxy_out[117];
    assign wire_6031 = lut_tile_2_5_chanxy_out[118];
    assign wire_6039 = lut_tile_2_5_chanxy_out[119];
    assign wire_6040 = lut_tile_2_5_chanxy_out[120];
    assign wire_6042 = lut_tile_2_5_chanxy_out[121];
    assign wire_6044 = lut_tile_2_5_chanxy_out[122];
    assign wire_6046 = lut_tile_2_5_chanxy_out[123];
    assign wire_6048 = lut_tile_2_5_chanxy_out[124];
    assign wire_6050 = lut_tile_2_5_chanxy_out[125];
    assign wire_6052 = lut_tile_2_5_chanxy_out[126];
    assign wire_6054 = lut_tile_2_5_chanxy_out[127];
    assign wire_6056 = lut_tile_2_5_chanxy_out[128];
    assign wire_6058 = lut_tile_2_5_chanxy_out[129];
    assign wire_6060 = lut_tile_2_5_chanxy_out[130];
    assign wire_6062 = lut_tile_2_5_chanxy_out[131];
    assign wire_6064 = lut_tile_2_5_chanxy_out[132];
    assign wire_6066 = lut_tile_2_5_chanxy_out[133];
    assign wire_6068 = lut_tile_2_5_chanxy_out[134];
    assign wire_6070 = lut_tile_2_5_chanxy_out[135];
    assign wire_6072 = lut_tile_2_5_chanxy_out[136];
    assign wire_6074 = lut_tile_2_5_chanxy_out[137];
    assign wire_6076 = lut_tile_2_5_chanxy_out[138];
    assign wire_6078 = lut_tile_2_5_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_3_1_chanxy_in = {wire_4758, wire_3161, wire_3157, wire_3156, wire_3105, wire_3104, wire_3051, wire_3050, wire_3014, wire_827, wire_453, wire_4750, wire_3199, wire_3155, wire_3154, wire_3101, wire_3100, wire_3049, wire_3048, wire_3022, wire_827, wire_453, wire_4742, wire_3197, wire_3153, wire_3152, wire_3099, wire_3098, wire_3045, wire_3044, wire_3030, wire_827, wire_453, wire_4734, wire_3195, wire_3149, wire_3148, wire_3097, wire_3096, wire_3043, wire_3042, wire_3038, wire_827, wire_453, wire_4726, wire_3193, wire_3147, wire_3146, wire_3093, wire_3092, wire_3046, wire_3041, wire_3040, wire_827, wire_449, wire_4718, wire_3191, wire_3145, wire_3144, wire_3091, wire_3090, wire_3054, wire_3037, wire_3036, wire_827, wire_449, wire_4710, wire_3189, wire_3141, wire_3140, wire_3089, wire_3088, wire_3062, wire_3035, wire_3034, wire_827, wire_449, wire_4702, wire_3187, wire_3139, wire_3138, wire_3085, wire_3084, wire_3070, wire_3033, wire_3032, wire_827, wire_449, wire_4694, wire_3185, wire_3137, wire_3136, wire_3083, wire_3082, wire_3078, wire_3029, wire_3028, wire_823, wire_449, wire_4686, wire_3183, wire_3133, wire_3132, wire_3086, wire_3081, wire_3080, wire_3027, wire_3026, wire_823, wire_449, wire_4678, wire_3181, wire_3131, wire_3130, wire_3094, wire_3077, wire_3076, wire_3025, wire_3024, wire_823, wire_449, wire_4670, wire_3179, wire_3129, wire_3128, wire_3102, wire_3075, wire_3074, wire_3021, wire_3020, wire_823, wire_449, wire_4662, wire_3177, wire_3125, wire_3124, wire_3110, wire_3073, wire_3072, wire_3019, wire_3018, wire_823, wire_445, wire_4654, wire_3175, wire_3123, wire_3122, wire_3118, wire_3069, wire_3068, wire_3017, wire_3016, wire_823, wire_445, wire_4646, wire_3173, wire_3126, wire_3121, wire_3120, wire_3067, wire_3066, wire_3013, wire_3012, wire_823, wire_445, wire_4638, wire_3171, wire_3134, wire_3117, wire_3116, wire_3065, wire_3064, wire_3011, wire_3010, wire_823, wire_445, wire_4630, wire_3169, wire_3142, wire_3115, wire_3114, wire_3061, wire_3060, wire_3009, wire_3008, wire_453, wire_445, wire_4622, wire_3167, wire_3150, wire_3113, wire_3112, wire_3059, wire_3058, wire_3005, wire_3004, wire_453, wire_445, wire_4614, wire_3165, wire_3158, wire_3109, wire_3108, wire_3057, wire_3056, wire_3003, wire_3002, wire_453, wire_445, wire_4606, wire_3163, wire_3107, wire_3106, wire_3053, wire_3052, wire_3006, wire_3001, wire_3000, wire_453, wire_445, wire_4879, wire_3519, wire_3479, wire_3478, wire_3427, wire_3426, wire_3373, wire_3372, wire_3320, wire_827, wire_453, wire_4877, wire_3481, wire_3477, wire_3476, wire_3472, wire_3423, wire_3422, wire_3371, wire_3370, wire_827, wire_453, wire_4875, wire_3483, wire_3475, wire_3474, wire_3464, wire_3421, wire_3420, wire_3367, wire_3366, wire_827, wire_453, wire_4873, wire_3485, wire_3471, wire_3470, wire_3456, wire_3419, wire_3418, wire_3365, wire_3364, wire_827, wire_453, wire_4871, wire_3487, wire_3469, wire_3468, wire_3448, wire_3415, wire_3414, wire_3363, wire_3362, wire_827, wire_449, wire_4869, wire_3489, wire_3467, wire_3466, wire_3440, wire_3413, wire_3412, wire_3359, wire_3358, wire_827, wire_449, wire_4867, wire_3491, wire_3463, wire_3462, wire_3432, wire_3411, wire_3410, wire_3357, wire_3356, wire_827, wire_449, wire_4865, wire_3493, wire_3461, wire_3460, wire_3424, wire_3407, wire_3406, wire_3355, wire_3354, wire_827, wire_449, wire_4863, wire_3495, wire_3459, wire_3458, wire_3416, wire_3405, wire_3404, wire_3351, wire_3350, wire_823, wire_449, wire_4861, wire_3497, wire_3455, wire_3454, wire_3408, wire_3403, wire_3402, wire_3349, wire_3348, wire_823, wire_449, wire_4859, wire_3499, wire_3453, wire_3452, wire_3400, wire_3399, wire_3398, wire_3347, wire_3346, wire_823, wire_449, wire_4857, wire_3501, wire_3451, wire_3450, wire_3397, wire_3396, wire_3392, wire_3343, wire_3342, wire_823, wire_449, wire_4855, wire_3503, wire_3447, wire_3446, wire_3395, wire_3394, wire_3384, wire_3341, wire_3340, wire_823, wire_445, wire_4853, wire_3505, wire_3445, wire_3444, wire_3391, wire_3390, wire_3376, wire_3339, wire_3338, wire_823, wire_445, wire_4851, wire_3507, wire_3443, wire_3442, wire_3389, wire_3388, wire_3368, wire_3335, wire_3334, wire_823, wire_445, wire_4849, wire_3509, wire_3439, wire_3438, wire_3387, wire_3386, wire_3360, wire_3333, wire_3332, wire_823, wire_445, wire_4847, wire_3511, wire_3437, wire_3436, wire_3383, wire_3382, wire_3352, wire_3331, wire_3330, wire_453, wire_445, wire_4845, wire_3513, wire_3435, wire_3434, wire_3381, wire_3380, wire_3344, wire_3327, wire_3326, wire_453, wire_445, wire_4843, wire_3515, wire_3431, wire_3430, wire_3379, wire_3378, wire_3336, wire_3325, wire_3324, wire_453, wire_445, wire_4841, wire_3517, wire_3429, wire_3428, wire_3375, wire_3374, wire_3328, wire_3323, wire_3322, wire_453, wire_445, wire_4559, wire_4438, wire_4519, wire_4518, wire_4459, wire_4458, wire_4843, wire_4839, wire_4838, wire_4773, wire_4772, wire_4744, wire_4707, wire_4706, wire_3519, wire_510, wire_502, wire_4479, wire_4478, wire_4433, wire_4432, wire_4353, wire_4352, wire_4557, wire_4430, wire_4845, wire_4825, wire_4824, wire_4799, wire_4798, wire_4736, wire_4651, wire_4650, wire_3517, wire_510, wire_502, wire_4517, wire_4516, wire_4477, wire_4476, wire_4537, wire_4350, wire_4497, wire_4496, wire_4847, wire_4811, wire_4810, wire_4785, wire_4784, wire_4755, wire_4754, wire_4728, wire_3515, wire_510, wire_502, wire_4425, wire_4424, wire_4457, wire_4456, wire_4345, wire_4344, wire_4555, wire_4422, wire_4849, wire_4837, wire_4836, wire_4771, wire_4770, wire_4720, wire_4699, wire_4698, wire_3513, wire_510, wire_502, wire_4535, wire_4342, wire_4495, wire_4494, wire_4515, wire_4514, wire_4455, wire_4454, wire_4851, wire_4823, wire_4822, wire_4797, wire_4796, wire_4712, wire_4643, wire_4642, wire_3511, wire_510, wire_452, wire_4337, wire_4336, wire_4533, wire_4334, wire_4475, wire_4474, wire_4417, wire_4416, wire_4853, wire_4809, wire_4808, wire_4783, wire_4782, wire_4747, wire_4746, wire_4704, wire_3509, wire_510, wire_452, wire_4493, wire_4492, wire_4553, wire_4414, wire_4513, wire_4512, wire_4453, wire_4452, wire_4855, wire_4835, wire_4834, wire_4769, wire_4768, wire_4696, wire_4691, wire_4690, wire_3507, wire_510, wire_452, wire_4473, wire_4472, wire_4409, wire_4408, wire_4329, wire_4328, wire_4551, wire_4406, wire_4857, wire_4821, wire_4820, wire_4795, wire_4794, wire_4688, wire_4635, wire_4634, wire_3505, wire_510, wire_452, wire_4511, wire_4510, wire_4471, wire_4470, wire_4531, wire_4326, wire_4491, wire_4490, wire_4859, wire_4807, wire_4806, wire_4781, wire_4780, wire_4739, wire_4738, wire_4680, wire_3503, wire_506, wire_452, wire_4401, wire_4400, wire_4451, wire_4450, wire_4321, wire_4320, wire_4549, wire_4398, wire_4861, wire_4833, wire_4832, wire_4767, wire_4766, wire_4683, wire_4682, wire_4672, wire_3501, wire_506, wire_452, wire_4529, wire_4318, wire_4489, wire_4488, wire_510, wire_4509, wire_4508, wire_510, wire_4449, wire_4448, wire_510, wire_4863, wire_4819, wire_4818, wire_4793, wire_4792, wire_4664, wire_4627, wire_4626, wire_3499, wire_506, wire_452, wire_4313, wire_4312, wire_510, wire_4527, wire_4310, wire_510, wire_4469, wire_4468, wire_510, wire_4393, wire_4392, wire_510, wire_4865, wire_4805, wire_4804, wire_4779, wire_4778, wire_4731, wire_4730, wire_4656, wire_3497, wire_506, wire_452, wire_4487, wire_4486, wire_510, wire_4547, wire_4390, wire_506, wire_4507, wire_4506, wire_506, wire_4447, wire_4446, wire_506, wire_4867, wire_4831, wire_4830, wire_4765, wire_4764, wire_4675, wire_4674, wire_4648, wire_3495, wire_506, wire_448, wire_4467, wire_4466, wire_506, wire_4385, wire_4384, wire_506, wire_4305, wire_4304, wire_506, wire_4545, wire_4382, wire_506, wire_4869, wire_4817, wire_4816, wire_4791, wire_4790, wire_4640, wire_4619, wire_4618, wire_3493, wire_506, wire_448, wire_4505, wire_4504, wire_506, wire_4465, wire_4464, wire_502, wire_4525, wire_4302, wire_502, wire_4485, wire_4484, wire_502, wire_4871, wire_4803, wire_4802, wire_4777, wire_4776, wire_4723, wire_4722, wire_4632, wire_3491, wire_506, wire_448, wire_4377, wire_4376, wire_502, wire_4445, wire_4444, wire_502, wire_4297, wire_4296, wire_502, wire_4543, wire_4374, wire_502, wire_4873, wire_4829, wire_4828, wire_4763, wire_4762, wire_4667, wire_4666, wire_4624, wire_3489, wire_506, wire_448, wire_4523, wire_4294, wire_502, wire_4483, wire_4482, wire_452, wire_4503, wire_4502, wire_452, wire_4443, wire_4442, wire_452, wire_4875, wire_4815, wire_4814, wire_4789, wire_4788, wire_4616, wire_4611, wire_4610, wire_3487, wire_502, wire_448, wire_4289, wire_4288, wire_452, wire_4521, wire_4286, wire_452, wire_4463, wire_4462, wire_452, wire_4369, wire_4368, wire_452, wire_4877, wire_4801, wire_4800, wire_4775, wire_4774, wire_4715, wire_4714, wire_4608, wire_3485, wire_502, wire_448, wire_4481, wire_4480, wire_452, wire_4541, wire_4366, wire_448, wire_4501, wire_4500, wire_448, wire_4441, wire_4440, wire_448, wire_4879, wire_4827, wire_4826, wire_4761, wire_4760, wire_4659, wire_4658, wire_4600, wire_3483, wire_502, wire_448, wire_4461, wire_4460, wire_448, wire_4361, wire_4360, wire_448, wire_4281, wire_4280, wire_448, wire_4539, wire_4358, wire_448, wire_4841, wire_4813, wire_4812, wire_4787, wire_4786, wire_4752, wire_4603, wire_4602, wire_3481, wire_502, wire_448, wire_4499, wire_4498, wire_448};
    // CHNAXY TOTAL: 860
    assign wire_3320 = lut_tile_3_1_chanxy_out[0];
    assign wire_3321 = lut_tile_3_1_chanxy_out[1];
    assign wire_3322 = lut_tile_3_1_chanxy_out[2];
    assign wire_3324 = lut_tile_3_1_chanxy_out[3];
    assign wire_3326 = lut_tile_3_1_chanxy_out[4];
    assign wire_3328 = lut_tile_3_1_chanxy_out[5];
    assign wire_3329 = lut_tile_3_1_chanxy_out[6];
    assign wire_3330 = lut_tile_3_1_chanxy_out[7];
    assign wire_3332 = lut_tile_3_1_chanxy_out[8];
    assign wire_3334 = lut_tile_3_1_chanxy_out[9];
    assign wire_3336 = lut_tile_3_1_chanxy_out[10];
    assign wire_3337 = lut_tile_3_1_chanxy_out[11];
    assign wire_3338 = lut_tile_3_1_chanxy_out[12];
    assign wire_3340 = lut_tile_3_1_chanxy_out[13];
    assign wire_3342 = lut_tile_3_1_chanxy_out[14];
    assign wire_3344 = lut_tile_3_1_chanxy_out[15];
    assign wire_3345 = lut_tile_3_1_chanxy_out[16];
    assign wire_3346 = lut_tile_3_1_chanxy_out[17];
    assign wire_3348 = lut_tile_3_1_chanxy_out[18];
    assign wire_3350 = lut_tile_3_1_chanxy_out[19];
    assign wire_3352 = lut_tile_3_1_chanxy_out[20];
    assign wire_3353 = lut_tile_3_1_chanxy_out[21];
    assign wire_3354 = lut_tile_3_1_chanxy_out[22];
    assign wire_3356 = lut_tile_3_1_chanxy_out[23];
    assign wire_3358 = lut_tile_3_1_chanxy_out[24];
    assign wire_3360 = lut_tile_3_1_chanxy_out[25];
    assign wire_3361 = lut_tile_3_1_chanxy_out[26];
    assign wire_3362 = lut_tile_3_1_chanxy_out[27];
    assign wire_3364 = lut_tile_3_1_chanxy_out[28];
    assign wire_3366 = lut_tile_3_1_chanxy_out[29];
    assign wire_3368 = lut_tile_3_1_chanxy_out[30];
    assign wire_3369 = lut_tile_3_1_chanxy_out[31];
    assign wire_3370 = lut_tile_3_1_chanxy_out[32];
    assign wire_3372 = lut_tile_3_1_chanxy_out[33];
    assign wire_3374 = lut_tile_3_1_chanxy_out[34];
    assign wire_3376 = lut_tile_3_1_chanxy_out[35];
    assign wire_3377 = lut_tile_3_1_chanxy_out[36];
    assign wire_3378 = lut_tile_3_1_chanxy_out[37];
    assign wire_3380 = lut_tile_3_1_chanxy_out[38];
    assign wire_3382 = lut_tile_3_1_chanxy_out[39];
    assign wire_3384 = lut_tile_3_1_chanxy_out[40];
    assign wire_3385 = lut_tile_3_1_chanxy_out[41];
    assign wire_3386 = lut_tile_3_1_chanxy_out[42];
    assign wire_3388 = lut_tile_3_1_chanxy_out[43];
    assign wire_3390 = lut_tile_3_1_chanxy_out[44];
    assign wire_3392 = lut_tile_3_1_chanxy_out[45];
    assign wire_3393 = lut_tile_3_1_chanxy_out[46];
    assign wire_3394 = lut_tile_3_1_chanxy_out[47];
    assign wire_3396 = lut_tile_3_1_chanxy_out[48];
    assign wire_3398 = lut_tile_3_1_chanxy_out[49];
    assign wire_3400 = lut_tile_3_1_chanxy_out[50];
    assign wire_3401 = lut_tile_3_1_chanxy_out[51];
    assign wire_3402 = lut_tile_3_1_chanxy_out[52];
    assign wire_3404 = lut_tile_3_1_chanxy_out[53];
    assign wire_3406 = lut_tile_3_1_chanxy_out[54];
    assign wire_3408 = lut_tile_3_1_chanxy_out[55];
    assign wire_3409 = lut_tile_3_1_chanxy_out[56];
    assign wire_3410 = lut_tile_3_1_chanxy_out[57];
    assign wire_3412 = lut_tile_3_1_chanxy_out[58];
    assign wire_3414 = lut_tile_3_1_chanxy_out[59];
    assign wire_3416 = lut_tile_3_1_chanxy_out[60];
    assign wire_3417 = lut_tile_3_1_chanxy_out[61];
    assign wire_3418 = lut_tile_3_1_chanxy_out[62];
    assign wire_3420 = lut_tile_3_1_chanxy_out[63];
    assign wire_3422 = lut_tile_3_1_chanxy_out[64];
    assign wire_3424 = lut_tile_3_1_chanxy_out[65];
    assign wire_3425 = lut_tile_3_1_chanxy_out[66];
    assign wire_3426 = lut_tile_3_1_chanxy_out[67];
    assign wire_3428 = lut_tile_3_1_chanxy_out[68];
    assign wire_3430 = lut_tile_3_1_chanxy_out[69];
    assign wire_3432 = lut_tile_3_1_chanxy_out[70];
    assign wire_3433 = lut_tile_3_1_chanxy_out[71];
    assign wire_3434 = lut_tile_3_1_chanxy_out[72];
    assign wire_3436 = lut_tile_3_1_chanxy_out[73];
    assign wire_3438 = lut_tile_3_1_chanxy_out[74];
    assign wire_3440 = lut_tile_3_1_chanxy_out[75];
    assign wire_3441 = lut_tile_3_1_chanxy_out[76];
    assign wire_3442 = lut_tile_3_1_chanxy_out[77];
    assign wire_3444 = lut_tile_3_1_chanxy_out[78];
    assign wire_3446 = lut_tile_3_1_chanxy_out[79];
    assign wire_3448 = lut_tile_3_1_chanxy_out[80];
    assign wire_3449 = lut_tile_3_1_chanxy_out[81];
    assign wire_3450 = lut_tile_3_1_chanxy_out[82];
    assign wire_3452 = lut_tile_3_1_chanxy_out[83];
    assign wire_3454 = lut_tile_3_1_chanxy_out[84];
    assign wire_3456 = lut_tile_3_1_chanxy_out[85];
    assign wire_3457 = lut_tile_3_1_chanxy_out[86];
    assign wire_3458 = lut_tile_3_1_chanxy_out[87];
    assign wire_3460 = lut_tile_3_1_chanxy_out[88];
    assign wire_3462 = lut_tile_3_1_chanxy_out[89];
    assign wire_3464 = lut_tile_3_1_chanxy_out[90];
    assign wire_3465 = lut_tile_3_1_chanxy_out[91];
    assign wire_3466 = lut_tile_3_1_chanxy_out[92];
    assign wire_3468 = lut_tile_3_1_chanxy_out[93];
    assign wire_3470 = lut_tile_3_1_chanxy_out[94];
    assign wire_3472 = lut_tile_3_1_chanxy_out[95];
    assign wire_3473 = lut_tile_3_1_chanxy_out[96];
    assign wire_3474 = lut_tile_3_1_chanxy_out[97];
    assign wire_3476 = lut_tile_3_1_chanxy_out[98];
    assign wire_3478 = lut_tile_3_1_chanxy_out[99];
    assign wire_4601 = lut_tile_3_1_chanxy_out[100];
    assign wire_4609 = lut_tile_3_1_chanxy_out[101];
    assign wire_4617 = lut_tile_3_1_chanxy_out[102];
    assign wire_4625 = lut_tile_3_1_chanxy_out[103];
    assign wire_4633 = lut_tile_3_1_chanxy_out[104];
    assign wire_4641 = lut_tile_3_1_chanxy_out[105];
    assign wire_4649 = lut_tile_3_1_chanxy_out[106];
    assign wire_4657 = lut_tile_3_1_chanxy_out[107];
    assign wire_4665 = lut_tile_3_1_chanxy_out[108];
    assign wire_4673 = lut_tile_3_1_chanxy_out[109];
    assign wire_4681 = lut_tile_3_1_chanxy_out[110];
    assign wire_4689 = lut_tile_3_1_chanxy_out[111];
    assign wire_4697 = lut_tile_3_1_chanxy_out[112];
    assign wire_4705 = lut_tile_3_1_chanxy_out[113];
    assign wire_4713 = lut_tile_3_1_chanxy_out[114];
    assign wire_4721 = lut_tile_3_1_chanxy_out[115];
    assign wire_4729 = lut_tile_3_1_chanxy_out[116];
    assign wire_4737 = lut_tile_3_1_chanxy_out[117];
    assign wire_4745 = lut_tile_3_1_chanxy_out[118];
    assign wire_4753 = lut_tile_3_1_chanxy_out[119];
    assign wire_4800 = lut_tile_3_1_chanxy_out[120];
    assign wire_4802 = lut_tile_3_1_chanxy_out[121];
    assign wire_4804 = lut_tile_3_1_chanxy_out[122];
    assign wire_4806 = lut_tile_3_1_chanxy_out[123];
    assign wire_4808 = lut_tile_3_1_chanxy_out[124];
    assign wire_4810 = lut_tile_3_1_chanxy_out[125];
    assign wire_4812 = lut_tile_3_1_chanxy_out[126];
    assign wire_4814 = lut_tile_3_1_chanxy_out[127];
    assign wire_4816 = lut_tile_3_1_chanxy_out[128];
    assign wire_4818 = lut_tile_3_1_chanxy_out[129];
    assign wire_4820 = lut_tile_3_1_chanxy_out[130];
    assign wire_4822 = lut_tile_3_1_chanxy_out[131];
    assign wire_4824 = lut_tile_3_1_chanxy_out[132];
    assign wire_4826 = lut_tile_3_1_chanxy_out[133];
    assign wire_4828 = lut_tile_3_1_chanxy_out[134];
    assign wire_4830 = lut_tile_3_1_chanxy_out[135];
    assign wire_4832 = lut_tile_3_1_chanxy_out[136];
    assign wire_4834 = lut_tile_3_1_chanxy_out[137];
    assign wire_4836 = lut_tile_3_1_chanxy_out[138];
    assign wire_4838 = lut_tile_3_1_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_3_2_chanxy_in = {wire_5072, wire_3201, wire_3199, wire_3198, wire_3107, wire_3106, wire_3053, wire_3052, wire_3008, wire_1203, wire_829, wire_5064, wire_3239, wire_3185, wire_3184, wire_3157, wire_3156, wire_3051, wire_3050, wire_3016, wire_1203, wire_829, wire_5056, wire_3237, wire_3171, wire_3170, wire_3155, wire_3154, wire_3101, wire_3100, wire_3024, wire_1203, wire_829, wire_5048, wire_3235, wire_3197, wire_3196, wire_3099, wire_3098, wire_3045, wire_3044, wire_3032, wire_1203, wire_829, wire_5040, wire_3233, wire_3183, wire_3182, wire_3149, wire_3148, wire_3043, wire_3042, wire_3040, wire_1203, wire_825, wire_5032, wire_3231, wire_3169, wire_3168, wire_3147, wire_3146, wire_3093, wire_3092, wire_3048, wire_1203, wire_825, wire_5024, wire_3229, wire_3195, wire_3194, wire_3091, wire_3090, wire_3056, wire_3037, wire_3036, wire_1203, wire_825, wire_5016, wire_3227, wire_3181, wire_3180, wire_3141, wire_3140, wire_3064, wire_3035, wire_3034, wire_1203, wire_825, wire_5008, wire_3225, wire_3167, wire_3166, wire_3139, wire_3138, wire_3085, wire_3084, wire_3072, wire_1199, wire_825, wire_5000, wire_3223, wire_3193, wire_3192, wire_3083, wire_3082, wire_3080, wire_3029, wire_3028, wire_1199, wire_825, wire_4992, wire_3221, wire_3179, wire_3178, wire_3133, wire_3132, wire_3088, wire_3027, wire_3026, wire_1199, wire_825, wire_4984, wire_3219, wire_3165, wire_3164, wire_3131, wire_3130, wire_3096, wire_3077, wire_3076, wire_1199, wire_825, wire_4976, wire_3217, wire_3191, wire_3190, wire_3104, wire_3075, wire_3074, wire_3021, wire_3020, wire_1199, wire_821, wire_4968, wire_3215, wire_3177, wire_3176, wire_3125, wire_3124, wire_3112, wire_3019, wire_3018, wire_1199, wire_821, wire_4960, wire_3213, wire_3163, wire_3162, wire_3123, wire_3122, wire_3120, wire_3069, wire_3068, wire_1199, wire_821, wire_4952, wire_3211, wire_3189, wire_3188, wire_3128, wire_3067, wire_3066, wire_3013, wire_3012, wire_1199, wire_821, wire_4944, wire_3209, wire_3175, wire_3174, wire_3136, wire_3117, wire_3116, wire_3011, wire_3010, wire_829, wire_821, wire_4936, wire_3207, wire_3161, wire_3160, wire_3144, wire_3115, wire_3114, wire_3061, wire_3060, wire_829, wire_821, wire_4928, wire_3205, wire_3187, wire_3186, wire_3152, wire_3059, wire_3058, wire_3005, wire_3004, wire_829, wire_821, wire_4920, wire_3203, wire_3173, wire_3172, wire_3109, wire_3108, wire_3003, wire_3002, wire_3000, wire_829, wire_821, wire_5199, wire_3559, wire_3507, wire_3506, wire_3479, wire_3478, wire_3373, wire_3372, wire_3322, wire_1203, wire_829, wire_5197, wire_3521, wire_3493, wire_3492, wire_3477, wire_3476, wire_3474, wire_3423, wire_3422, wire_1203, wire_829, wire_5195, wire_3523, wire_3519, wire_3518, wire_3466, wire_3421, wire_3420, wire_3367, wire_3366, wire_1203, wire_829, wire_5193, wire_3525, wire_3505, wire_3504, wire_3471, wire_3470, wire_3458, wire_3365, wire_3364, wire_1203, wire_829, wire_5191, wire_3527, wire_3491, wire_3490, wire_3469, wire_3468, wire_3450, wire_3415, wire_3414, wire_1203, wire_825, wire_5189, wire_3529, wire_3517, wire_3516, wire_3442, wire_3413, wire_3412, wire_3359, wire_3358, wire_1203, wire_825, wire_5187, wire_3531, wire_3503, wire_3502, wire_3463, wire_3462, wire_3434, wire_3357, wire_3356, wire_1203, wire_825, wire_5185, wire_3533, wire_3489, wire_3488, wire_3461, wire_3460, wire_3426, wire_3407, wire_3406, wire_1203, wire_825, wire_5183, wire_3535, wire_3515, wire_3514, wire_3418, wire_3405, wire_3404, wire_3351, wire_3350, wire_1199, wire_825, wire_5181, wire_3537, wire_3501, wire_3500, wire_3455, wire_3454, wire_3410, wire_3349, wire_3348, wire_1199, wire_825, wire_5179, wire_3539, wire_3487, wire_3486, wire_3453, wire_3452, wire_3402, wire_3399, wire_3398, wire_1199, wire_825, wire_5177, wire_3541, wire_3513, wire_3512, wire_3397, wire_3396, wire_3394, wire_3343, wire_3342, wire_1199, wire_825, wire_5175, wire_3543, wire_3499, wire_3498, wire_3447, wire_3446, wire_3386, wire_3341, wire_3340, wire_1199, wire_821, wire_5173, wire_3545, wire_3485, wire_3484, wire_3445, wire_3444, wire_3391, wire_3390, wire_3378, wire_1199, wire_821, wire_5171, wire_3547, wire_3511, wire_3510, wire_3389, wire_3388, wire_3370, wire_3335, wire_3334, wire_1199, wire_821, wire_5169, wire_3549, wire_3497, wire_3496, wire_3439, wire_3438, wire_3362, wire_3333, wire_3332, wire_1199, wire_821, wire_5167, wire_3551, wire_3483, wire_3482, wire_3437, wire_3436, wire_3383, wire_3382, wire_3354, wire_829, wire_821, wire_5165, wire_3553, wire_3509, wire_3508, wire_3381, wire_3380, wire_3346, wire_3327, wire_3326, wire_829, wire_821, wire_5163, wire_3555, wire_3495, wire_3494, wire_3431, wire_3430, wire_3338, wire_3325, wire_3324, wire_829, wire_821, wire_5161, wire_3557, wire_3481, wire_3480, wire_3429, wire_3428, wire_3375, wire_3374, wire_3330, wire_829, wire_821, wire_4877, wire_4839, wire_4838, wire_4773, wire_4772, wire_4752, wire_4707, wire_4706, wire_3472, wire_886, wire_878, wire_4875, wire_4825, wire_4824, wire_4799, wire_4798, wire_4651, wire_4650, wire_4600, wire_3464, wire_886, wire_878, wire_4873, wire_4811, wire_4810, wire_4785, wire_4784, wire_4755, wire_4754, wire_4608, wire_3456, wire_886, wire_878, wire_4871, wire_4837, wire_4836, wire_4771, wire_4770, wire_4699, wire_4698, wire_4616, wire_3448, wire_886, wire_878, wire_4869, wire_4823, wire_4822, wire_4797, wire_4796, wire_4643, wire_4642, wire_4624, wire_3440, wire_886, wire_828, wire_4867, wire_4809, wire_4808, wire_4783, wire_4782, wire_4747, wire_4746, wire_4632, wire_3432, wire_886, wire_828, wire_4865, wire_4835, wire_4834, wire_4769, wire_4768, wire_4691, wire_4690, wire_4640, wire_3424, wire_886, wire_828, wire_4863, wire_4821, wire_4820, wire_4795, wire_4794, wire_4648, wire_4635, wire_4634, wire_3416, wire_886, wire_828, wire_4861, wire_4807, wire_4806, wire_4781, wire_4780, wire_4739, wire_4738, wire_4656, wire_3408, wire_882, wire_828, wire_4859, wire_4833, wire_4832, wire_4767, wire_4766, wire_4683, wire_4682, wire_4664, wire_3400, wire_882, wire_828, wire_4857, wire_4819, wire_4818, wire_4793, wire_4792, wire_4672, wire_4627, wire_4626, wire_3392, wire_882, wire_828, wire_4855, wire_4805, wire_4804, wire_4779, wire_4778, wire_4731, wire_4730, wire_4680, wire_3384, wire_882, wire_828, wire_4853, wire_4831, wire_4830, wire_4765, wire_4764, wire_4688, wire_4675, wire_4674, wire_3376, wire_882, wire_824, wire_4851, wire_4817, wire_4816, wire_4791, wire_4790, wire_4696, wire_4619, wire_4618, wire_3368, wire_882, wire_824, wire_4849, wire_4803, wire_4802, wire_4777, wire_4776, wire_4723, wire_4722, wire_4704, wire_3360, wire_882, wire_824, wire_4847, wire_4829, wire_4828, wire_4763, wire_4762, wire_4712, wire_4667, wire_4666, wire_3352, wire_882, wire_824, wire_4845, wire_4815, wire_4814, wire_4789, wire_4788, wire_4720, wire_4611, wire_4610, wire_3344, wire_878, wire_824, wire_4843, wire_4801, wire_4800, wire_4775, wire_4774, wire_4728, wire_4715, wire_4714, wire_3336, wire_878, wire_824, wire_4841, wire_4827, wire_4826, wire_4761, wire_4760, wire_4736, wire_4659, wire_4658, wire_3328, wire_878, wire_824, wire_4879, wire_4813, wire_4812, wire_4787, wire_4786, wire_4744, wire_4603, wire_4602, wire_3320, wire_878, wire_824, wire_5163, wire_5147, wire_5146, wire_5119, wire_5118, wire_5066, wire_4973, wire_4972, wire_3559, wire_886, wire_878, wire_5165, wire_5133, wire_5132, wire_5105, wire_5104, wire_5077, wire_5076, wire_5058, wire_3557, wire_886, wire_878, wire_5167, wire_5159, wire_5158, wire_5091, wire_5090, wire_5050, wire_5021, wire_5020, wire_3555, wire_886, wire_878, wire_5169, wire_5145, wire_5144, wire_5117, wire_5116, wire_5042, wire_4965, wire_4964, wire_3553, wire_886, wire_878, wire_5171, wire_5131, wire_5130, wire_5103, wire_5102, wire_5069, wire_5068, wire_5034, wire_3551, wire_886, wire_828, wire_5173, wire_5157, wire_5156, wire_5089, wire_5088, wire_5026, wire_5013, wire_5012, wire_3549, wire_886, wire_828, wire_5175, wire_5143, wire_5142, wire_5115, wire_5114, wire_5018, wire_4957, wire_4956, wire_3547, wire_886, wire_828, wire_5177, wire_5129, wire_5128, wire_5101, wire_5100, wire_5061, wire_5060, wire_5010, wire_3545, wire_886, wire_828, wire_5179, wire_5155, wire_5154, wire_5087, wire_5086, wire_5005, wire_5004, wire_5002, wire_3543, wire_882, wire_828, wire_5181, wire_5141, wire_5140, wire_5113, wire_5112, wire_4994, wire_4949, wire_4948, wire_3541, wire_882, wire_828, wire_5183, wire_5127, wire_5126, wire_5099, wire_5098, wire_5053, wire_5052, wire_4986, wire_3539, wire_882, wire_828, wire_5185, wire_5153, wire_5152, wire_5085, wire_5084, wire_4997, wire_4996, wire_4978, wire_3537, wire_882, wire_828, wire_5187, wire_5139, wire_5138, wire_5111, wire_5110, wire_4970, wire_4941, wire_4940, wire_3535, wire_882, wire_824, wire_5189, wire_5125, wire_5124, wire_5097, wire_5096, wire_5045, wire_5044, wire_4962, wire_3533, wire_882, wire_824, wire_5191, wire_5151, wire_5150, wire_5083, wire_5082, wire_4989, wire_4988, wire_4954, wire_3531, wire_882, wire_824, wire_5193, wire_5137, wire_5136, wire_5109, wire_5108, wire_4946, wire_4933, wire_4932, wire_3529, wire_882, wire_824, wire_5195, wire_5123, wire_5122, wire_5095, wire_5094, wire_5037, wire_5036, wire_4938, wire_3527, wire_878, wire_824, wire_5197, wire_5149, wire_5148, wire_5081, wire_5080, wire_4981, wire_4980, wire_4930, wire_3525, wire_878, wire_824, wire_5199, wire_5135, wire_5134, wire_5107, wire_5106, wire_4925, wire_4924, wire_4922, wire_3523, wire_878, wire_824, wire_5161, wire_5121, wire_5120, wire_5093, wire_5092, wire_5074, wire_5029, wire_5028, wire_3521, wire_878, wire_824};
    // CHNAXY TOTAL: 880
    assign wire_3323 = lut_tile_3_2_chanxy_out[0];
    assign wire_3331 = lut_tile_3_2_chanxy_out[1];
    assign wire_3339 = lut_tile_3_2_chanxy_out[2];
    assign wire_3347 = lut_tile_3_2_chanxy_out[3];
    assign wire_3355 = lut_tile_3_2_chanxy_out[4];
    assign wire_3363 = lut_tile_3_2_chanxy_out[5];
    assign wire_3371 = lut_tile_3_2_chanxy_out[6];
    assign wire_3379 = lut_tile_3_2_chanxy_out[7];
    assign wire_3387 = lut_tile_3_2_chanxy_out[8];
    assign wire_3395 = lut_tile_3_2_chanxy_out[9];
    assign wire_3403 = lut_tile_3_2_chanxy_out[10];
    assign wire_3411 = lut_tile_3_2_chanxy_out[11];
    assign wire_3419 = lut_tile_3_2_chanxy_out[12];
    assign wire_3427 = lut_tile_3_2_chanxy_out[13];
    assign wire_3435 = lut_tile_3_2_chanxy_out[14];
    assign wire_3443 = lut_tile_3_2_chanxy_out[15];
    assign wire_3451 = lut_tile_3_2_chanxy_out[16];
    assign wire_3459 = lut_tile_3_2_chanxy_out[17];
    assign wire_3467 = lut_tile_3_2_chanxy_out[18];
    assign wire_3475 = lut_tile_3_2_chanxy_out[19];
    assign wire_3480 = lut_tile_3_2_chanxy_out[20];
    assign wire_3482 = lut_tile_3_2_chanxy_out[21];
    assign wire_3484 = lut_tile_3_2_chanxy_out[22];
    assign wire_3486 = lut_tile_3_2_chanxy_out[23];
    assign wire_3488 = lut_tile_3_2_chanxy_out[24];
    assign wire_3490 = lut_tile_3_2_chanxy_out[25];
    assign wire_3492 = lut_tile_3_2_chanxy_out[26];
    assign wire_3494 = lut_tile_3_2_chanxy_out[27];
    assign wire_3496 = lut_tile_3_2_chanxy_out[28];
    assign wire_3498 = lut_tile_3_2_chanxy_out[29];
    assign wire_3500 = lut_tile_3_2_chanxy_out[30];
    assign wire_3502 = lut_tile_3_2_chanxy_out[31];
    assign wire_3504 = lut_tile_3_2_chanxy_out[32];
    assign wire_3506 = lut_tile_3_2_chanxy_out[33];
    assign wire_3508 = lut_tile_3_2_chanxy_out[34];
    assign wire_3510 = lut_tile_3_2_chanxy_out[35];
    assign wire_3512 = lut_tile_3_2_chanxy_out[36];
    assign wire_3514 = lut_tile_3_2_chanxy_out[37];
    assign wire_3516 = lut_tile_3_2_chanxy_out[38];
    assign wire_3518 = lut_tile_3_2_chanxy_out[39];
    assign wire_4923 = lut_tile_3_2_chanxy_out[40];
    assign wire_4931 = lut_tile_3_2_chanxy_out[41];
    assign wire_4939 = lut_tile_3_2_chanxy_out[42];
    assign wire_4947 = lut_tile_3_2_chanxy_out[43];
    assign wire_4955 = lut_tile_3_2_chanxy_out[44];
    assign wire_4963 = lut_tile_3_2_chanxy_out[45];
    assign wire_4971 = lut_tile_3_2_chanxy_out[46];
    assign wire_4979 = lut_tile_3_2_chanxy_out[47];
    assign wire_4987 = lut_tile_3_2_chanxy_out[48];
    assign wire_4995 = lut_tile_3_2_chanxy_out[49];
    assign wire_5003 = lut_tile_3_2_chanxy_out[50];
    assign wire_5011 = lut_tile_3_2_chanxy_out[51];
    assign wire_5019 = lut_tile_3_2_chanxy_out[52];
    assign wire_5027 = lut_tile_3_2_chanxy_out[53];
    assign wire_5035 = lut_tile_3_2_chanxy_out[54];
    assign wire_5043 = lut_tile_3_2_chanxy_out[55];
    assign wire_5051 = lut_tile_3_2_chanxy_out[56];
    assign wire_5059 = lut_tile_3_2_chanxy_out[57];
    assign wire_5067 = lut_tile_3_2_chanxy_out[58];
    assign wire_5075 = lut_tile_3_2_chanxy_out[59];
    assign wire_5120 = lut_tile_3_2_chanxy_out[60];
    assign wire_5122 = lut_tile_3_2_chanxy_out[61];
    assign wire_5124 = lut_tile_3_2_chanxy_out[62];
    assign wire_5126 = lut_tile_3_2_chanxy_out[63];
    assign wire_5128 = lut_tile_3_2_chanxy_out[64];
    assign wire_5130 = lut_tile_3_2_chanxy_out[65];
    assign wire_5132 = lut_tile_3_2_chanxy_out[66];
    assign wire_5134 = lut_tile_3_2_chanxy_out[67];
    assign wire_5136 = lut_tile_3_2_chanxy_out[68];
    assign wire_5138 = lut_tile_3_2_chanxy_out[69];
    assign wire_5140 = lut_tile_3_2_chanxy_out[70];
    assign wire_5142 = lut_tile_3_2_chanxy_out[71];
    assign wire_5144 = lut_tile_3_2_chanxy_out[72];
    assign wire_5146 = lut_tile_3_2_chanxy_out[73];
    assign wire_5148 = lut_tile_3_2_chanxy_out[74];
    assign wire_5150 = lut_tile_3_2_chanxy_out[75];
    assign wire_5152 = lut_tile_3_2_chanxy_out[76];
    assign wire_5154 = lut_tile_3_2_chanxy_out[77];
    assign wire_5156 = lut_tile_3_2_chanxy_out[78];
    assign wire_5158 = lut_tile_3_2_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_3_3_chanxy_in = {wire_5394, wire_3241, wire_3227, wire_3226, wire_3199, wire_3198, wire_3053, wire_3052, wire_3010, wire_1579, wire_1205, wire_5386, wire_3279, wire_3213, wire_3212, wire_3185, wire_3184, wire_3157, wire_3156, wire_3018, wire_1579, wire_1205, wire_5378, wire_3277, wire_3239, wire_3238, wire_3171, wire_3170, wire_3101, wire_3100, wire_3026, wire_1579, wire_1205, wire_5370, wire_3275, wire_3225, wire_3224, wire_3197, wire_3196, wire_3045, wire_3044, wire_3034, wire_1579, wire_1205, wire_5362, wire_3273, wire_3211, wire_3210, wire_3183, wire_3182, wire_3149, wire_3148, wire_3042, wire_1579, wire_1201, wire_5354, wire_3271, wire_3237, wire_3236, wire_3169, wire_3168, wire_3093, wire_3092, wire_3050, wire_1579, wire_1201, wire_5346, wire_3269, wire_3223, wire_3222, wire_3195, wire_3194, wire_3058, wire_3037, wire_3036, wire_1579, wire_1201, wire_5338, wire_3267, wire_3209, wire_3208, wire_3181, wire_3180, wire_3141, wire_3140, wire_3066, wire_1579, wire_1201, wire_5330, wire_3265, wire_3235, wire_3234, wire_3167, wire_3166, wire_3085, wire_3084, wire_3074, wire_1575, wire_1201, wire_5322, wire_3263, wire_3221, wire_3220, wire_3193, wire_3192, wire_3082, wire_3029, wire_3028, wire_1575, wire_1201, wire_5314, wire_3261, wire_3207, wire_3206, wire_3179, wire_3178, wire_3133, wire_3132, wire_3090, wire_1575, wire_1201, wire_5306, wire_3259, wire_3233, wire_3232, wire_3165, wire_3164, wire_3098, wire_3077, wire_3076, wire_1575, wire_1201, wire_5298, wire_3257, wire_3219, wire_3218, wire_3191, wire_3190, wire_3106, wire_3021, wire_3020, wire_1575, wire_1197, wire_5290, wire_3255, wire_3205, wire_3204, wire_3177, wire_3176, wire_3125, wire_3124, wire_3114, wire_1575, wire_1197, wire_5282, wire_3253, wire_3231, wire_3230, wire_3163, wire_3162, wire_3122, wire_3069, wire_3068, wire_1575, wire_1197, wire_5274, wire_3251, wire_3217, wire_3216, wire_3189, wire_3188, wire_3130, wire_3013, wire_3012, wire_1575, wire_1197, wire_5266, wire_3249, wire_3203, wire_3202, wire_3175, wire_3174, wire_3138, wire_3117, wire_3116, wire_1205, wire_1197, wire_5258, wire_3247, wire_3229, wire_3228, wire_3161, wire_3160, wire_3146, wire_3061, wire_3060, wire_1205, wire_1197, wire_5250, wire_3245, wire_3215, wire_3214, wire_3187, wire_3186, wire_3154, wire_3005, wire_3004, wire_1205, wire_1197, wire_5242, wire_3243, wire_3201, wire_3200, wire_3173, wire_3172, wire_3109, wire_3108, wire_3002, wire_1205, wire_1197, wire_5519, wire_3599, wire_3533, wire_3532, wire_3507, wire_3506, wire_3479, wire_3478, wire_3324, wire_1579, wire_1205, wire_5517, wire_3561, wire_3559, wire_3558, wire_3493, wire_3492, wire_3476, wire_3423, wire_3422, wire_1579, wire_1205, wire_5515, wire_3563, wire_3545, wire_3544, wire_3519, wire_3518, wire_3468, wire_3367, wire_3366, wire_1579, wire_1205, wire_5513, wire_3565, wire_3531, wire_3530, wire_3505, wire_3504, wire_3471, wire_3470, wire_3460, wire_1579, wire_1205, wire_5511, wire_3567, wire_3557, wire_3556, wire_3491, wire_3490, wire_3452, wire_3415, wire_3414, wire_1579, wire_1201, wire_5509, wire_3569, wire_3543, wire_3542, wire_3517, wire_3516, wire_3444, wire_3359, wire_3358, wire_1579, wire_1201, wire_5507, wire_3571, wire_3529, wire_3528, wire_3503, wire_3502, wire_3463, wire_3462, wire_3436, wire_1579, wire_1201, wire_5505, wire_3573, wire_3555, wire_3554, wire_3489, wire_3488, wire_3428, wire_3407, wire_3406, wire_1579, wire_1201, wire_5503, wire_3575, wire_3541, wire_3540, wire_3515, wire_3514, wire_3420, wire_3351, wire_3350, wire_1575, wire_1201, wire_5501, wire_3577, wire_3527, wire_3526, wire_3501, wire_3500, wire_3455, wire_3454, wire_3412, wire_1575, wire_1201, wire_5499, wire_3579, wire_3553, wire_3552, wire_3487, wire_3486, wire_3404, wire_3399, wire_3398, wire_1575, wire_1201, wire_5497, wire_3581, wire_3539, wire_3538, wire_3513, wire_3512, wire_3396, wire_3343, wire_3342, wire_1575, wire_1201, wire_5495, wire_3583, wire_3525, wire_3524, wire_3499, wire_3498, wire_3447, wire_3446, wire_3388, wire_1575, wire_1197, wire_5493, wire_3585, wire_3551, wire_3550, wire_3485, wire_3484, wire_3391, wire_3390, wire_3380, wire_1575, wire_1197, wire_5491, wire_3587, wire_3537, wire_3536, wire_3511, wire_3510, wire_3372, wire_3335, wire_3334, wire_1575, wire_1197, wire_5489, wire_3589, wire_3523, wire_3522, wire_3497, wire_3496, wire_3439, wire_3438, wire_3364, wire_1575, wire_1197, wire_5487, wire_3591, wire_3549, wire_3548, wire_3483, wire_3482, wire_3383, wire_3382, wire_3356, wire_1205, wire_1197, wire_5485, wire_3593, wire_3535, wire_3534, wire_3509, wire_3508, wire_3348, wire_3327, wire_3326, wire_1205, wire_1197, wire_5483, wire_3595, wire_3521, wire_3520, wire_3495, wire_3494, wire_3431, wire_3430, wire_3340, wire_1205, wire_1197, wire_5481, wire_3597, wire_3547, wire_3546, wire_3481, wire_3480, wire_3375, wire_3374, wire_3332, wire_1205, wire_1197, wire_5197, wire_5147, wire_5146, wire_5119, wire_5118, wire_5074, wire_4973, wire_4972, wire_3474, wire_1262, wire_1254, wire_5195, wire_5133, wire_5132, wire_5105, wire_5104, wire_5077, wire_5076, wire_4922, wire_3466, wire_1262, wire_1254, wire_5193, wire_5159, wire_5158, wire_5091, wire_5090, wire_5021, wire_5020, wire_4930, wire_3458, wire_1262, wire_1254, wire_5191, wire_5145, wire_5144, wire_5117, wire_5116, wire_4965, wire_4964, wire_4938, wire_3450, wire_1262, wire_1254, wire_5189, wire_5131, wire_5130, wire_5103, wire_5102, wire_5069, wire_5068, wire_4946, wire_3442, wire_1262, wire_1204, wire_5187, wire_5157, wire_5156, wire_5089, wire_5088, wire_5013, wire_5012, wire_4954, wire_3434, wire_1262, wire_1204, wire_5185, wire_5143, wire_5142, wire_5115, wire_5114, wire_4962, wire_4957, wire_4956, wire_3426, wire_1262, wire_1204, wire_5183, wire_5129, wire_5128, wire_5101, wire_5100, wire_5061, wire_5060, wire_4970, wire_3418, wire_1262, wire_1204, wire_5181, wire_5155, wire_5154, wire_5087, wire_5086, wire_5005, wire_5004, wire_4978, wire_3410, wire_1258, wire_1204, wire_5179, wire_5141, wire_5140, wire_5113, wire_5112, wire_4986, wire_4949, wire_4948, wire_3402, wire_1258, wire_1204, wire_5177, wire_5127, wire_5126, wire_5099, wire_5098, wire_5053, wire_5052, wire_4994, wire_3394, wire_1258, wire_1204, wire_5175, wire_5153, wire_5152, wire_5085, wire_5084, wire_5002, wire_4997, wire_4996, wire_3386, wire_1258, wire_1204, wire_5173, wire_5139, wire_5138, wire_5111, wire_5110, wire_5010, wire_4941, wire_4940, wire_3378, wire_1258, wire_1200, wire_5171, wire_5125, wire_5124, wire_5097, wire_5096, wire_5045, wire_5044, wire_5018, wire_3370, wire_1258, wire_1200, wire_5169, wire_5151, wire_5150, wire_5083, wire_5082, wire_5026, wire_4989, wire_4988, wire_3362, wire_1258, wire_1200, wire_5167, wire_5137, wire_5136, wire_5109, wire_5108, wire_5034, wire_4933, wire_4932, wire_3354, wire_1258, wire_1200, wire_5165, wire_5123, wire_5122, wire_5095, wire_5094, wire_5042, wire_5037, wire_5036, wire_3346, wire_1254, wire_1200, wire_5163, wire_5149, wire_5148, wire_5081, wire_5080, wire_5050, wire_4981, wire_4980, wire_3338, wire_1254, wire_1200, wire_5161, wire_5135, wire_5134, wire_5107, wire_5106, wire_5058, wire_4925, wire_4924, wire_3330, wire_1254, wire_1200, wire_5199, wire_5121, wire_5120, wire_5093, wire_5092, wire_5066, wire_5029, wire_5028, wire_3322, wire_1254, wire_1200, wire_5483, wire_5453, wire_5452, wire_5427, wire_5426, wire_5399, wire_5398, wire_5388, wire_3599, wire_1262, wire_1254, wire_5485, wire_5479, wire_5478, wire_5413, wire_5412, wire_5380, wire_5343, wire_5342, wire_3597, wire_1262, wire_1254, wire_5487, wire_5465, wire_5464, wire_5439, wire_5438, wire_5372, wire_5287, wire_5286, wire_3595, wire_1262, wire_1254, wire_5489, wire_5451, wire_5450, wire_5425, wire_5424, wire_5391, wire_5390, wire_5364, wire_3593, wire_1262, wire_1254, wire_5491, wire_5477, wire_5476, wire_5411, wire_5410, wire_5356, wire_5335, wire_5334, wire_3591, wire_1262, wire_1204, wire_5493, wire_5463, wire_5462, wire_5437, wire_5436, wire_5348, wire_5279, wire_5278, wire_3589, wire_1262, wire_1204, wire_5495, wire_5449, wire_5448, wire_5423, wire_5422, wire_5383, wire_5382, wire_5340, wire_3587, wire_1262, wire_1204, wire_5497, wire_5475, wire_5474, wire_5409, wire_5408, wire_5332, wire_5327, wire_5326, wire_3585, wire_1262, wire_1204, wire_5499, wire_5461, wire_5460, wire_5435, wire_5434, wire_5324, wire_5271, wire_5270, wire_3583, wire_1258, wire_1204, wire_5501, wire_5447, wire_5446, wire_5421, wire_5420, wire_5375, wire_5374, wire_5316, wire_3581, wire_1258, wire_1204, wire_5503, wire_5473, wire_5472, wire_5407, wire_5406, wire_5319, wire_5318, wire_5308, wire_3579, wire_1258, wire_1204, wire_5505, wire_5459, wire_5458, wire_5433, wire_5432, wire_5300, wire_5263, wire_5262, wire_3577, wire_1258, wire_1204, wire_5507, wire_5445, wire_5444, wire_5419, wire_5418, wire_5367, wire_5366, wire_5292, wire_3575, wire_1258, wire_1200, wire_5509, wire_5471, wire_5470, wire_5405, wire_5404, wire_5311, wire_5310, wire_5284, wire_3573, wire_1258, wire_1200, wire_5511, wire_5457, wire_5456, wire_5431, wire_5430, wire_5276, wire_5255, wire_5254, wire_3571, wire_1258, wire_1200, wire_5513, wire_5443, wire_5442, wire_5417, wire_5416, wire_5359, wire_5358, wire_5268, wire_3569, wire_1258, wire_1200, wire_5515, wire_5469, wire_5468, wire_5403, wire_5402, wire_5303, wire_5302, wire_5260, wire_3567, wire_1254, wire_1200, wire_5517, wire_5455, wire_5454, wire_5429, wire_5428, wire_5252, wire_5247, wire_5246, wire_3565, wire_1254, wire_1200, wire_5519, wire_5441, wire_5440, wire_5415, wire_5414, wire_5351, wire_5350, wire_5244, wire_3563, wire_1254, wire_1200, wire_5481, wire_5467, wire_5466, wire_5401, wire_5400, wire_5396, wire_5295, wire_5294, wire_3561, wire_1254, wire_1200};
    // CHNAXY TOTAL: 880
    assign wire_3325 = lut_tile_3_3_chanxy_out[0];
    assign wire_3333 = lut_tile_3_3_chanxy_out[1];
    assign wire_3341 = lut_tile_3_3_chanxy_out[2];
    assign wire_3349 = lut_tile_3_3_chanxy_out[3];
    assign wire_3357 = lut_tile_3_3_chanxy_out[4];
    assign wire_3365 = lut_tile_3_3_chanxy_out[5];
    assign wire_3373 = lut_tile_3_3_chanxy_out[6];
    assign wire_3381 = lut_tile_3_3_chanxy_out[7];
    assign wire_3389 = lut_tile_3_3_chanxy_out[8];
    assign wire_3397 = lut_tile_3_3_chanxy_out[9];
    assign wire_3405 = lut_tile_3_3_chanxy_out[10];
    assign wire_3413 = lut_tile_3_3_chanxy_out[11];
    assign wire_3421 = lut_tile_3_3_chanxy_out[12];
    assign wire_3429 = lut_tile_3_3_chanxy_out[13];
    assign wire_3437 = lut_tile_3_3_chanxy_out[14];
    assign wire_3445 = lut_tile_3_3_chanxy_out[15];
    assign wire_3453 = lut_tile_3_3_chanxy_out[16];
    assign wire_3461 = lut_tile_3_3_chanxy_out[17];
    assign wire_3469 = lut_tile_3_3_chanxy_out[18];
    assign wire_3477 = lut_tile_3_3_chanxy_out[19];
    assign wire_3520 = lut_tile_3_3_chanxy_out[20];
    assign wire_3522 = lut_tile_3_3_chanxy_out[21];
    assign wire_3524 = lut_tile_3_3_chanxy_out[22];
    assign wire_3526 = lut_tile_3_3_chanxy_out[23];
    assign wire_3528 = lut_tile_3_3_chanxy_out[24];
    assign wire_3530 = lut_tile_3_3_chanxy_out[25];
    assign wire_3532 = lut_tile_3_3_chanxy_out[26];
    assign wire_3534 = lut_tile_3_3_chanxy_out[27];
    assign wire_3536 = lut_tile_3_3_chanxy_out[28];
    assign wire_3538 = lut_tile_3_3_chanxy_out[29];
    assign wire_3540 = lut_tile_3_3_chanxy_out[30];
    assign wire_3542 = lut_tile_3_3_chanxy_out[31];
    assign wire_3544 = lut_tile_3_3_chanxy_out[32];
    assign wire_3546 = lut_tile_3_3_chanxy_out[33];
    assign wire_3548 = lut_tile_3_3_chanxy_out[34];
    assign wire_3550 = lut_tile_3_3_chanxy_out[35];
    assign wire_3552 = lut_tile_3_3_chanxy_out[36];
    assign wire_3554 = lut_tile_3_3_chanxy_out[37];
    assign wire_3556 = lut_tile_3_3_chanxy_out[38];
    assign wire_3558 = lut_tile_3_3_chanxy_out[39];
    assign wire_5245 = lut_tile_3_3_chanxy_out[40];
    assign wire_5253 = lut_tile_3_3_chanxy_out[41];
    assign wire_5261 = lut_tile_3_3_chanxy_out[42];
    assign wire_5269 = lut_tile_3_3_chanxy_out[43];
    assign wire_5277 = lut_tile_3_3_chanxy_out[44];
    assign wire_5285 = lut_tile_3_3_chanxy_out[45];
    assign wire_5293 = lut_tile_3_3_chanxy_out[46];
    assign wire_5301 = lut_tile_3_3_chanxy_out[47];
    assign wire_5309 = lut_tile_3_3_chanxy_out[48];
    assign wire_5317 = lut_tile_3_3_chanxy_out[49];
    assign wire_5325 = lut_tile_3_3_chanxy_out[50];
    assign wire_5333 = lut_tile_3_3_chanxy_out[51];
    assign wire_5341 = lut_tile_3_3_chanxy_out[52];
    assign wire_5349 = lut_tile_3_3_chanxy_out[53];
    assign wire_5357 = lut_tile_3_3_chanxy_out[54];
    assign wire_5365 = lut_tile_3_3_chanxy_out[55];
    assign wire_5373 = lut_tile_3_3_chanxy_out[56];
    assign wire_5381 = lut_tile_3_3_chanxy_out[57];
    assign wire_5389 = lut_tile_3_3_chanxy_out[58];
    assign wire_5397 = lut_tile_3_3_chanxy_out[59];
    assign wire_5440 = lut_tile_3_3_chanxy_out[60];
    assign wire_5442 = lut_tile_3_3_chanxy_out[61];
    assign wire_5444 = lut_tile_3_3_chanxy_out[62];
    assign wire_5446 = lut_tile_3_3_chanxy_out[63];
    assign wire_5448 = lut_tile_3_3_chanxy_out[64];
    assign wire_5450 = lut_tile_3_3_chanxy_out[65];
    assign wire_5452 = lut_tile_3_3_chanxy_out[66];
    assign wire_5454 = lut_tile_3_3_chanxy_out[67];
    assign wire_5456 = lut_tile_3_3_chanxy_out[68];
    assign wire_5458 = lut_tile_3_3_chanxy_out[69];
    assign wire_5460 = lut_tile_3_3_chanxy_out[70];
    assign wire_5462 = lut_tile_3_3_chanxy_out[71];
    assign wire_5464 = lut_tile_3_3_chanxy_out[72];
    assign wire_5466 = lut_tile_3_3_chanxy_out[73];
    assign wire_5468 = lut_tile_3_3_chanxy_out[74];
    assign wire_5470 = lut_tile_3_3_chanxy_out[75];
    assign wire_5472 = lut_tile_3_3_chanxy_out[76];
    assign wire_5474 = lut_tile_3_3_chanxy_out[77];
    assign wire_5476 = lut_tile_3_3_chanxy_out[78];
    assign wire_5478 = lut_tile_3_3_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_3_4_chanxy_in = {wire_5716, wire_3281, wire_3253, wire_3252, wire_3227, wire_3226, wire_3199, wire_3198, wire_3012, wire_1955, wire_1581, wire_5708, wire_3319, wire_3279, wire_3278, wire_3213, wire_3212, wire_3185, wire_3184, wire_3020, wire_1955, wire_1581, wire_5700, wire_3317, wire_3265, wire_3264, wire_3239, wire_3238, wire_3171, wire_3170, wire_3028, wire_1955, wire_1581, wire_5692, wire_3315, wire_3251, wire_3250, wire_3225, wire_3224, wire_3197, wire_3196, wire_3036, wire_1955, wire_1581, wire_5684, wire_3313, wire_3277, wire_3276, wire_3211, wire_3210, wire_3183, wire_3182, wire_3044, wire_1955, wire_1577, wire_5676, wire_3311, wire_3263, wire_3262, wire_3237, wire_3236, wire_3169, wire_3168, wire_3052, wire_1955, wire_1577, wire_5668, wire_3309, wire_3249, wire_3248, wire_3223, wire_3222, wire_3195, wire_3194, wire_3060, wire_1955, wire_1577, wire_5660, wire_3307, wire_3275, wire_3274, wire_3209, wire_3208, wire_3181, wire_3180, wire_3068, wire_1955, wire_1577, wire_5652, wire_3305, wire_3261, wire_3260, wire_3235, wire_3234, wire_3167, wire_3166, wire_3076, wire_1951, wire_1577, wire_5644, wire_3303, wire_3247, wire_3246, wire_3221, wire_3220, wire_3193, wire_3192, wire_3084, wire_1951, wire_1577, wire_5636, wire_3301, wire_3273, wire_3272, wire_3207, wire_3206, wire_3179, wire_3178, wire_3092, wire_1951, wire_1577, wire_5628, wire_3299, wire_3259, wire_3258, wire_3233, wire_3232, wire_3165, wire_3164, wire_3100, wire_1951, wire_1577, wire_5620, wire_3297, wire_3245, wire_3244, wire_3219, wire_3218, wire_3191, wire_3190, wire_3108, wire_1951, wire_1573, wire_5612, wire_3295, wire_3271, wire_3270, wire_3205, wire_3204, wire_3177, wire_3176, wire_3116, wire_1951, wire_1573, wire_5604, wire_3293, wire_3257, wire_3256, wire_3231, wire_3230, wire_3163, wire_3162, wire_3124, wire_1951, wire_1573, wire_5596, wire_3291, wire_3243, wire_3242, wire_3217, wire_3216, wire_3189, wire_3188, wire_3132, wire_1951, wire_1573, wire_5588, wire_3289, wire_3269, wire_3268, wire_3203, wire_3202, wire_3175, wire_3174, wire_3140, wire_1581, wire_1573, wire_5580, wire_3287, wire_3255, wire_3254, wire_3229, wire_3228, wire_3161, wire_3160, wire_3148, wire_1581, wire_1573, wire_5572, wire_3285, wire_3241, wire_3240, wire_3215, wire_3214, wire_3187, wire_3186, wire_3156, wire_1581, wire_1573, wire_5564, wire_3283, wire_3267, wire_3266, wire_3201, wire_3200, wire_3173, wire_3172, wire_3004, wire_1581, wire_1573, wire_5839, wire_3639, wire_3599, wire_3598, wire_3533, wire_3532, wire_3507, wire_3506, wire_3326, wire_1955, wire_1581, wire_5837, wire_3601, wire_3585, wire_3584, wire_3559, wire_3558, wire_3493, wire_3492, wire_3478, wire_1955, wire_1581, wire_5835, wire_3603, wire_3571, wire_3570, wire_3545, wire_3544, wire_3519, wire_3518, wire_3470, wire_1955, wire_1581, wire_5833, wire_3605, wire_3597, wire_3596, wire_3531, wire_3530, wire_3505, wire_3504, wire_3462, wire_1955, wire_1581, wire_5831, wire_3607, wire_3583, wire_3582, wire_3557, wire_3556, wire_3491, wire_3490, wire_3454, wire_1955, wire_1577, wire_5829, wire_3609, wire_3569, wire_3568, wire_3543, wire_3542, wire_3517, wire_3516, wire_3446, wire_1955, wire_1577, wire_5827, wire_3611, wire_3595, wire_3594, wire_3529, wire_3528, wire_3503, wire_3502, wire_3438, wire_1955, wire_1577, wire_5825, wire_3613, wire_3581, wire_3580, wire_3555, wire_3554, wire_3489, wire_3488, wire_3430, wire_1955, wire_1577, wire_5823, wire_3615, wire_3567, wire_3566, wire_3541, wire_3540, wire_3515, wire_3514, wire_3422, wire_1951, wire_1577, wire_5821, wire_3617, wire_3593, wire_3592, wire_3527, wire_3526, wire_3501, wire_3500, wire_3414, wire_1951, wire_1577, wire_5819, wire_3619, wire_3579, wire_3578, wire_3553, wire_3552, wire_3487, wire_3486, wire_3406, wire_1951, wire_1577, wire_5817, wire_3621, wire_3565, wire_3564, wire_3539, wire_3538, wire_3513, wire_3512, wire_3398, wire_1951, wire_1577, wire_5815, wire_3623, wire_3591, wire_3590, wire_3525, wire_3524, wire_3499, wire_3498, wire_3390, wire_1951, wire_1573, wire_5813, wire_3625, wire_3577, wire_3576, wire_3551, wire_3550, wire_3485, wire_3484, wire_3382, wire_1951, wire_1573, wire_5811, wire_3627, wire_3563, wire_3562, wire_3537, wire_3536, wire_3511, wire_3510, wire_3374, wire_1951, wire_1573, wire_5809, wire_3629, wire_3589, wire_3588, wire_3523, wire_3522, wire_3497, wire_3496, wire_3366, wire_1951, wire_1573, wire_5807, wire_3631, wire_3575, wire_3574, wire_3549, wire_3548, wire_3483, wire_3482, wire_3358, wire_1581, wire_1573, wire_5805, wire_3633, wire_3561, wire_3560, wire_3535, wire_3534, wire_3509, wire_3508, wire_3350, wire_1581, wire_1573, wire_5803, wire_3635, wire_3587, wire_3586, wire_3521, wire_3520, wire_3495, wire_3494, wire_3342, wire_1581, wire_1573, wire_5801, wire_3637, wire_3573, wire_3572, wire_3547, wire_3546, wire_3481, wire_3480, wire_3334, wire_1581, wire_1573, wire_5517, wire_5453, wire_5452, wire_5427, wire_5426, wire_5399, wire_5398, wire_5396, wire_3476, wire_1638, wire_1630, wire_5515, wire_5479, wire_5478, wire_5413, wire_5412, wire_5343, wire_5342, wire_5244, wire_3468, wire_1638, wire_1630, wire_5513, wire_5465, wire_5464, wire_5439, wire_5438, wire_5287, wire_5286, wire_5252, wire_3460, wire_1638, wire_1630, wire_5511, wire_5451, wire_5450, wire_5425, wire_5424, wire_5391, wire_5390, wire_5260, wire_3452, wire_1638, wire_1630, wire_5509, wire_5477, wire_5476, wire_5411, wire_5410, wire_5335, wire_5334, wire_5268, wire_3444, wire_1638, wire_1580, wire_5507, wire_5463, wire_5462, wire_5437, wire_5436, wire_5279, wire_5278, wire_5276, wire_3436, wire_1638, wire_1580, wire_5505, wire_5449, wire_5448, wire_5423, wire_5422, wire_5383, wire_5382, wire_5284, wire_3428, wire_1638, wire_1580, wire_5503, wire_5475, wire_5474, wire_5409, wire_5408, wire_5327, wire_5326, wire_5292, wire_3420, wire_1638, wire_1580, wire_5501, wire_5461, wire_5460, wire_5435, wire_5434, wire_5300, wire_5271, wire_5270, wire_3412, wire_1634, wire_1580, wire_5499, wire_5447, wire_5446, wire_5421, wire_5420, wire_5375, wire_5374, wire_5308, wire_3404, wire_1634, wire_1580, wire_5497, wire_5473, wire_5472, wire_5407, wire_5406, wire_5319, wire_5318, wire_5316, wire_3396, wire_1634, wire_1580, wire_5495, wire_5459, wire_5458, wire_5433, wire_5432, wire_5324, wire_5263, wire_5262, wire_3388, wire_1634, wire_1580, wire_5493, wire_5445, wire_5444, wire_5419, wire_5418, wire_5367, wire_5366, wire_5332, wire_3380, wire_1634, wire_1576, wire_5491, wire_5471, wire_5470, wire_5405, wire_5404, wire_5340, wire_5311, wire_5310, wire_3372, wire_1634, wire_1576, wire_5489, wire_5457, wire_5456, wire_5431, wire_5430, wire_5348, wire_5255, wire_5254, wire_3364, wire_1634, wire_1576, wire_5487, wire_5443, wire_5442, wire_5417, wire_5416, wire_5359, wire_5358, wire_5356, wire_3356, wire_1634, wire_1576, wire_5485, wire_5469, wire_5468, wire_5403, wire_5402, wire_5364, wire_5303, wire_5302, wire_3348, wire_1630, wire_1576, wire_5483, wire_5455, wire_5454, wire_5429, wire_5428, wire_5372, wire_5247, wire_5246, wire_3340, wire_1630, wire_1576, wire_5481, wire_5441, wire_5440, wire_5415, wire_5414, wire_5380, wire_5351, wire_5350, wire_3332, wire_1630, wire_1576, wire_5519, wire_5467, wire_5466, wire_5401, wire_5400, wire_5388, wire_5295, wire_5294, wire_3324, wire_1630, wire_1576, wire_5803, wire_5799, wire_5798, wire_5733, wire_5732, wire_5710, wire_5665, wire_5664, wire_3639, wire_1638, wire_1630, wire_5805, wire_5785, wire_5784, wire_5759, wire_5758, wire_5702, wire_5609, wire_5608, wire_3637, wire_1638, wire_1630, wire_5807, wire_5771, wire_5770, wire_5745, wire_5744, wire_5713, wire_5712, wire_5694, wire_3635, wire_1638, wire_1630, wire_5809, wire_5797, wire_5796, wire_5731, wire_5730, wire_5686, wire_5657, wire_5656, wire_3633, wire_1638, wire_1630, wire_5811, wire_5783, wire_5782, wire_5757, wire_5756, wire_5678, wire_5601, wire_5600, wire_3631, wire_1638, wire_1580, wire_5813, wire_5769, wire_5768, wire_5743, wire_5742, wire_5705, wire_5704, wire_5670, wire_3629, wire_1638, wire_1580, wire_5815, wire_5795, wire_5794, wire_5729, wire_5728, wire_5662, wire_5649, wire_5648, wire_3627, wire_1638, wire_1580, wire_5817, wire_5781, wire_5780, wire_5755, wire_5754, wire_5654, wire_5593, wire_5592, wire_3625, wire_1638, wire_1580, wire_5819, wire_5767, wire_5766, wire_5741, wire_5740, wire_5697, wire_5696, wire_5646, wire_3623, wire_1634, wire_1580, wire_5821, wire_5793, wire_5792, wire_5727, wire_5726, wire_5641, wire_5640, wire_5638, wire_3621, wire_1634, wire_1580, wire_5823, wire_5779, wire_5778, wire_5753, wire_5752, wire_5630, wire_5585, wire_5584, wire_3619, wire_1634, wire_1580, wire_5825, wire_5765, wire_5764, wire_5739, wire_5738, wire_5689, wire_5688, wire_5622, wire_3617, wire_1634, wire_1580, wire_5827, wire_5791, wire_5790, wire_5725, wire_5724, wire_5633, wire_5632, wire_5614, wire_3615, wire_1634, wire_1576, wire_5829, wire_5777, wire_5776, wire_5751, wire_5750, wire_5606, wire_5577, wire_5576, wire_3613, wire_1634, wire_1576, wire_5831, wire_5763, wire_5762, wire_5737, wire_5736, wire_5681, wire_5680, wire_5598, wire_3611, wire_1634, wire_1576, wire_5833, wire_5789, wire_5788, wire_5723, wire_5722, wire_5625, wire_5624, wire_5590, wire_3609, wire_1634, wire_1576, wire_5835, wire_5775, wire_5774, wire_5749, wire_5748, wire_5582, wire_5569, wire_5568, wire_3607, wire_1630, wire_1576, wire_5837, wire_5761, wire_5760, wire_5735, wire_5734, wire_5673, wire_5672, wire_5574, wire_3605, wire_1630, wire_1576, wire_5839, wire_5787, wire_5786, wire_5721, wire_5720, wire_5617, wire_5616, wire_5566, wire_3603, wire_1630, wire_1576, wire_5801, wire_5773, wire_5772, wire_5747, wire_5746, wire_5718, wire_5561, wire_5560, wire_3601, wire_1630, wire_1576};
    // CHNAXY TOTAL: 880
    assign wire_3327 = lut_tile_3_4_chanxy_out[0];
    assign wire_3335 = lut_tile_3_4_chanxy_out[1];
    assign wire_3343 = lut_tile_3_4_chanxy_out[2];
    assign wire_3351 = lut_tile_3_4_chanxy_out[3];
    assign wire_3359 = lut_tile_3_4_chanxy_out[4];
    assign wire_3367 = lut_tile_3_4_chanxy_out[5];
    assign wire_3375 = lut_tile_3_4_chanxy_out[6];
    assign wire_3383 = lut_tile_3_4_chanxy_out[7];
    assign wire_3391 = lut_tile_3_4_chanxy_out[8];
    assign wire_3399 = lut_tile_3_4_chanxy_out[9];
    assign wire_3407 = lut_tile_3_4_chanxy_out[10];
    assign wire_3415 = lut_tile_3_4_chanxy_out[11];
    assign wire_3423 = lut_tile_3_4_chanxy_out[12];
    assign wire_3431 = lut_tile_3_4_chanxy_out[13];
    assign wire_3439 = lut_tile_3_4_chanxy_out[14];
    assign wire_3447 = lut_tile_3_4_chanxy_out[15];
    assign wire_3455 = lut_tile_3_4_chanxy_out[16];
    assign wire_3463 = lut_tile_3_4_chanxy_out[17];
    assign wire_3471 = lut_tile_3_4_chanxy_out[18];
    assign wire_3479 = lut_tile_3_4_chanxy_out[19];
    assign wire_3560 = lut_tile_3_4_chanxy_out[20];
    assign wire_3562 = lut_tile_3_4_chanxy_out[21];
    assign wire_3564 = lut_tile_3_4_chanxy_out[22];
    assign wire_3566 = lut_tile_3_4_chanxy_out[23];
    assign wire_3568 = lut_tile_3_4_chanxy_out[24];
    assign wire_3570 = lut_tile_3_4_chanxy_out[25];
    assign wire_3572 = lut_tile_3_4_chanxy_out[26];
    assign wire_3574 = lut_tile_3_4_chanxy_out[27];
    assign wire_3576 = lut_tile_3_4_chanxy_out[28];
    assign wire_3578 = lut_tile_3_4_chanxy_out[29];
    assign wire_3580 = lut_tile_3_4_chanxy_out[30];
    assign wire_3582 = lut_tile_3_4_chanxy_out[31];
    assign wire_3584 = lut_tile_3_4_chanxy_out[32];
    assign wire_3586 = lut_tile_3_4_chanxy_out[33];
    assign wire_3588 = lut_tile_3_4_chanxy_out[34];
    assign wire_3590 = lut_tile_3_4_chanxy_out[35];
    assign wire_3592 = lut_tile_3_4_chanxy_out[36];
    assign wire_3594 = lut_tile_3_4_chanxy_out[37];
    assign wire_3596 = lut_tile_3_4_chanxy_out[38];
    assign wire_3598 = lut_tile_3_4_chanxy_out[39];
    assign wire_5567 = lut_tile_3_4_chanxy_out[40];
    assign wire_5575 = lut_tile_3_4_chanxy_out[41];
    assign wire_5583 = lut_tile_3_4_chanxy_out[42];
    assign wire_5591 = lut_tile_3_4_chanxy_out[43];
    assign wire_5599 = lut_tile_3_4_chanxy_out[44];
    assign wire_5607 = lut_tile_3_4_chanxy_out[45];
    assign wire_5615 = lut_tile_3_4_chanxy_out[46];
    assign wire_5623 = lut_tile_3_4_chanxy_out[47];
    assign wire_5631 = lut_tile_3_4_chanxy_out[48];
    assign wire_5639 = lut_tile_3_4_chanxy_out[49];
    assign wire_5647 = lut_tile_3_4_chanxy_out[50];
    assign wire_5655 = lut_tile_3_4_chanxy_out[51];
    assign wire_5663 = lut_tile_3_4_chanxy_out[52];
    assign wire_5671 = lut_tile_3_4_chanxy_out[53];
    assign wire_5679 = lut_tile_3_4_chanxy_out[54];
    assign wire_5687 = lut_tile_3_4_chanxy_out[55];
    assign wire_5695 = lut_tile_3_4_chanxy_out[56];
    assign wire_5703 = lut_tile_3_4_chanxy_out[57];
    assign wire_5711 = lut_tile_3_4_chanxy_out[58];
    assign wire_5719 = lut_tile_3_4_chanxy_out[59];
    assign wire_5760 = lut_tile_3_4_chanxy_out[60];
    assign wire_5762 = lut_tile_3_4_chanxy_out[61];
    assign wire_5764 = lut_tile_3_4_chanxy_out[62];
    assign wire_5766 = lut_tile_3_4_chanxy_out[63];
    assign wire_5768 = lut_tile_3_4_chanxy_out[64];
    assign wire_5770 = lut_tile_3_4_chanxy_out[65];
    assign wire_5772 = lut_tile_3_4_chanxy_out[66];
    assign wire_5774 = lut_tile_3_4_chanxy_out[67];
    assign wire_5776 = lut_tile_3_4_chanxy_out[68];
    assign wire_5778 = lut_tile_3_4_chanxy_out[69];
    assign wire_5780 = lut_tile_3_4_chanxy_out[70];
    assign wire_5782 = lut_tile_3_4_chanxy_out[71];
    assign wire_5784 = lut_tile_3_4_chanxy_out[72];
    assign wire_5786 = lut_tile_3_4_chanxy_out[73];
    assign wire_5788 = lut_tile_3_4_chanxy_out[74];
    assign wire_5790 = lut_tile_3_4_chanxy_out[75];
    assign wire_5792 = lut_tile_3_4_chanxy_out[76];
    assign wire_5794 = lut_tile_3_4_chanxy_out[77];
    assign wire_5796 = lut_tile_3_4_chanxy_out[78];
    assign wire_5798 = lut_tile_3_4_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_3_5_chanxy_in = {wire_6038, wire_3198, wire_3188, wire_3178, wire_3168, wire_2259, wire_2253, wire_2244, wire_1957, wire_6030, wire_3318, wire_3308, wire_3298, wire_3288, wire_2259, wire_2253, wire_2244, wire_1957, wire_6022, wire_3278, wire_3268, wire_3258, wire_3248, wire_2259, wire_2253, wire_2244, wire_1957, wire_6014, wire_3238, wire_3228, wire_3218, wire_3208, wire_2259, wire_2253, wire_2244, wire_1957, wire_6006, wire_3196, wire_3186, wire_3176, wire_3166, wire_2259, wire_2250, wire_2244, wire_1953, wire_5998, wire_3316, wire_3306, wire_3296, wire_3286, wire_2259, wire_2250, wire_2244, wire_1953, wire_5990, wire_3276, wire_3266, wire_3256, wire_3246, wire_2259, wire_2250, wire_2244, wire_1953, wire_5982, wire_3236, wire_3226, wire_3216, wire_3206, wire_2259, wire_2250, wire_2244, wire_1953, wire_5974, wire_3194, wire_3184, wire_3174, wire_3164, wire_2256, wire_2250, wire_2241, wire_1953, wire_5966, wire_3314, wire_3304, wire_3294, wire_3284, wire_2256, wire_2250, wire_2241, wire_1953, wire_5958, wire_3274, wire_3264, wire_3254, wire_3244, wire_2256, wire_2250, wire_2241, wire_1953, wire_5950, wire_3234, wire_3224, wire_3214, wire_3204, wire_2256, wire_2250, wire_2241, wire_1953, wire_5942, wire_3192, wire_3182, wire_3172, wire_3162, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_5934, wire_3312, wire_3302, wire_3292, wire_3282, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_5926, wire_3272, wire_3262, wire_3252, wire_3242, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_5918, wire_3232, wire_3222, wire_3212, wire_3202, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_5910, wire_3190, wire_3180, wire_3170, wire_3160, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_5902, wire_3310, wire_3300, wire_3290, wire_3280, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_5894, wire_3270, wire_3260, wire_3250, wire_3240, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_5886, wire_3230, wire_3220, wire_3210, wire_3200, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_6159, wire_3638, wire_3628, wire_3618, wire_3608, wire_2259, wire_2253, wire_2244, wire_1957, wire_6157, wire_3598, wire_3588, wire_3578, wire_3568, wire_2259, wire_2253, wire_2244, wire_1957, wire_6155, wire_3558, wire_3548, wire_3538, wire_3528, wire_2259, wire_2253, wire_2244, wire_1957, wire_6153, wire_3518, wire_3508, wire_3498, wire_3488, wire_2259, wire_2253, wire_2244, wire_1957, wire_6151, wire_3636, wire_3626, wire_3616, wire_3606, wire_2259, wire_2250, wire_2244, wire_1953, wire_6149, wire_3596, wire_3586, wire_3576, wire_3566, wire_2259, wire_2250, wire_2244, wire_1953, wire_6147, wire_3556, wire_3546, wire_3536, wire_3526, wire_2259, wire_2250, wire_2244, wire_1953, wire_6145, wire_3516, wire_3506, wire_3496, wire_3486, wire_2259, wire_2250, wire_2244, wire_1953, wire_6143, wire_3634, wire_3624, wire_3614, wire_3604, wire_2256, wire_2250, wire_2241, wire_1953, wire_6141, wire_3594, wire_3584, wire_3574, wire_3564, wire_2256, wire_2250, wire_2241, wire_1953, wire_6139, wire_3554, wire_3544, wire_3534, wire_3524, wire_2256, wire_2250, wire_2241, wire_1953, wire_6137, wire_3514, wire_3504, wire_3494, wire_3484, wire_2256, wire_2250, wire_2241, wire_1953, wire_6135, wire_3632, wire_3622, wire_3612, wire_3602, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_6133, wire_3592, wire_3582, wire_3572, wire_3562, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_6131, wire_3552, wire_3542, wire_3532, wire_3522, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_6129, wire_3512, wire_3502, wire_3492, wire_3482, wire_2262, wire_2256, wire_2247, wire_2241, wire_1949, wire_6127, wire_3630, wire_3620, wire_3610, wire_3600, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_6125, wire_3590, wire_3580, wire_3570, wire_3560, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_6123, wire_3550, wire_3540, wire_3530, wire_3520, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_6121, wire_3510, wire_3500, wire_3490, wire_3480, wire_2262, wire_2253, wire_2247, wire_1957, wire_1949, wire_6119, wire_6118, wire_5837, wire_5799, wire_5798, wire_5733, wire_5732, wire_5718, wire_5665, wire_5664, wire_3478, wire_2014, wire_2006, wire_5955, wire_5954, wire_5835, wire_5785, wire_5784, wire_5759, wire_5758, wire_5609, wire_5608, wire_5566, wire_3470, wire_2014, wire_2006, wire_6097, wire_6096, wire_5833, wire_5771, wire_5770, wire_5745, wire_5744, wire_5713, wire_5712, wire_5574, wire_3462, wire_2014, wire_2006, wire_6137, wire_5944, wire_5831, wire_5797, wire_5796, wire_5731, wire_5730, wire_5657, wire_5656, wire_5582, wire_3454, wire_2014, wire_2006, wire_6157, wire_6024, wire_5829, wire_5783, wire_5782, wire_5757, wire_5756, wire_5601, wire_5600, wire_5590, wire_3446, wire_2014, wire_1956, wire_6075, wire_6074, wire_5827, wire_5769, wire_5768, wire_5743, wire_5742, wire_5705, wire_5704, wire_5598, wire_3438, wire_2014, wire_1956, wire_6113, wire_6112, wire_5825, wire_5795, wire_5794, wire_5729, wire_5728, wire_5649, wire_5648, wire_5606, wire_3430, wire_2014, wire_1956, wire_5931, wire_5930, wire_5823, wire_5781, wire_5780, wire_5755, wire_5754, wire_5614, wire_5593, wire_5592, wire_3422, wire_2014, wire_1956, wire_6091, wire_6090, wire_5821, wire_5767, wire_5766, wire_5741, wire_5740, wire_5697, wire_5696, wire_5622, wire_3414, wire_2010, wire_1956, wire_6131, wire_5920, wire_5819, wire_5793, wire_5792, wire_5727, wire_5726, wire_5641, wire_5640, wire_5630, wire_3406, wire_2010, wire_1956, wire_6151, wire_6000, wire_2014, wire_5817, wire_5779, wire_5778, wire_5753, wire_5752, wire_5638, wire_5585, wire_5584, wire_3398, wire_2010, wire_1956, wire_6069, wire_6068, wire_2014, wire_5815, wire_5765, wire_5764, wire_5739, wire_5738, wire_5689, wire_5688, wire_5646, wire_3390, wire_2010, wire_1956, wire_6107, wire_6106, wire_2010, wire_5813, wire_5791, wire_5790, wire_5725, wire_5724, wire_5654, wire_5633, wire_5632, wire_3382, wire_2010, wire_1952, wire_5907, wire_5906, wire_2010, wire_5811, wire_5777, wire_5776, wire_5751, wire_5750, wire_5662, wire_5577, wire_5576, wire_3374, wire_2010, wire_1952, wire_6085, wire_6084, wire_2006, wire_5809, wire_5763, wire_5762, wire_5737, wire_5736, wire_5681, wire_5680, wire_5670, wire_3366, wire_2010, wire_1952, wire_6125, wire_5896, wire_2006, wire_5807, wire_5789, wire_5788, wire_5723, wire_5722, wire_5678, wire_5625, wire_5624, wire_3358, wire_2010, wire_1952, wire_6145, wire_5976, wire_1956, wire_5805, wire_5775, wire_5774, wire_5749, wire_5748, wire_5686, wire_5569, wire_5568, wire_3350, wire_2006, wire_1952, wire_6063, wire_6062, wire_1956, wire_5803, wire_5761, wire_5760, wire_5735, wire_5734, wire_5694, wire_5673, wire_5672, wire_3342, wire_2006, wire_1952, wire_6101, wire_6100, wire_1952, wire_5801, wire_5787, wire_5786, wire_5721, wire_5720, wire_5702, wire_5617, wire_5616, wire_3334, wire_2006, wire_1952, wire_5883, wire_5882, wire_1952, wire_5839, wire_5773, wire_5772, wire_5747, wire_5746, wire_5710, wire_5561, wire_5560, wire_3326, wire_2006, wire_1952, wire_6059, wire_6058, wire_6159, wire_6032, wire_6057, wire_6056, wire_6027, wire_6026, wire_5939, wire_5938, wire_6019, wire_6018, wire_6053, wire_6052, wire_6153, wire_6008, wire_6051, wire_6050, wire_6003, wire_6002, wire_5915, wire_5914, wire_2014, wire_5995, wire_5994, wire_2014, wire_6047, wire_6046, wire_2010, wire_6147, wire_5984, wire_2010, wire_6045, wire_6044, wire_2006, wire_5979, wire_5978, wire_2006, wire_5891, wire_5890, wire_1956, wire_5971, wire_5970, wire_1956, wire_6041, wire_6040, wire_1952, wire_6141, wire_5960, wire_1952, wire_6079, wire_6078, wire_6117, wire_6116, wire_6077, wire_6076, wire_6095, wire_6094, wire_6135, wire_5936, wire_6093, wire_6092, wire_6073, wire_6072, wire_6111, wire_6110, wire_6071, wire_6070, wire_6089, wire_6088, wire_6129, wire_5912, wire_2014, wire_6087, wire_6086, wire_2014, wire_6067, wire_6066, wire_2010, wire_6105, wire_6104, wire_2010, wire_6065, wire_6064, wire_2006, wire_6083, wire_6082, wire_2006, wire_6123, wire_5888, wire_1956, wire_6081, wire_6080, wire_1956, wire_6061, wire_6060, wire_1952, wire_6099, wire_6098, wire_1952, wire_6035, wire_6034, wire_6139, wire_5952, wire_5947, wire_5946, wire_6055, wire_6054, wire_6115, wire_6114, wire_6155, wire_6016, wire_6011, wire_6010, wire_6133, wire_5928, wire_5923, wire_5922, wire_6049, wire_6048, wire_6109, wire_6108, wire_2014, wire_6149, wire_5992, wire_2014, wire_5987, wire_5986, wire_2010, wire_6127, wire_5904, wire_2010, wire_5899, wire_5898, wire_2006, wire_6043, wire_6042, wire_2006, wire_6103, wire_6102, wire_1956, wire_6143, wire_5968, wire_1956, wire_5963, wire_5962, wire_1952, wire_6121, wire_5880, wire_1952};
    // CHNAXY TOTAL: 796
    assign wire_3481 = lut_tile_3_5_chanxy_out[0];
    assign wire_3483 = lut_tile_3_5_chanxy_out[1];
    assign wire_3485 = lut_tile_3_5_chanxy_out[2];
    assign wire_3487 = lut_tile_3_5_chanxy_out[3];
    assign wire_3489 = lut_tile_3_5_chanxy_out[4];
    assign wire_3491 = lut_tile_3_5_chanxy_out[5];
    assign wire_3493 = lut_tile_3_5_chanxy_out[6];
    assign wire_3495 = lut_tile_3_5_chanxy_out[7];
    assign wire_3497 = lut_tile_3_5_chanxy_out[8];
    assign wire_3499 = lut_tile_3_5_chanxy_out[9];
    assign wire_3501 = lut_tile_3_5_chanxy_out[10];
    assign wire_3503 = lut_tile_3_5_chanxy_out[11];
    assign wire_3505 = lut_tile_3_5_chanxy_out[12];
    assign wire_3507 = lut_tile_3_5_chanxy_out[13];
    assign wire_3509 = lut_tile_3_5_chanxy_out[14];
    assign wire_3511 = lut_tile_3_5_chanxy_out[15];
    assign wire_3513 = lut_tile_3_5_chanxy_out[16];
    assign wire_3515 = lut_tile_3_5_chanxy_out[17];
    assign wire_3517 = lut_tile_3_5_chanxy_out[18];
    assign wire_3519 = lut_tile_3_5_chanxy_out[19];
    assign wire_3521 = lut_tile_3_5_chanxy_out[20];
    assign wire_3523 = lut_tile_3_5_chanxy_out[21];
    assign wire_3525 = lut_tile_3_5_chanxy_out[22];
    assign wire_3527 = lut_tile_3_5_chanxy_out[23];
    assign wire_3529 = lut_tile_3_5_chanxy_out[24];
    assign wire_3531 = lut_tile_3_5_chanxy_out[25];
    assign wire_3533 = lut_tile_3_5_chanxy_out[26];
    assign wire_3535 = lut_tile_3_5_chanxy_out[27];
    assign wire_3537 = lut_tile_3_5_chanxy_out[28];
    assign wire_3539 = lut_tile_3_5_chanxy_out[29];
    assign wire_3541 = lut_tile_3_5_chanxy_out[30];
    assign wire_3543 = lut_tile_3_5_chanxy_out[31];
    assign wire_3545 = lut_tile_3_5_chanxy_out[32];
    assign wire_3547 = lut_tile_3_5_chanxy_out[33];
    assign wire_3549 = lut_tile_3_5_chanxy_out[34];
    assign wire_3551 = lut_tile_3_5_chanxy_out[35];
    assign wire_3553 = lut_tile_3_5_chanxy_out[36];
    assign wire_3555 = lut_tile_3_5_chanxy_out[37];
    assign wire_3557 = lut_tile_3_5_chanxy_out[38];
    assign wire_3559 = lut_tile_3_5_chanxy_out[39];
    assign wire_3561 = lut_tile_3_5_chanxy_out[40];
    assign wire_3563 = lut_tile_3_5_chanxy_out[41];
    assign wire_3565 = lut_tile_3_5_chanxy_out[42];
    assign wire_3567 = lut_tile_3_5_chanxy_out[43];
    assign wire_3569 = lut_tile_3_5_chanxy_out[44];
    assign wire_3571 = lut_tile_3_5_chanxy_out[45];
    assign wire_3573 = lut_tile_3_5_chanxy_out[46];
    assign wire_3575 = lut_tile_3_5_chanxy_out[47];
    assign wire_3577 = lut_tile_3_5_chanxy_out[48];
    assign wire_3579 = lut_tile_3_5_chanxy_out[49];
    assign wire_3581 = lut_tile_3_5_chanxy_out[50];
    assign wire_3583 = lut_tile_3_5_chanxy_out[51];
    assign wire_3585 = lut_tile_3_5_chanxy_out[52];
    assign wire_3587 = lut_tile_3_5_chanxy_out[53];
    assign wire_3589 = lut_tile_3_5_chanxy_out[54];
    assign wire_3591 = lut_tile_3_5_chanxy_out[55];
    assign wire_3593 = lut_tile_3_5_chanxy_out[56];
    assign wire_3595 = lut_tile_3_5_chanxy_out[57];
    assign wire_3597 = lut_tile_3_5_chanxy_out[58];
    assign wire_3599 = lut_tile_3_5_chanxy_out[59];
    assign wire_3600 = lut_tile_3_5_chanxy_out[60];
    assign wire_3601 = lut_tile_3_5_chanxy_out[61];
    assign wire_3602 = lut_tile_3_5_chanxy_out[62];
    assign wire_3603 = lut_tile_3_5_chanxy_out[63];
    assign wire_3604 = lut_tile_3_5_chanxy_out[64];
    assign wire_3605 = lut_tile_3_5_chanxy_out[65];
    assign wire_3606 = lut_tile_3_5_chanxy_out[66];
    assign wire_3607 = lut_tile_3_5_chanxy_out[67];
    assign wire_3608 = lut_tile_3_5_chanxy_out[68];
    assign wire_3609 = lut_tile_3_5_chanxy_out[69];
    assign wire_3610 = lut_tile_3_5_chanxy_out[70];
    assign wire_3611 = lut_tile_3_5_chanxy_out[71];
    assign wire_3612 = lut_tile_3_5_chanxy_out[72];
    assign wire_3613 = lut_tile_3_5_chanxy_out[73];
    assign wire_3614 = lut_tile_3_5_chanxy_out[74];
    assign wire_3615 = lut_tile_3_5_chanxy_out[75];
    assign wire_3616 = lut_tile_3_5_chanxy_out[76];
    assign wire_3617 = lut_tile_3_5_chanxy_out[77];
    assign wire_3618 = lut_tile_3_5_chanxy_out[78];
    assign wire_3619 = lut_tile_3_5_chanxy_out[79];
    assign wire_3620 = lut_tile_3_5_chanxy_out[80];
    assign wire_3621 = lut_tile_3_5_chanxy_out[81];
    assign wire_3622 = lut_tile_3_5_chanxy_out[82];
    assign wire_3623 = lut_tile_3_5_chanxy_out[83];
    assign wire_3624 = lut_tile_3_5_chanxy_out[84];
    assign wire_3625 = lut_tile_3_5_chanxy_out[85];
    assign wire_3626 = lut_tile_3_5_chanxy_out[86];
    assign wire_3627 = lut_tile_3_5_chanxy_out[87];
    assign wire_3628 = lut_tile_3_5_chanxy_out[88];
    assign wire_3629 = lut_tile_3_5_chanxy_out[89];
    assign wire_3630 = lut_tile_3_5_chanxy_out[90];
    assign wire_3631 = lut_tile_3_5_chanxy_out[91];
    assign wire_3632 = lut_tile_3_5_chanxy_out[92];
    assign wire_3633 = lut_tile_3_5_chanxy_out[93];
    assign wire_3634 = lut_tile_3_5_chanxy_out[94];
    assign wire_3635 = lut_tile_3_5_chanxy_out[95];
    assign wire_3636 = lut_tile_3_5_chanxy_out[96];
    assign wire_3637 = lut_tile_3_5_chanxy_out[97];
    assign wire_3638 = lut_tile_3_5_chanxy_out[98];
    assign wire_3639 = lut_tile_3_5_chanxy_out[99];
    assign wire_5881 = lut_tile_3_5_chanxy_out[100];
    assign wire_5889 = lut_tile_3_5_chanxy_out[101];
    assign wire_5897 = lut_tile_3_5_chanxy_out[102];
    assign wire_5905 = lut_tile_3_5_chanxy_out[103];
    assign wire_5913 = lut_tile_3_5_chanxy_out[104];
    assign wire_5921 = lut_tile_3_5_chanxy_out[105];
    assign wire_5929 = lut_tile_3_5_chanxy_out[106];
    assign wire_5937 = lut_tile_3_5_chanxy_out[107];
    assign wire_5945 = lut_tile_3_5_chanxy_out[108];
    assign wire_5953 = lut_tile_3_5_chanxy_out[109];
    assign wire_5961 = lut_tile_3_5_chanxy_out[110];
    assign wire_5969 = lut_tile_3_5_chanxy_out[111];
    assign wire_5977 = lut_tile_3_5_chanxy_out[112];
    assign wire_5985 = lut_tile_3_5_chanxy_out[113];
    assign wire_5993 = lut_tile_3_5_chanxy_out[114];
    assign wire_6001 = lut_tile_3_5_chanxy_out[115];
    assign wire_6009 = lut_tile_3_5_chanxy_out[116];
    assign wire_6017 = lut_tile_3_5_chanxy_out[117];
    assign wire_6025 = lut_tile_3_5_chanxy_out[118];
    assign wire_6033 = lut_tile_3_5_chanxy_out[119];
    assign wire_6080 = lut_tile_3_5_chanxy_out[120];
    assign wire_6082 = lut_tile_3_5_chanxy_out[121];
    assign wire_6084 = lut_tile_3_5_chanxy_out[122];
    assign wire_6086 = lut_tile_3_5_chanxy_out[123];
    assign wire_6088 = lut_tile_3_5_chanxy_out[124];
    assign wire_6090 = lut_tile_3_5_chanxy_out[125];
    assign wire_6092 = lut_tile_3_5_chanxy_out[126];
    assign wire_6094 = lut_tile_3_5_chanxy_out[127];
    assign wire_6096 = lut_tile_3_5_chanxy_out[128];
    assign wire_6098 = lut_tile_3_5_chanxy_out[129];
    assign wire_6100 = lut_tile_3_5_chanxy_out[130];
    assign wire_6102 = lut_tile_3_5_chanxy_out[131];
    assign wire_6104 = lut_tile_3_5_chanxy_out[132];
    assign wire_6106 = lut_tile_3_5_chanxy_out[133];
    assign wire_6108 = lut_tile_3_5_chanxy_out[134];
    assign wire_6110 = lut_tile_3_5_chanxy_out[135];
    assign wire_6112 = lut_tile_3_5_chanxy_out[136];
    assign wire_6114 = lut_tile_3_5_chanxy_out[137];
    assign wire_6116 = lut_tile_3_5_chanxy_out[138];
    assign wire_6118 = lut_tile_3_5_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_4_1_chanxy_in = {wire_4752, wire_3481, wire_3479, wire_3478, wire_3427, wire_3426, wire_3373, wire_3372, wire_3328, wire_883, wire_509, wire_4744, wire_3519, wire_3477, wire_3476, wire_3423, wire_3422, wire_3371, wire_3370, wire_3336, wire_883, wire_509, wire_4736, wire_3517, wire_3475, wire_3474, wire_3421, wire_3420, wire_3367, wire_3366, wire_3344, wire_883, wire_509, wire_4728, wire_3515, wire_3471, wire_3470, wire_3419, wire_3418, wire_3365, wire_3364, wire_3352, wire_883, wire_509, wire_4720, wire_3513, wire_3469, wire_3468, wire_3415, wire_3414, wire_3363, wire_3362, wire_3360, wire_883, wire_505, wire_4712, wire_3511, wire_3467, wire_3466, wire_3413, wire_3412, wire_3368, wire_3359, wire_3358, wire_883, wire_505, wire_4704, wire_3509, wire_3463, wire_3462, wire_3411, wire_3410, wire_3376, wire_3357, wire_3356, wire_883, wire_505, wire_4696, wire_3507, wire_3461, wire_3460, wire_3407, wire_3406, wire_3384, wire_3355, wire_3354, wire_883, wire_505, wire_4688, wire_3505, wire_3459, wire_3458, wire_3405, wire_3404, wire_3392, wire_3351, wire_3350, wire_879, wire_505, wire_4680, wire_3503, wire_3455, wire_3454, wire_3403, wire_3402, wire_3400, wire_3349, wire_3348, wire_879, wire_505, wire_4672, wire_3501, wire_3453, wire_3452, wire_3408, wire_3399, wire_3398, wire_3347, wire_3346, wire_879, wire_505, wire_4664, wire_3499, wire_3451, wire_3450, wire_3416, wire_3397, wire_3396, wire_3343, wire_3342, wire_879, wire_505, wire_4656, wire_3497, wire_3447, wire_3446, wire_3424, wire_3395, wire_3394, wire_3341, wire_3340, wire_879, wire_501, wire_4648, wire_3495, wire_3445, wire_3444, wire_3432, wire_3391, wire_3390, wire_3339, wire_3338, wire_879, wire_501, wire_4640, wire_3493, wire_3443, wire_3442, wire_3440, wire_3389, wire_3388, wire_3335, wire_3334, wire_879, wire_501, wire_4632, wire_3491, wire_3448, wire_3439, wire_3438, wire_3387, wire_3386, wire_3333, wire_3332, wire_879, wire_501, wire_4624, wire_3489, wire_3456, wire_3437, wire_3436, wire_3383, wire_3382, wire_3331, wire_3330, wire_509, wire_501, wire_4616, wire_3487, wire_3464, wire_3435, wire_3434, wire_3381, wire_3380, wire_3327, wire_3326, wire_509, wire_501, wire_4608, wire_3485, wire_3472, wire_3431, wire_3430, wire_3379, wire_3378, wire_3325, wire_3324, wire_509, wire_501, wire_4600, wire_3483, wire_3429, wire_3428, wire_3375, wire_3374, wire_3323, wire_3322, wire_3320, wire_509, wire_501, wire_4919, wire_3839, wire_3799, wire_3798, wire_3745, wire_3744, wire_3693, wire_3692, wire_3642, wire_883, wire_509, wire_4917, wire_3801, wire_3797, wire_3796, wire_3794, wire_3743, wire_3742, wire_3689, wire_3688, wire_883, wire_509, wire_4915, wire_3803, wire_3793, wire_3792, wire_3786, wire_3741, wire_3740, wire_3687, wire_3686, wire_883, wire_509, wire_4913, wire_3805, wire_3791, wire_3790, wire_3778, wire_3737, wire_3736, wire_3685, wire_3684, wire_883, wire_509, wire_4911, wire_3807, wire_3789, wire_3788, wire_3770, wire_3735, wire_3734, wire_3681, wire_3680, wire_883, wire_505, wire_4909, wire_3809, wire_3785, wire_3784, wire_3762, wire_3733, wire_3732, wire_3679, wire_3678, wire_883, wire_505, wire_4907, wire_3811, wire_3783, wire_3782, wire_3754, wire_3729, wire_3728, wire_3677, wire_3676, wire_883, wire_505, wire_4905, wire_3813, wire_3781, wire_3780, wire_3746, wire_3727, wire_3726, wire_3673, wire_3672, wire_883, wire_505, wire_4903, wire_3815, wire_3777, wire_3776, wire_3738, wire_3725, wire_3724, wire_3671, wire_3670, wire_879, wire_505, wire_4901, wire_3817, wire_3775, wire_3774, wire_3730, wire_3721, wire_3720, wire_3669, wire_3668, wire_879, wire_505, wire_4899, wire_3819, wire_3773, wire_3772, wire_3722, wire_3719, wire_3718, wire_3665, wire_3664, wire_879, wire_505, wire_4897, wire_3821, wire_3769, wire_3768, wire_3717, wire_3716, wire_3714, wire_3663, wire_3662, wire_879, wire_505, wire_4895, wire_3823, wire_3767, wire_3766, wire_3713, wire_3712, wire_3706, wire_3661, wire_3660, wire_879, wire_501, wire_4893, wire_3825, wire_3765, wire_3764, wire_3711, wire_3710, wire_3698, wire_3657, wire_3656, wire_879, wire_501, wire_4891, wire_3827, wire_3761, wire_3760, wire_3709, wire_3708, wire_3690, wire_3655, wire_3654, wire_879, wire_501, wire_4889, wire_3829, wire_3759, wire_3758, wire_3705, wire_3704, wire_3682, wire_3653, wire_3652, wire_879, wire_501, wire_4887, wire_3831, wire_3757, wire_3756, wire_3703, wire_3702, wire_3674, wire_3649, wire_3648, wire_509, wire_501, wire_4885, wire_3833, wire_3753, wire_3752, wire_3701, wire_3700, wire_3666, wire_3647, wire_3646, wire_509, wire_501, wire_4883, wire_3835, wire_3751, wire_3750, wire_3697, wire_3696, wire_3658, wire_3645, wire_3644, wire_509, wire_501, wire_4881, wire_3837, wire_3749, wire_3748, wire_3695, wire_3694, wire_3650, wire_3641, wire_3640, wire_509, wire_501, wire_4559, wire_4558, wire_4519, wire_4518, wire_4883, wire_4867, wire_4866, wire_4839, wire_4838, wire_4773, wire_4772, wire_4746, wire_3839, wire_566, wire_558, wire_4459, wire_4458, wire_4479, wire_4478, wire_4599, wire_4432, wire_4579, wire_4352, wire_4885, wire_4853, wire_4852, wire_4825, wire_4824, wire_4799, wire_4798, wire_4738, wire_3837, wire_566, wire_558, wire_4557, wire_4556, wire_4517, wire_4516, wire_4477, wire_4476, wire_4537, wire_4536, wire_4887, wire_4879, wire_4878, wire_4811, wire_4810, wire_4785, wire_4784, wire_4730, wire_3835, wire_566, wire_558, wire_4497, wire_4496, wire_4597, wire_4424, wire_4457, wire_4456, wire_4577, wire_4344, wire_4889, wire_4865, wire_4864, wire_4837, wire_4836, wire_4771, wire_4770, wire_4722, wire_3833, wire_566, wire_558, wire_4555, wire_4554, wire_4535, wire_4534, wire_4495, wire_4494, wire_4515, wire_4514, wire_4891, wire_4851, wire_4850, wire_4823, wire_4822, wire_4797, wire_4796, wire_4714, wire_3831, wire_566, wire_508, wire_4455, wire_4454, wire_4575, wire_4336, wire_4533, wire_4532, wire_4475, wire_4474, wire_4893, wire_4877, wire_4876, wire_4809, wire_4808, wire_4783, wire_4782, wire_4706, wire_3829, wire_566, wire_508, wire_4595, wire_4416, wire_4493, wire_4492, wire_4553, wire_4552, wire_4513, wire_4512, wire_4895, wire_4863, wire_4862, wire_4835, wire_4834, wire_4769, wire_4768, wire_4698, wire_3827, wire_566, wire_508, wire_4453, wire_4452, wire_4473, wire_4472, wire_4593, wire_4408, wire_4573, wire_4328, wire_4897, wire_4849, wire_4848, wire_4821, wire_4820, wire_4795, wire_4794, wire_4690, wire_3825, wire_566, wire_508, wire_4551, wire_4550, wire_4511, wire_4510, wire_4471, wire_4470, wire_4531, wire_4530, wire_4899, wire_4875, wire_4874, wire_4807, wire_4806, wire_4781, wire_4780, wire_4682, wire_3823, wire_562, wire_508, wire_4491, wire_4490, wire_4591, wire_4400, wire_4451, wire_4450, wire_4571, wire_4320, wire_4901, wire_4861, wire_4860, wire_4833, wire_4832, wire_4767, wire_4766, wire_4674, wire_3821, wire_562, wire_508, wire_4549, wire_4548, wire_4529, wire_4528, wire_4489, wire_4488, wire_566, wire_4509, wire_4508, wire_566, wire_4903, wire_4847, wire_4846, wire_4819, wire_4818, wire_4793, wire_4792, wire_4666, wire_3819, wire_562, wire_508, wire_4449, wire_4448, wire_566, wire_4569, wire_4312, wire_566, wire_4527, wire_4526, wire_566, wire_4469, wire_4468, wire_566, wire_4905, wire_4873, wire_4872, wire_4805, wire_4804, wire_4779, wire_4778, wire_4658, wire_3817, wire_562, wire_508, wire_4589, wire_4392, wire_566, wire_4487, wire_4486, wire_566, wire_4547, wire_4546, wire_562, wire_4507, wire_4506, wire_562, wire_4907, wire_4859, wire_4858, wire_4831, wire_4830, wire_4765, wire_4764, wire_4650, wire_3815, wire_562, wire_504, wire_4447, wire_4446, wire_562, wire_4467, wire_4466, wire_562, wire_4587, wire_4384, wire_562, wire_4567, wire_4304, wire_562, wire_4909, wire_4845, wire_4844, wire_4817, wire_4816, wire_4791, wire_4790, wire_4642, wire_3813, wire_562, wire_504, wire_4545, wire_4544, wire_562, wire_4505, wire_4504, wire_562, wire_4465, wire_4464, wire_558, wire_4525, wire_4524, wire_558, wire_4911, wire_4871, wire_4870, wire_4803, wire_4802, wire_4777, wire_4776, wire_4634, wire_3811, wire_562, wire_504, wire_4485, wire_4484, wire_558, wire_4585, wire_4376, wire_558, wire_4445, wire_4444, wire_558, wire_4565, wire_4296, wire_558, wire_4913, wire_4857, wire_4856, wire_4829, wire_4828, wire_4763, wire_4762, wire_4626, wire_3809, wire_562, wire_504, wire_4543, wire_4542, wire_558, wire_4523, wire_4522, wire_558, wire_4483, wire_4482, wire_508, wire_4503, wire_4502, wire_508, wire_4915, wire_4843, wire_4842, wire_4815, wire_4814, wire_4789, wire_4788, wire_4618, wire_3807, wire_558, wire_504, wire_4443, wire_4442, wire_508, wire_4563, wire_4288, wire_508, wire_4521, wire_4520, wire_508, wire_4463, wire_4462, wire_508, wire_4917, wire_4869, wire_4868, wire_4801, wire_4800, wire_4775, wire_4774, wire_4610, wire_3805, wire_558, wire_504, wire_4583, wire_4368, wire_508, wire_4481, wire_4480, wire_508, wire_4541, wire_4540, wire_504, wire_4501, wire_4500, wire_504, wire_4919, wire_4855, wire_4854, wire_4827, wire_4826, wire_4761, wire_4760, wire_4602, wire_3803, wire_558, wire_504, wire_4441, wire_4440, wire_504, wire_4461, wire_4460, wire_504, wire_4581, wire_4360, wire_504, wire_4561, wire_4280, wire_504, wire_4881, wire_4841, wire_4840, wire_4813, wire_4812, wire_4787, wire_4786, wire_4754, wire_3801, wire_558, wire_504, wire_4539, wire_4538, wire_504, wire_4499, wire_4498, wire_504};
    // CHNAXY TOTAL: 860
    assign wire_3640 = lut_tile_4_1_chanxy_out[0];
    assign wire_3642 = lut_tile_4_1_chanxy_out[1];
    assign wire_3643 = lut_tile_4_1_chanxy_out[2];
    assign wire_3644 = lut_tile_4_1_chanxy_out[3];
    assign wire_3646 = lut_tile_4_1_chanxy_out[4];
    assign wire_3648 = lut_tile_4_1_chanxy_out[5];
    assign wire_3650 = lut_tile_4_1_chanxy_out[6];
    assign wire_3651 = lut_tile_4_1_chanxy_out[7];
    assign wire_3652 = lut_tile_4_1_chanxy_out[8];
    assign wire_3654 = lut_tile_4_1_chanxy_out[9];
    assign wire_3656 = lut_tile_4_1_chanxy_out[10];
    assign wire_3658 = lut_tile_4_1_chanxy_out[11];
    assign wire_3659 = lut_tile_4_1_chanxy_out[12];
    assign wire_3660 = lut_tile_4_1_chanxy_out[13];
    assign wire_3662 = lut_tile_4_1_chanxy_out[14];
    assign wire_3664 = lut_tile_4_1_chanxy_out[15];
    assign wire_3666 = lut_tile_4_1_chanxy_out[16];
    assign wire_3667 = lut_tile_4_1_chanxy_out[17];
    assign wire_3668 = lut_tile_4_1_chanxy_out[18];
    assign wire_3670 = lut_tile_4_1_chanxy_out[19];
    assign wire_3672 = lut_tile_4_1_chanxy_out[20];
    assign wire_3674 = lut_tile_4_1_chanxy_out[21];
    assign wire_3675 = lut_tile_4_1_chanxy_out[22];
    assign wire_3676 = lut_tile_4_1_chanxy_out[23];
    assign wire_3678 = lut_tile_4_1_chanxy_out[24];
    assign wire_3680 = lut_tile_4_1_chanxy_out[25];
    assign wire_3682 = lut_tile_4_1_chanxy_out[26];
    assign wire_3683 = lut_tile_4_1_chanxy_out[27];
    assign wire_3684 = lut_tile_4_1_chanxy_out[28];
    assign wire_3686 = lut_tile_4_1_chanxy_out[29];
    assign wire_3688 = lut_tile_4_1_chanxy_out[30];
    assign wire_3690 = lut_tile_4_1_chanxy_out[31];
    assign wire_3691 = lut_tile_4_1_chanxy_out[32];
    assign wire_3692 = lut_tile_4_1_chanxy_out[33];
    assign wire_3694 = lut_tile_4_1_chanxy_out[34];
    assign wire_3696 = lut_tile_4_1_chanxy_out[35];
    assign wire_3698 = lut_tile_4_1_chanxy_out[36];
    assign wire_3699 = lut_tile_4_1_chanxy_out[37];
    assign wire_3700 = lut_tile_4_1_chanxy_out[38];
    assign wire_3702 = lut_tile_4_1_chanxy_out[39];
    assign wire_3704 = lut_tile_4_1_chanxy_out[40];
    assign wire_3706 = lut_tile_4_1_chanxy_out[41];
    assign wire_3707 = lut_tile_4_1_chanxy_out[42];
    assign wire_3708 = lut_tile_4_1_chanxy_out[43];
    assign wire_3710 = lut_tile_4_1_chanxy_out[44];
    assign wire_3712 = lut_tile_4_1_chanxy_out[45];
    assign wire_3714 = lut_tile_4_1_chanxy_out[46];
    assign wire_3715 = lut_tile_4_1_chanxy_out[47];
    assign wire_3716 = lut_tile_4_1_chanxy_out[48];
    assign wire_3718 = lut_tile_4_1_chanxy_out[49];
    assign wire_3720 = lut_tile_4_1_chanxy_out[50];
    assign wire_3722 = lut_tile_4_1_chanxy_out[51];
    assign wire_3723 = lut_tile_4_1_chanxy_out[52];
    assign wire_3724 = lut_tile_4_1_chanxy_out[53];
    assign wire_3726 = lut_tile_4_1_chanxy_out[54];
    assign wire_3728 = lut_tile_4_1_chanxy_out[55];
    assign wire_3730 = lut_tile_4_1_chanxy_out[56];
    assign wire_3731 = lut_tile_4_1_chanxy_out[57];
    assign wire_3732 = lut_tile_4_1_chanxy_out[58];
    assign wire_3734 = lut_tile_4_1_chanxy_out[59];
    assign wire_3736 = lut_tile_4_1_chanxy_out[60];
    assign wire_3738 = lut_tile_4_1_chanxy_out[61];
    assign wire_3739 = lut_tile_4_1_chanxy_out[62];
    assign wire_3740 = lut_tile_4_1_chanxy_out[63];
    assign wire_3742 = lut_tile_4_1_chanxy_out[64];
    assign wire_3744 = lut_tile_4_1_chanxy_out[65];
    assign wire_3746 = lut_tile_4_1_chanxy_out[66];
    assign wire_3747 = lut_tile_4_1_chanxy_out[67];
    assign wire_3748 = lut_tile_4_1_chanxy_out[68];
    assign wire_3750 = lut_tile_4_1_chanxy_out[69];
    assign wire_3752 = lut_tile_4_1_chanxy_out[70];
    assign wire_3754 = lut_tile_4_1_chanxy_out[71];
    assign wire_3755 = lut_tile_4_1_chanxy_out[72];
    assign wire_3756 = lut_tile_4_1_chanxy_out[73];
    assign wire_3758 = lut_tile_4_1_chanxy_out[74];
    assign wire_3760 = lut_tile_4_1_chanxy_out[75];
    assign wire_3762 = lut_tile_4_1_chanxy_out[76];
    assign wire_3763 = lut_tile_4_1_chanxy_out[77];
    assign wire_3764 = lut_tile_4_1_chanxy_out[78];
    assign wire_3766 = lut_tile_4_1_chanxy_out[79];
    assign wire_3768 = lut_tile_4_1_chanxy_out[80];
    assign wire_3770 = lut_tile_4_1_chanxy_out[81];
    assign wire_3771 = lut_tile_4_1_chanxy_out[82];
    assign wire_3772 = lut_tile_4_1_chanxy_out[83];
    assign wire_3774 = lut_tile_4_1_chanxy_out[84];
    assign wire_3776 = lut_tile_4_1_chanxy_out[85];
    assign wire_3778 = lut_tile_4_1_chanxy_out[86];
    assign wire_3779 = lut_tile_4_1_chanxy_out[87];
    assign wire_3780 = lut_tile_4_1_chanxy_out[88];
    assign wire_3782 = lut_tile_4_1_chanxy_out[89];
    assign wire_3784 = lut_tile_4_1_chanxy_out[90];
    assign wire_3786 = lut_tile_4_1_chanxy_out[91];
    assign wire_3787 = lut_tile_4_1_chanxy_out[92];
    assign wire_3788 = lut_tile_4_1_chanxy_out[93];
    assign wire_3790 = lut_tile_4_1_chanxy_out[94];
    assign wire_3792 = lut_tile_4_1_chanxy_out[95];
    assign wire_3794 = lut_tile_4_1_chanxy_out[96];
    assign wire_3795 = lut_tile_4_1_chanxy_out[97];
    assign wire_3796 = lut_tile_4_1_chanxy_out[98];
    assign wire_3798 = lut_tile_4_1_chanxy_out[99];
    assign wire_4603 = lut_tile_4_1_chanxy_out[100];
    assign wire_4611 = lut_tile_4_1_chanxy_out[101];
    assign wire_4619 = lut_tile_4_1_chanxy_out[102];
    assign wire_4627 = lut_tile_4_1_chanxy_out[103];
    assign wire_4635 = lut_tile_4_1_chanxy_out[104];
    assign wire_4643 = lut_tile_4_1_chanxy_out[105];
    assign wire_4651 = lut_tile_4_1_chanxy_out[106];
    assign wire_4659 = lut_tile_4_1_chanxy_out[107];
    assign wire_4667 = lut_tile_4_1_chanxy_out[108];
    assign wire_4675 = lut_tile_4_1_chanxy_out[109];
    assign wire_4683 = lut_tile_4_1_chanxy_out[110];
    assign wire_4691 = lut_tile_4_1_chanxy_out[111];
    assign wire_4699 = lut_tile_4_1_chanxy_out[112];
    assign wire_4707 = lut_tile_4_1_chanxy_out[113];
    assign wire_4715 = lut_tile_4_1_chanxy_out[114];
    assign wire_4723 = lut_tile_4_1_chanxy_out[115];
    assign wire_4731 = lut_tile_4_1_chanxy_out[116];
    assign wire_4739 = lut_tile_4_1_chanxy_out[117];
    assign wire_4747 = lut_tile_4_1_chanxy_out[118];
    assign wire_4755 = lut_tile_4_1_chanxy_out[119];
    assign wire_4840 = lut_tile_4_1_chanxy_out[120];
    assign wire_4842 = lut_tile_4_1_chanxy_out[121];
    assign wire_4844 = lut_tile_4_1_chanxy_out[122];
    assign wire_4846 = lut_tile_4_1_chanxy_out[123];
    assign wire_4848 = lut_tile_4_1_chanxy_out[124];
    assign wire_4850 = lut_tile_4_1_chanxy_out[125];
    assign wire_4852 = lut_tile_4_1_chanxy_out[126];
    assign wire_4854 = lut_tile_4_1_chanxy_out[127];
    assign wire_4856 = lut_tile_4_1_chanxy_out[128];
    assign wire_4858 = lut_tile_4_1_chanxy_out[129];
    assign wire_4860 = lut_tile_4_1_chanxy_out[130];
    assign wire_4862 = lut_tile_4_1_chanxy_out[131];
    assign wire_4864 = lut_tile_4_1_chanxy_out[132];
    assign wire_4866 = lut_tile_4_1_chanxy_out[133];
    assign wire_4868 = lut_tile_4_1_chanxy_out[134];
    assign wire_4870 = lut_tile_4_1_chanxy_out[135];
    assign wire_4872 = lut_tile_4_1_chanxy_out[136];
    assign wire_4874 = lut_tile_4_1_chanxy_out[137];
    assign wire_4876 = lut_tile_4_1_chanxy_out[138];
    assign wire_4878 = lut_tile_4_1_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_4_2_chanxy_in = {wire_5074, wire_3521, wire_3507, wire_3506, wire_3479, wire_3478, wire_3373, wire_3372, wire_3330, wire_1259, wire_885, wire_5066, wire_3559, wire_3493, wire_3492, wire_3477, wire_3476, wire_3423, wire_3422, wire_3338, wire_1259, wire_885, wire_5058, wire_3557, wire_3519, wire_3518, wire_3421, wire_3420, wire_3367, wire_3366, wire_3346, wire_1259, wire_885, wire_5050, wire_3555, wire_3505, wire_3504, wire_3471, wire_3470, wire_3365, wire_3364, wire_3354, wire_1259, wire_885, wire_5042, wire_3553, wire_3491, wire_3490, wire_3469, wire_3468, wire_3415, wire_3414, wire_3362, wire_1259, wire_881, wire_5034, wire_3551, wire_3517, wire_3516, wire_3413, wire_3412, wire_3370, wire_3359, wire_3358, wire_1259, wire_881, wire_5026, wire_3549, wire_3503, wire_3502, wire_3463, wire_3462, wire_3378, wire_3357, wire_3356, wire_1259, wire_881, wire_5018, wire_3547, wire_3489, wire_3488, wire_3461, wire_3460, wire_3407, wire_3406, wire_3386, wire_1259, wire_881, wire_5010, wire_3545, wire_3515, wire_3514, wire_3405, wire_3404, wire_3394, wire_3351, wire_3350, wire_1255, wire_881, wire_5002, wire_3543, wire_3501, wire_3500, wire_3455, wire_3454, wire_3402, wire_3349, wire_3348, wire_1255, wire_881, wire_4994, wire_3541, wire_3487, wire_3486, wire_3453, wire_3452, wire_3410, wire_3399, wire_3398, wire_1255, wire_881, wire_4986, wire_3539, wire_3513, wire_3512, wire_3418, wire_3397, wire_3396, wire_3343, wire_3342, wire_1255, wire_881, wire_4978, wire_3537, wire_3499, wire_3498, wire_3447, wire_3446, wire_3426, wire_3341, wire_3340, wire_1255, wire_877, wire_4970, wire_3535, wire_3485, wire_3484, wire_3445, wire_3444, wire_3434, wire_3391, wire_3390, wire_1255, wire_877, wire_4962, wire_3533, wire_3511, wire_3510, wire_3442, wire_3389, wire_3388, wire_3335, wire_3334, wire_1255, wire_877, wire_4954, wire_3531, wire_3497, wire_3496, wire_3450, wire_3439, wire_3438, wire_3333, wire_3332, wire_1255, wire_877, wire_4946, wire_3529, wire_3483, wire_3482, wire_3458, wire_3437, wire_3436, wire_3383, wire_3382, wire_885, wire_877, wire_4938, wire_3527, wire_3509, wire_3508, wire_3466, wire_3381, wire_3380, wire_3327, wire_3326, wire_885, wire_877, wire_4930, wire_3525, wire_3495, wire_3494, wire_3474, wire_3431, wire_3430, wire_3325, wire_3324, wire_885, wire_877, wire_4922, wire_3523, wire_3481, wire_3480, wire_3429, wire_3428, wire_3375, wire_3374, wire_3322, wire_885, wire_877, wire_5239, wire_3879, wire_3813, wire_3812, wire_3799, wire_3798, wire_3745, wire_3744, wire_3644, wire_1259, wire_885, wire_5237, wire_3841, wire_3839, wire_3838, wire_3796, wire_3743, wire_3742, wire_3689, wire_3688, wire_1259, wire_885, wire_5235, wire_3843, wire_3825, wire_3824, wire_3793, wire_3792, wire_3788, wire_3687, wire_3686, wire_1259, wire_885, wire_5233, wire_3845, wire_3811, wire_3810, wire_3791, wire_3790, wire_3780, wire_3737, wire_3736, wire_1259, wire_885, wire_5231, wire_3847, wire_3837, wire_3836, wire_3772, wire_3735, wire_3734, wire_3681, wire_3680, wire_1259, wire_881, wire_5229, wire_3849, wire_3823, wire_3822, wire_3785, wire_3784, wire_3764, wire_3679, wire_3678, wire_1259, wire_881, wire_5227, wire_3851, wire_3809, wire_3808, wire_3783, wire_3782, wire_3756, wire_3729, wire_3728, wire_1259, wire_881, wire_5225, wire_3853, wire_3835, wire_3834, wire_3748, wire_3727, wire_3726, wire_3673, wire_3672, wire_1259, wire_881, wire_5223, wire_3855, wire_3821, wire_3820, wire_3777, wire_3776, wire_3740, wire_3671, wire_3670, wire_1255, wire_881, wire_5221, wire_3857, wire_3807, wire_3806, wire_3775, wire_3774, wire_3732, wire_3721, wire_3720, wire_1255, wire_881, wire_5219, wire_3859, wire_3833, wire_3832, wire_3724, wire_3719, wire_3718, wire_3665, wire_3664, wire_1255, wire_881, wire_5217, wire_3861, wire_3819, wire_3818, wire_3769, wire_3768, wire_3716, wire_3663, wire_3662, wire_1255, wire_881, wire_5215, wire_3863, wire_3805, wire_3804, wire_3767, wire_3766, wire_3713, wire_3712, wire_3708, wire_1255, wire_877, wire_5213, wire_3865, wire_3831, wire_3830, wire_3711, wire_3710, wire_3700, wire_3657, wire_3656, wire_1255, wire_877, wire_5211, wire_3867, wire_3817, wire_3816, wire_3761, wire_3760, wire_3692, wire_3655, wire_3654, wire_1255, wire_877, wire_5209, wire_3869, wire_3803, wire_3802, wire_3759, wire_3758, wire_3705, wire_3704, wire_3684, wire_1255, wire_877, wire_5207, wire_3871, wire_3829, wire_3828, wire_3703, wire_3702, wire_3676, wire_3649, wire_3648, wire_885, wire_877, wire_5205, wire_3873, wire_3815, wire_3814, wire_3753, wire_3752, wire_3668, wire_3647, wire_3646, wire_885, wire_877, wire_5203, wire_3875, wire_3801, wire_3800, wire_3751, wire_3750, wire_3697, wire_3696, wire_3660, wire_885, wire_877, wire_5201, wire_3877, wire_3827, wire_3826, wire_3695, wire_3694, wire_3652, wire_3641, wire_3640, wire_885, wire_877, wire_4917, wire_4867, wire_4866, wire_4839, wire_4838, wire_4773, wire_4772, wire_4754, wire_3794, wire_942, wire_934, wire_4915, wire_4853, wire_4852, wire_4825, wire_4824, wire_4799, wire_4798, wire_4602, wire_3786, wire_942, wire_934, wire_4913, wire_4879, wire_4878, wire_4811, wire_4810, wire_4785, wire_4784, wire_4610, wire_3778, wire_942, wire_934, wire_4911, wire_4865, wire_4864, wire_4837, wire_4836, wire_4771, wire_4770, wire_4618, wire_3770, wire_942, wire_934, wire_4909, wire_4851, wire_4850, wire_4823, wire_4822, wire_4797, wire_4796, wire_4626, wire_3762, wire_942, wire_884, wire_4907, wire_4877, wire_4876, wire_4809, wire_4808, wire_4783, wire_4782, wire_4634, wire_3754, wire_942, wire_884, wire_4905, wire_4863, wire_4862, wire_4835, wire_4834, wire_4769, wire_4768, wire_4642, wire_3746, wire_942, wire_884, wire_4903, wire_4849, wire_4848, wire_4821, wire_4820, wire_4795, wire_4794, wire_4650, wire_3738, wire_942, wire_884, wire_4901, wire_4875, wire_4874, wire_4807, wire_4806, wire_4781, wire_4780, wire_4658, wire_3730, wire_938, wire_884, wire_4899, wire_4861, wire_4860, wire_4833, wire_4832, wire_4767, wire_4766, wire_4666, wire_3722, wire_938, wire_884, wire_4897, wire_4847, wire_4846, wire_4819, wire_4818, wire_4793, wire_4792, wire_4674, wire_3714, wire_938, wire_884, wire_4895, wire_4873, wire_4872, wire_4805, wire_4804, wire_4779, wire_4778, wire_4682, wire_3706, wire_938, wire_884, wire_4893, wire_4859, wire_4858, wire_4831, wire_4830, wire_4765, wire_4764, wire_4690, wire_3698, wire_938, wire_880, wire_4891, wire_4845, wire_4844, wire_4817, wire_4816, wire_4791, wire_4790, wire_4698, wire_3690, wire_938, wire_880, wire_4889, wire_4871, wire_4870, wire_4803, wire_4802, wire_4777, wire_4776, wire_4706, wire_3682, wire_938, wire_880, wire_4887, wire_4857, wire_4856, wire_4829, wire_4828, wire_4763, wire_4762, wire_4714, wire_3674, wire_938, wire_880, wire_4885, wire_4843, wire_4842, wire_4815, wire_4814, wire_4789, wire_4788, wire_4722, wire_3666, wire_934, wire_880, wire_4883, wire_4869, wire_4868, wire_4801, wire_4800, wire_4775, wire_4774, wire_4730, wire_3658, wire_934, wire_880, wire_4881, wire_4855, wire_4854, wire_4827, wire_4826, wire_4761, wire_4760, wire_4738, wire_3650, wire_934, wire_880, wire_4919, wire_4841, wire_4840, wire_4813, wire_4812, wire_4787, wire_4786, wire_4746, wire_3642, wire_934, wire_880, wire_5203, wire_5173, wire_5172, wire_5147, wire_5146, wire_5119, wire_5118, wire_5068, wire_3879, wire_942, wire_934, wire_5205, wire_5199, wire_5198, wire_5133, wire_5132, wire_5105, wire_5104, wire_5060, wire_3877, wire_942, wire_934, wire_5207, wire_5185, wire_5184, wire_5159, wire_5158, wire_5091, wire_5090, wire_5052, wire_3875, wire_942, wire_934, wire_5209, wire_5171, wire_5170, wire_5145, wire_5144, wire_5117, wire_5116, wire_5044, wire_3873, wire_942, wire_934, wire_5211, wire_5197, wire_5196, wire_5131, wire_5130, wire_5103, wire_5102, wire_5036, wire_3871, wire_942, wire_884, wire_5213, wire_5183, wire_5182, wire_5157, wire_5156, wire_5089, wire_5088, wire_5028, wire_3869, wire_942, wire_884, wire_5215, wire_5169, wire_5168, wire_5143, wire_5142, wire_5115, wire_5114, wire_5020, wire_3867, wire_942, wire_884, wire_5217, wire_5195, wire_5194, wire_5129, wire_5128, wire_5101, wire_5100, wire_5012, wire_3865, wire_942, wire_884, wire_5219, wire_5181, wire_5180, wire_5155, wire_5154, wire_5087, wire_5086, wire_5004, wire_3863, wire_938, wire_884, wire_5221, wire_5167, wire_5166, wire_5141, wire_5140, wire_5113, wire_5112, wire_4996, wire_3861, wire_938, wire_884, wire_5223, wire_5193, wire_5192, wire_5127, wire_5126, wire_5099, wire_5098, wire_4988, wire_3859, wire_938, wire_884, wire_5225, wire_5179, wire_5178, wire_5153, wire_5152, wire_5085, wire_5084, wire_4980, wire_3857, wire_938, wire_884, wire_5227, wire_5165, wire_5164, wire_5139, wire_5138, wire_5111, wire_5110, wire_4972, wire_3855, wire_938, wire_880, wire_5229, wire_5191, wire_5190, wire_5125, wire_5124, wire_5097, wire_5096, wire_4964, wire_3853, wire_938, wire_880, wire_5231, wire_5177, wire_5176, wire_5151, wire_5150, wire_5083, wire_5082, wire_4956, wire_3851, wire_938, wire_880, wire_5233, wire_5163, wire_5162, wire_5137, wire_5136, wire_5109, wire_5108, wire_4948, wire_3849, wire_938, wire_880, wire_5235, wire_5189, wire_5188, wire_5123, wire_5122, wire_5095, wire_5094, wire_4940, wire_3847, wire_934, wire_880, wire_5237, wire_5175, wire_5174, wire_5149, wire_5148, wire_5081, wire_5080, wire_4932, wire_3845, wire_934, wire_880, wire_5239, wire_5161, wire_5160, wire_5135, wire_5134, wire_5107, wire_5106, wire_4924, wire_3843, wire_934, wire_880, wire_5201, wire_5187, wire_5186, wire_5121, wire_5120, wire_5093, wire_5092, wire_5076, wire_3841, wire_934, wire_880};
    // CHNAXY TOTAL: 880
    assign wire_3645 = lut_tile_4_2_chanxy_out[0];
    assign wire_3653 = lut_tile_4_2_chanxy_out[1];
    assign wire_3661 = lut_tile_4_2_chanxy_out[2];
    assign wire_3669 = lut_tile_4_2_chanxy_out[3];
    assign wire_3677 = lut_tile_4_2_chanxy_out[4];
    assign wire_3685 = lut_tile_4_2_chanxy_out[5];
    assign wire_3693 = lut_tile_4_2_chanxy_out[6];
    assign wire_3701 = lut_tile_4_2_chanxy_out[7];
    assign wire_3709 = lut_tile_4_2_chanxy_out[8];
    assign wire_3717 = lut_tile_4_2_chanxy_out[9];
    assign wire_3725 = lut_tile_4_2_chanxy_out[10];
    assign wire_3733 = lut_tile_4_2_chanxy_out[11];
    assign wire_3741 = lut_tile_4_2_chanxy_out[12];
    assign wire_3749 = lut_tile_4_2_chanxy_out[13];
    assign wire_3757 = lut_tile_4_2_chanxy_out[14];
    assign wire_3765 = lut_tile_4_2_chanxy_out[15];
    assign wire_3773 = lut_tile_4_2_chanxy_out[16];
    assign wire_3781 = lut_tile_4_2_chanxy_out[17];
    assign wire_3789 = lut_tile_4_2_chanxy_out[18];
    assign wire_3797 = lut_tile_4_2_chanxy_out[19];
    assign wire_3800 = lut_tile_4_2_chanxy_out[20];
    assign wire_3802 = lut_tile_4_2_chanxy_out[21];
    assign wire_3804 = lut_tile_4_2_chanxy_out[22];
    assign wire_3806 = lut_tile_4_2_chanxy_out[23];
    assign wire_3808 = lut_tile_4_2_chanxy_out[24];
    assign wire_3810 = lut_tile_4_2_chanxy_out[25];
    assign wire_3812 = lut_tile_4_2_chanxy_out[26];
    assign wire_3814 = lut_tile_4_2_chanxy_out[27];
    assign wire_3816 = lut_tile_4_2_chanxy_out[28];
    assign wire_3818 = lut_tile_4_2_chanxy_out[29];
    assign wire_3820 = lut_tile_4_2_chanxy_out[30];
    assign wire_3822 = lut_tile_4_2_chanxy_out[31];
    assign wire_3824 = lut_tile_4_2_chanxy_out[32];
    assign wire_3826 = lut_tile_4_2_chanxy_out[33];
    assign wire_3828 = lut_tile_4_2_chanxy_out[34];
    assign wire_3830 = lut_tile_4_2_chanxy_out[35];
    assign wire_3832 = lut_tile_4_2_chanxy_out[36];
    assign wire_3834 = lut_tile_4_2_chanxy_out[37];
    assign wire_3836 = lut_tile_4_2_chanxy_out[38];
    assign wire_3838 = lut_tile_4_2_chanxy_out[39];
    assign wire_4925 = lut_tile_4_2_chanxy_out[40];
    assign wire_4933 = lut_tile_4_2_chanxy_out[41];
    assign wire_4941 = lut_tile_4_2_chanxy_out[42];
    assign wire_4949 = lut_tile_4_2_chanxy_out[43];
    assign wire_4957 = lut_tile_4_2_chanxy_out[44];
    assign wire_4965 = lut_tile_4_2_chanxy_out[45];
    assign wire_4973 = lut_tile_4_2_chanxy_out[46];
    assign wire_4981 = lut_tile_4_2_chanxy_out[47];
    assign wire_4989 = lut_tile_4_2_chanxy_out[48];
    assign wire_4997 = lut_tile_4_2_chanxy_out[49];
    assign wire_5005 = lut_tile_4_2_chanxy_out[50];
    assign wire_5013 = lut_tile_4_2_chanxy_out[51];
    assign wire_5021 = lut_tile_4_2_chanxy_out[52];
    assign wire_5029 = lut_tile_4_2_chanxy_out[53];
    assign wire_5037 = lut_tile_4_2_chanxy_out[54];
    assign wire_5045 = lut_tile_4_2_chanxy_out[55];
    assign wire_5053 = lut_tile_4_2_chanxy_out[56];
    assign wire_5061 = lut_tile_4_2_chanxy_out[57];
    assign wire_5069 = lut_tile_4_2_chanxy_out[58];
    assign wire_5077 = lut_tile_4_2_chanxy_out[59];
    assign wire_5160 = lut_tile_4_2_chanxy_out[60];
    assign wire_5162 = lut_tile_4_2_chanxy_out[61];
    assign wire_5164 = lut_tile_4_2_chanxy_out[62];
    assign wire_5166 = lut_tile_4_2_chanxy_out[63];
    assign wire_5168 = lut_tile_4_2_chanxy_out[64];
    assign wire_5170 = lut_tile_4_2_chanxy_out[65];
    assign wire_5172 = lut_tile_4_2_chanxy_out[66];
    assign wire_5174 = lut_tile_4_2_chanxy_out[67];
    assign wire_5176 = lut_tile_4_2_chanxy_out[68];
    assign wire_5178 = lut_tile_4_2_chanxy_out[69];
    assign wire_5180 = lut_tile_4_2_chanxy_out[70];
    assign wire_5182 = lut_tile_4_2_chanxy_out[71];
    assign wire_5184 = lut_tile_4_2_chanxy_out[72];
    assign wire_5186 = lut_tile_4_2_chanxy_out[73];
    assign wire_5188 = lut_tile_4_2_chanxy_out[74];
    assign wire_5190 = lut_tile_4_2_chanxy_out[75];
    assign wire_5192 = lut_tile_4_2_chanxy_out[76];
    assign wire_5194 = lut_tile_4_2_chanxy_out[77];
    assign wire_5196 = lut_tile_4_2_chanxy_out[78];
    assign wire_5198 = lut_tile_4_2_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_4_3_chanxy_in = {wire_5396, wire_3561, wire_3533, wire_3532, wire_3507, wire_3506, wire_3479, wire_3478, wire_3332, wire_1635, wire_1261, wire_5388, wire_3599, wire_3559, wire_3558, wire_3493, wire_3492, wire_3423, wire_3422, wire_3340, wire_1635, wire_1261, wire_5380, wire_3597, wire_3545, wire_3544, wire_3519, wire_3518, wire_3367, wire_3366, wire_3348, wire_1635, wire_1261, wire_5372, wire_3595, wire_3531, wire_3530, wire_3505, wire_3504, wire_3471, wire_3470, wire_3356, wire_1635, wire_1261, wire_5364, wire_3593, wire_3557, wire_3556, wire_3491, wire_3490, wire_3415, wire_3414, wire_3364, wire_1635, wire_1257, wire_5356, wire_3591, wire_3543, wire_3542, wire_3517, wire_3516, wire_3372, wire_3359, wire_3358, wire_1635, wire_1257, wire_5348, wire_3589, wire_3529, wire_3528, wire_3503, wire_3502, wire_3463, wire_3462, wire_3380, wire_1635, wire_1257, wire_5340, wire_3587, wire_3555, wire_3554, wire_3489, wire_3488, wire_3407, wire_3406, wire_3388, wire_1635, wire_1257, wire_5332, wire_3585, wire_3541, wire_3540, wire_3515, wire_3514, wire_3396, wire_3351, wire_3350, wire_1631, wire_1257, wire_5324, wire_3583, wire_3527, wire_3526, wire_3501, wire_3500, wire_3455, wire_3454, wire_3404, wire_1631, wire_1257, wire_5316, wire_3581, wire_3553, wire_3552, wire_3487, wire_3486, wire_3412, wire_3399, wire_3398, wire_1631, wire_1257, wire_5308, wire_3579, wire_3539, wire_3538, wire_3513, wire_3512, wire_3420, wire_3343, wire_3342, wire_1631, wire_1257, wire_5300, wire_3577, wire_3525, wire_3524, wire_3499, wire_3498, wire_3447, wire_3446, wire_3428, wire_1631, wire_1253, wire_5292, wire_3575, wire_3551, wire_3550, wire_3485, wire_3484, wire_3436, wire_3391, wire_3390, wire_1631, wire_1253, wire_5284, wire_3573, wire_3537, wire_3536, wire_3511, wire_3510, wire_3444, wire_3335, wire_3334, wire_1631, wire_1253, wire_5276, wire_3571, wire_3523, wire_3522, wire_3497, wire_3496, wire_3452, wire_3439, wire_3438, wire_1631, wire_1253, wire_5268, wire_3569, wire_3549, wire_3548, wire_3483, wire_3482, wire_3460, wire_3383, wire_3382, wire_1261, wire_1253, wire_5260, wire_3567, wire_3535, wire_3534, wire_3509, wire_3508, wire_3468, wire_3327, wire_3326, wire_1261, wire_1253, wire_5252, wire_3565, wire_3521, wire_3520, wire_3495, wire_3494, wire_3476, wire_3431, wire_3430, wire_1261, wire_1253, wire_5244, wire_3563, wire_3547, wire_3546, wire_3481, wire_3480, wire_3375, wire_3374, wire_3324, wire_1261, wire_1253, wire_5559, wire_3919, wire_3879, wire_3878, wire_3813, wire_3812, wire_3745, wire_3744, wire_3646, wire_1635, wire_1261, wire_5557, wire_3881, wire_3865, wire_3864, wire_3839, wire_3838, wire_3798, wire_3689, wire_3688, wire_1635, wire_1261, wire_5555, wire_3883, wire_3851, wire_3850, wire_3825, wire_3824, wire_3793, wire_3792, wire_3790, wire_1635, wire_1261, wire_5553, wire_3885, wire_3877, wire_3876, wire_3811, wire_3810, wire_3782, wire_3737, wire_3736, wire_1635, wire_1261, wire_5551, wire_3887, wire_3863, wire_3862, wire_3837, wire_3836, wire_3774, wire_3681, wire_3680, wire_1635, wire_1257, wire_5549, wire_3889, wire_3849, wire_3848, wire_3823, wire_3822, wire_3785, wire_3784, wire_3766, wire_1635, wire_1257, wire_5547, wire_3891, wire_3875, wire_3874, wire_3809, wire_3808, wire_3758, wire_3729, wire_3728, wire_1635, wire_1257, wire_5545, wire_3893, wire_3861, wire_3860, wire_3835, wire_3834, wire_3750, wire_3673, wire_3672, wire_1635, wire_1257, wire_5543, wire_3895, wire_3847, wire_3846, wire_3821, wire_3820, wire_3777, wire_3776, wire_3742, wire_1631, wire_1257, wire_5541, wire_3897, wire_3873, wire_3872, wire_3807, wire_3806, wire_3734, wire_3721, wire_3720, wire_1631, wire_1257, wire_5539, wire_3899, wire_3859, wire_3858, wire_3833, wire_3832, wire_3726, wire_3665, wire_3664, wire_1631, wire_1257, wire_5537, wire_3901, wire_3845, wire_3844, wire_3819, wire_3818, wire_3769, wire_3768, wire_3718, wire_1631, wire_1257, wire_5535, wire_3903, wire_3871, wire_3870, wire_3805, wire_3804, wire_3713, wire_3712, wire_3710, wire_1631, wire_1253, wire_5533, wire_3905, wire_3857, wire_3856, wire_3831, wire_3830, wire_3702, wire_3657, wire_3656, wire_1631, wire_1253, wire_5531, wire_3907, wire_3843, wire_3842, wire_3817, wire_3816, wire_3761, wire_3760, wire_3694, wire_1631, wire_1253, wire_5529, wire_3909, wire_3869, wire_3868, wire_3803, wire_3802, wire_3705, wire_3704, wire_3686, wire_1631, wire_1253, wire_5527, wire_3911, wire_3855, wire_3854, wire_3829, wire_3828, wire_3678, wire_3649, wire_3648, wire_1261, wire_1253, wire_5525, wire_3913, wire_3841, wire_3840, wire_3815, wire_3814, wire_3753, wire_3752, wire_3670, wire_1261, wire_1253, wire_5523, wire_3915, wire_3867, wire_3866, wire_3801, wire_3800, wire_3697, wire_3696, wire_3662, wire_1261, wire_1253, wire_5521, wire_3917, wire_3853, wire_3852, wire_3827, wire_3826, wire_3654, wire_3641, wire_3640, wire_1261, wire_1253, wire_5237, wire_5173, wire_5172, wire_5147, wire_5146, wire_5119, wire_5118, wire_5076, wire_3796, wire_1318, wire_1310, wire_5235, wire_5199, wire_5198, wire_5133, wire_5132, wire_5105, wire_5104, wire_4924, wire_3788, wire_1318, wire_1310, wire_5233, wire_5185, wire_5184, wire_5159, wire_5158, wire_5091, wire_5090, wire_4932, wire_3780, wire_1318, wire_1310, wire_5231, wire_5171, wire_5170, wire_5145, wire_5144, wire_5117, wire_5116, wire_4940, wire_3772, wire_1318, wire_1310, wire_5229, wire_5197, wire_5196, wire_5131, wire_5130, wire_5103, wire_5102, wire_4948, wire_3764, wire_1318, wire_1260, wire_5227, wire_5183, wire_5182, wire_5157, wire_5156, wire_5089, wire_5088, wire_4956, wire_3756, wire_1318, wire_1260, wire_5225, wire_5169, wire_5168, wire_5143, wire_5142, wire_5115, wire_5114, wire_4964, wire_3748, wire_1318, wire_1260, wire_5223, wire_5195, wire_5194, wire_5129, wire_5128, wire_5101, wire_5100, wire_4972, wire_3740, wire_1318, wire_1260, wire_5221, wire_5181, wire_5180, wire_5155, wire_5154, wire_5087, wire_5086, wire_4980, wire_3732, wire_1314, wire_1260, wire_5219, wire_5167, wire_5166, wire_5141, wire_5140, wire_5113, wire_5112, wire_4988, wire_3724, wire_1314, wire_1260, wire_5217, wire_5193, wire_5192, wire_5127, wire_5126, wire_5099, wire_5098, wire_4996, wire_3716, wire_1314, wire_1260, wire_5215, wire_5179, wire_5178, wire_5153, wire_5152, wire_5085, wire_5084, wire_5004, wire_3708, wire_1314, wire_1260, wire_5213, wire_5165, wire_5164, wire_5139, wire_5138, wire_5111, wire_5110, wire_5012, wire_3700, wire_1314, wire_1256, wire_5211, wire_5191, wire_5190, wire_5125, wire_5124, wire_5097, wire_5096, wire_5020, wire_3692, wire_1314, wire_1256, wire_5209, wire_5177, wire_5176, wire_5151, wire_5150, wire_5083, wire_5082, wire_5028, wire_3684, wire_1314, wire_1256, wire_5207, wire_5163, wire_5162, wire_5137, wire_5136, wire_5109, wire_5108, wire_5036, wire_3676, wire_1314, wire_1256, wire_5205, wire_5189, wire_5188, wire_5123, wire_5122, wire_5095, wire_5094, wire_5044, wire_3668, wire_1310, wire_1256, wire_5203, wire_5175, wire_5174, wire_5149, wire_5148, wire_5081, wire_5080, wire_5052, wire_3660, wire_1310, wire_1256, wire_5201, wire_5161, wire_5160, wire_5135, wire_5134, wire_5107, wire_5106, wire_5060, wire_3652, wire_1310, wire_1256, wire_5239, wire_5187, wire_5186, wire_5121, wire_5120, wire_5093, wire_5092, wire_5068, wire_3644, wire_1310, wire_1256, wire_5523, wire_5519, wire_5518, wire_5453, wire_5452, wire_5427, wire_5426, wire_5390, wire_3919, wire_1318, wire_1310, wire_5525, wire_5505, wire_5504, wire_5479, wire_5478, wire_5413, wire_5412, wire_5382, wire_3917, wire_1318, wire_1310, wire_5527, wire_5491, wire_5490, wire_5465, wire_5464, wire_5439, wire_5438, wire_5374, wire_3915, wire_1318, wire_1310, wire_5529, wire_5517, wire_5516, wire_5451, wire_5450, wire_5425, wire_5424, wire_5366, wire_3913, wire_1318, wire_1310, wire_5531, wire_5503, wire_5502, wire_5477, wire_5476, wire_5411, wire_5410, wire_5358, wire_3911, wire_1318, wire_1260, wire_5533, wire_5489, wire_5488, wire_5463, wire_5462, wire_5437, wire_5436, wire_5350, wire_3909, wire_1318, wire_1260, wire_5535, wire_5515, wire_5514, wire_5449, wire_5448, wire_5423, wire_5422, wire_5342, wire_3907, wire_1318, wire_1260, wire_5537, wire_5501, wire_5500, wire_5475, wire_5474, wire_5409, wire_5408, wire_5334, wire_3905, wire_1318, wire_1260, wire_5539, wire_5487, wire_5486, wire_5461, wire_5460, wire_5435, wire_5434, wire_5326, wire_3903, wire_1314, wire_1260, wire_5541, wire_5513, wire_5512, wire_5447, wire_5446, wire_5421, wire_5420, wire_5318, wire_3901, wire_1314, wire_1260, wire_5543, wire_5499, wire_5498, wire_5473, wire_5472, wire_5407, wire_5406, wire_5310, wire_3899, wire_1314, wire_1260, wire_5545, wire_5485, wire_5484, wire_5459, wire_5458, wire_5433, wire_5432, wire_5302, wire_3897, wire_1314, wire_1260, wire_5547, wire_5511, wire_5510, wire_5445, wire_5444, wire_5419, wire_5418, wire_5294, wire_3895, wire_1314, wire_1256, wire_5549, wire_5497, wire_5496, wire_5471, wire_5470, wire_5405, wire_5404, wire_5286, wire_3893, wire_1314, wire_1256, wire_5551, wire_5483, wire_5482, wire_5457, wire_5456, wire_5431, wire_5430, wire_5278, wire_3891, wire_1314, wire_1256, wire_5553, wire_5509, wire_5508, wire_5443, wire_5442, wire_5417, wire_5416, wire_5270, wire_3889, wire_1314, wire_1256, wire_5555, wire_5495, wire_5494, wire_5469, wire_5468, wire_5403, wire_5402, wire_5262, wire_3887, wire_1310, wire_1256, wire_5557, wire_5481, wire_5480, wire_5455, wire_5454, wire_5429, wire_5428, wire_5254, wire_3885, wire_1310, wire_1256, wire_5559, wire_5507, wire_5506, wire_5441, wire_5440, wire_5415, wire_5414, wire_5246, wire_3883, wire_1310, wire_1256, wire_5521, wire_5493, wire_5492, wire_5467, wire_5466, wire_5401, wire_5400, wire_5398, wire_3881, wire_1310, wire_1256};
    // CHNAXY TOTAL: 880
    assign wire_3647 = lut_tile_4_3_chanxy_out[0];
    assign wire_3655 = lut_tile_4_3_chanxy_out[1];
    assign wire_3663 = lut_tile_4_3_chanxy_out[2];
    assign wire_3671 = lut_tile_4_3_chanxy_out[3];
    assign wire_3679 = lut_tile_4_3_chanxy_out[4];
    assign wire_3687 = lut_tile_4_3_chanxy_out[5];
    assign wire_3695 = lut_tile_4_3_chanxy_out[6];
    assign wire_3703 = lut_tile_4_3_chanxy_out[7];
    assign wire_3711 = lut_tile_4_3_chanxy_out[8];
    assign wire_3719 = lut_tile_4_3_chanxy_out[9];
    assign wire_3727 = lut_tile_4_3_chanxy_out[10];
    assign wire_3735 = lut_tile_4_3_chanxy_out[11];
    assign wire_3743 = lut_tile_4_3_chanxy_out[12];
    assign wire_3751 = lut_tile_4_3_chanxy_out[13];
    assign wire_3759 = lut_tile_4_3_chanxy_out[14];
    assign wire_3767 = lut_tile_4_3_chanxy_out[15];
    assign wire_3775 = lut_tile_4_3_chanxy_out[16];
    assign wire_3783 = lut_tile_4_3_chanxy_out[17];
    assign wire_3791 = lut_tile_4_3_chanxy_out[18];
    assign wire_3799 = lut_tile_4_3_chanxy_out[19];
    assign wire_3840 = lut_tile_4_3_chanxy_out[20];
    assign wire_3842 = lut_tile_4_3_chanxy_out[21];
    assign wire_3844 = lut_tile_4_3_chanxy_out[22];
    assign wire_3846 = lut_tile_4_3_chanxy_out[23];
    assign wire_3848 = lut_tile_4_3_chanxy_out[24];
    assign wire_3850 = lut_tile_4_3_chanxy_out[25];
    assign wire_3852 = lut_tile_4_3_chanxy_out[26];
    assign wire_3854 = lut_tile_4_3_chanxy_out[27];
    assign wire_3856 = lut_tile_4_3_chanxy_out[28];
    assign wire_3858 = lut_tile_4_3_chanxy_out[29];
    assign wire_3860 = lut_tile_4_3_chanxy_out[30];
    assign wire_3862 = lut_tile_4_3_chanxy_out[31];
    assign wire_3864 = lut_tile_4_3_chanxy_out[32];
    assign wire_3866 = lut_tile_4_3_chanxy_out[33];
    assign wire_3868 = lut_tile_4_3_chanxy_out[34];
    assign wire_3870 = lut_tile_4_3_chanxy_out[35];
    assign wire_3872 = lut_tile_4_3_chanxy_out[36];
    assign wire_3874 = lut_tile_4_3_chanxy_out[37];
    assign wire_3876 = lut_tile_4_3_chanxy_out[38];
    assign wire_3878 = lut_tile_4_3_chanxy_out[39];
    assign wire_5247 = lut_tile_4_3_chanxy_out[40];
    assign wire_5255 = lut_tile_4_3_chanxy_out[41];
    assign wire_5263 = lut_tile_4_3_chanxy_out[42];
    assign wire_5271 = lut_tile_4_3_chanxy_out[43];
    assign wire_5279 = lut_tile_4_3_chanxy_out[44];
    assign wire_5287 = lut_tile_4_3_chanxy_out[45];
    assign wire_5295 = lut_tile_4_3_chanxy_out[46];
    assign wire_5303 = lut_tile_4_3_chanxy_out[47];
    assign wire_5311 = lut_tile_4_3_chanxy_out[48];
    assign wire_5319 = lut_tile_4_3_chanxy_out[49];
    assign wire_5327 = lut_tile_4_3_chanxy_out[50];
    assign wire_5335 = lut_tile_4_3_chanxy_out[51];
    assign wire_5343 = lut_tile_4_3_chanxy_out[52];
    assign wire_5351 = lut_tile_4_3_chanxy_out[53];
    assign wire_5359 = lut_tile_4_3_chanxy_out[54];
    assign wire_5367 = lut_tile_4_3_chanxy_out[55];
    assign wire_5375 = lut_tile_4_3_chanxy_out[56];
    assign wire_5383 = lut_tile_4_3_chanxy_out[57];
    assign wire_5391 = lut_tile_4_3_chanxy_out[58];
    assign wire_5399 = lut_tile_4_3_chanxy_out[59];
    assign wire_5480 = lut_tile_4_3_chanxy_out[60];
    assign wire_5482 = lut_tile_4_3_chanxy_out[61];
    assign wire_5484 = lut_tile_4_3_chanxy_out[62];
    assign wire_5486 = lut_tile_4_3_chanxy_out[63];
    assign wire_5488 = lut_tile_4_3_chanxy_out[64];
    assign wire_5490 = lut_tile_4_3_chanxy_out[65];
    assign wire_5492 = lut_tile_4_3_chanxy_out[66];
    assign wire_5494 = lut_tile_4_3_chanxy_out[67];
    assign wire_5496 = lut_tile_4_3_chanxy_out[68];
    assign wire_5498 = lut_tile_4_3_chanxy_out[69];
    assign wire_5500 = lut_tile_4_3_chanxy_out[70];
    assign wire_5502 = lut_tile_4_3_chanxy_out[71];
    assign wire_5504 = lut_tile_4_3_chanxy_out[72];
    assign wire_5506 = lut_tile_4_3_chanxy_out[73];
    assign wire_5508 = lut_tile_4_3_chanxy_out[74];
    assign wire_5510 = lut_tile_4_3_chanxy_out[75];
    assign wire_5512 = lut_tile_4_3_chanxy_out[76];
    assign wire_5514 = lut_tile_4_3_chanxy_out[77];
    assign wire_5516 = lut_tile_4_3_chanxy_out[78];
    assign wire_5518 = lut_tile_4_3_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_4_4_chanxy_in = {wire_5718, wire_3601, wire_3599, wire_3598, wire_3533, wire_3532, wire_3507, wire_3506, wire_3334, wire_2011, wire_1637, wire_5710, wire_3639, wire_3585, wire_3584, wire_3559, wire_3558, wire_3493, wire_3492, wire_3342, wire_2011, wire_1637, wire_5702, wire_3637, wire_3571, wire_3570, wire_3545, wire_3544, wire_3519, wire_3518, wire_3350, wire_2011, wire_1637, wire_5694, wire_3635, wire_3597, wire_3596, wire_3531, wire_3530, wire_3505, wire_3504, wire_3358, wire_2011, wire_1637, wire_5686, wire_3633, wire_3583, wire_3582, wire_3557, wire_3556, wire_3491, wire_3490, wire_3366, wire_2011, wire_1633, wire_5678, wire_3631, wire_3569, wire_3568, wire_3543, wire_3542, wire_3517, wire_3516, wire_3374, wire_2011, wire_1633, wire_5670, wire_3629, wire_3595, wire_3594, wire_3529, wire_3528, wire_3503, wire_3502, wire_3382, wire_2011, wire_1633, wire_5662, wire_3627, wire_3581, wire_3580, wire_3555, wire_3554, wire_3489, wire_3488, wire_3390, wire_2011, wire_1633, wire_5654, wire_3625, wire_3567, wire_3566, wire_3541, wire_3540, wire_3515, wire_3514, wire_3398, wire_2007, wire_1633, wire_5646, wire_3623, wire_3593, wire_3592, wire_3527, wire_3526, wire_3501, wire_3500, wire_3406, wire_2007, wire_1633, wire_5638, wire_3621, wire_3579, wire_3578, wire_3553, wire_3552, wire_3487, wire_3486, wire_3414, wire_2007, wire_1633, wire_5630, wire_3619, wire_3565, wire_3564, wire_3539, wire_3538, wire_3513, wire_3512, wire_3422, wire_2007, wire_1633, wire_5622, wire_3617, wire_3591, wire_3590, wire_3525, wire_3524, wire_3499, wire_3498, wire_3430, wire_2007, wire_1629, wire_5614, wire_3615, wire_3577, wire_3576, wire_3551, wire_3550, wire_3485, wire_3484, wire_3438, wire_2007, wire_1629, wire_5606, wire_3613, wire_3563, wire_3562, wire_3537, wire_3536, wire_3511, wire_3510, wire_3446, wire_2007, wire_1629, wire_5598, wire_3611, wire_3589, wire_3588, wire_3523, wire_3522, wire_3497, wire_3496, wire_3454, wire_2007, wire_1629, wire_5590, wire_3609, wire_3575, wire_3574, wire_3549, wire_3548, wire_3483, wire_3482, wire_3462, wire_1637, wire_1629, wire_5582, wire_3607, wire_3561, wire_3560, wire_3535, wire_3534, wire_3509, wire_3508, wire_3470, wire_1637, wire_1629, wire_5574, wire_3605, wire_3587, wire_3586, wire_3521, wire_3520, wire_3495, wire_3494, wire_3478, wire_1637, wire_1629, wire_5566, wire_3603, wire_3573, wire_3572, wire_3547, wire_3546, wire_3481, wire_3480, wire_3326, wire_1637, wire_1629, wire_5879, wire_3959, wire_3919, wire_3918, wire_3853, wire_3852, wire_3827, wire_3826, wire_3640, wire_2011, wire_1637, wire_5877, wire_3921, wire_3905, wire_3904, wire_3879, wire_3878, wire_3813, wire_3812, wire_3792, wire_2011, wire_1637, wire_5875, wire_3923, wire_3891, wire_3890, wire_3865, wire_3864, wire_3839, wire_3838, wire_3784, wire_2011, wire_1637, wire_5873, wire_3925, wire_3917, wire_3916, wire_3851, wire_3850, wire_3825, wire_3824, wire_3776, wire_2011, wire_1637, wire_5871, wire_3927, wire_3903, wire_3902, wire_3877, wire_3876, wire_3811, wire_3810, wire_3768, wire_2011, wire_1633, wire_5869, wire_3929, wire_3889, wire_3888, wire_3863, wire_3862, wire_3837, wire_3836, wire_3760, wire_2011, wire_1633, wire_5867, wire_3931, wire_3915, wire_3914, wire_3849, wire_3848, wire_3823, wire_3822, wire_3752, wire_2011, wire_1633, wire_5865, wire_3933, wire_3901, wire_3900, wire_3875, wire_3874, wire_3809, wire_3808, wire_3744, wire_2011, wire_1633, wire_5863, wire_3935, wire_3887, wire_3886, wire_3861, wire_3860, wire_3835, wire_3834, wire_3736, wire_2007, wire_1633, wire_5861, wire_3937, wire_3913, wire_3912, wire_3847, wire_3846, wire_3821, wire_3820, wire_3728, wire_2007, wire_1633, wire_5859, wire_3939, wire_3899, wire_3898, wire_3873, wire_3872, wire_3807, wire_3806, wire_3720, wire_2007, wire_1633, wire_5857, wire_3941, wire_3885, wire_3884, wire_3859, wire_3858, wire_3833, wire_3832, wire_3712, wire_2007, wire_1633, wire_5855, wire_3943, wire_3911, wire_3910, wire_3845, wire_3844, wire_3819, wire_3818, wire_3704, wire_2007, wire_1629, wire_5853, wire_3945, wire_3897, wire_3896, wire_3871, wire_3870, wire_3805, wire_3804, wire_3696, wire_2007, wire_1629, wire_5851, wire_3947, wire_3883, wire_3882, wire_3857, wire_3856, wire_3831, wire_3830, wire_3688, wire_2007, wire_1629, wire_5849, wire_3949, wire_3909, wire_3908, wire_3843, wire_3842, wire_3817, wire_3816, wire_3680, wire_2007, wire_1629, wire_5847, wire_3951, wire_3895, wire_3894, wire_3869, wire_3868, wire_3803, wire_3802, wire_3672, wire_1637, wire_1629, wire_5845, wire_3953, wire_3881, wire_3880, wire_3855, wire_3854, wire_3829, wire_3828, wire_3664, wire_1637, wire_1629, wire_5843, wire_3955, wire_3907, wire_3906, wire_3841, wire_3840, wire_3815, wire_3814, wire_3656, wire_1637, wire_1629, wire_5841, wire_3957, wire_3893, wire_3892, wire_3867, wire_3866, wire_3801, wire_3800, wire_3648, wire_1637, wire_1629, wire_5557, wire_5519, wire_5518, wire_5453, wire_5452, wire_5427, wire_5426, wire_5398, wire_3798, wire_1694, wire_1686, wire_5555, wire_5505, wire_5504, wire_5479, wire_5478, wire_5413, wire_5412, wire_5246, wire_3790, wire_1694, wire_1686, wire_5553, wire_5491, wire_5490, wire_5465, wire_5464, wire_5439, wire_5438, wire_5254, wire_3782, wire_1694, wire_1686, wire_5551, wire_5517, wire_5516, wire_5451, wire_5450, wire_5425, wire_5424, wire_5262, wire_3774, wire_1694, wire_1686, wire_5549, wire_5503, wire_5502, wire_5477, wire_5476, wire_5411, wire_5410, wire_5270, wire_3766, wire_1694, wire_1636, wire_5547, wire_5489, wire_5488, wire_5463, wire_5462, wire_5437, wire_5436, wire_5278, wire_3758, wire_1694, wire_1636, wire_5545, wire_5515, wire_5514, wire_5449, wire_5448, wire_5423, wire_5422, wire_5286, wire_3750, wire_1694, wire_1636, wire_5543, wire_5501, wire_5500, wire_5475, wire_5474, wire_5409, wire_5408, wire_5294, wire_3742, wire_1694, wire_1636, wire_5541, wire_5487, wire_5486, wire_5461, wire_5460, wire_5435, wire_5434, wire_5302, wire_3734, wire_1690, wire_1636, wire_5539, wire_5513, wire_5512, wire_5447, wire_5446, wire_5421, wire_5420, wire_5310, wire_3726, wire_1690, wire_1636, wire_5537, wire_5499, wire_5498, wire_5473, wire_5472, wire_5407, wire_5406, wire_5318, wire_3718, wire_1690, wire_1636, wire_5535, wire_5485, wire_5484, wire_5459, wire_5458, wire_5433, wire_5432, wire_5326, wire_3710, wire_1690, wire_1636, wire_5533, wire_5511, wire_5510, wire_5445, wire_5444, wire_5419, wire_5418, wire_5334, wire_3702, wire_1690, wire_1632, wire_5531, wire_5497, wire_5496, wire_5471, wire_5470, wire_5405, wire_5404, wire_5342, wire_3694, wire_1690, wire_1632, wire_5529, wire_5483, wire_5482, wire_5457, wire_5456, wire_5431, wire_5430, wire_5350, wire_3686, wire_1690, wire_1632, wire_5527, wire_5509, wire_5508, wire_5443, wire_5442, wire_5417, wire_5416, wire_5358, wire_3678, wire_1690, wire_1632, wire_5525, wire_5495, wire_5494, wire_5469, wire_5468, wire_5403, wire_5402, wire_5366, wire_3670, wire_1686, wire_1632, wire_5523, wire_5481, wire_5480, wire_5455, wire_5454, wire_5429, wire_5428, wire_5374, wire_3662, wire_1686, wire_1632, wire_5521, wire_5507, wire_5506, wire_5441, wire_5440, wire_5415, wire_5414, wire_5382, wire_3654, wire_1686, wire_1632, wire_5559, wire_5493, wire_5492, wire_5467, wire_5466, wire_5401, wire_5400, wire_5390, wire_3646, wire_1686, wire_1632, wire_5843, wire_5839, wire_5838, wire_5773, wire_5772, wire_5747, wire_5746, wire_5704, wire_3959, wire_1694, wire_1686, wire_5845, wire_5825, wire_5824, wire_5799, wire_5798, wire_5733, wire_5732, wire_5696, wire_3957, wire_1694, wire_1686, wire_5847, wire_5811, wire_5810, wire_5785, wire_5784, wire_5759, wire_5758, wire_5688, wire_3955, wire_1694, wire_1686, wire_5849, wire_5837, wire_5836, wire_5771, wire_5770, wire_5745, wire_5744, wire_5680, wire_3953, wire_1694, wire_1686, wire_5851, wire_5823, wire_5822, wire_5797, wire_5796, wire_5731, wire_5730, wire_5672, wire_3951, wire_1694, wire_1636, wire_5853, wire_5809, wire_5808, wire_5783, wire_5782, wire_5757, wire_5756, wire_5664, wire_3949, wire_1694, wire_1636, wire_5855, wire_5835, wire_5834, wire_5769, wire_5768, wire_5743, wire_5742, wire_5656, wire_3947, wire_1694, wire_1636, wire_5857, wire_5821, wire_5820, wire_5795, wire_5794, wire_5729, wire_5728, wire_5648, wire_3945, wire_1694, wire_1636, wire_5859, wire_5807, wire_5806, wire_5781, wire_5780, wire_5755, wire_5754, wire_5640, wire_3943, wire_1690, wire_1636, wire_5861, wire_5833, wire_5832, wire_5767, wire_5766, wire_5741, wire_5740, wire_5632, wire_3941, wire_1690, wire_1636, wire_5863, wire_5819, wire_5818, wire_5793, wire_5792, wire_5727, wire_5726, wire_5624, wire_3939, wire_1690, wire_1636, wire_5865, wire_5805, wire_5804, wire_5779, wire_5778, wire_5753, wire_5752, wire_5616, wire_3937, wire_1690, wire_1636, wire_5867, wire_5831, wire_5830, wire_5765, wire_5764, wire_5739, wire_5738, wire_5608, wire_3935, wire_1690, wire_1632, wire_5869, wire_5817, wire_5816, wire_5791, wire_5790, wire_5725, wire_5724, wire_5600, wire_3933, wire_1690, wire_1632, wire_5871, wire_5803, wire_5802, wire_5777, wire_5776, wire_5751, wire_5750, wire_5592, wire_3931, wire_1690, wire_1632, wire_5873, wire_5829, wire_5828, wire_5763, wire_5762, wire_5737, wire_5736, wire_5584, wire_3929, wire_1690, wire_1632, wire_5875, wire_5815, wire_5814, wire_5789, wire_5788, wire_5723, wire_5722, wire_5576, wire_3927, wire_1686, wire_1632, wire_5877, wire_5801, wire_5800, wire_5775, wire_5774, wire_5749, wire_5748, wire_5568, wire_3925, wire_1686, wire_1632, wire_5879, wire_5827, wire_5826, wire_5761, wire_5760, wire_5735, wire_5734, wire_5560, wire_3923, wire_1686, wire_1632, wire_5841, wire_5813, wire_5812, wire_5787, wire_5786, wire_5721, wire_5720, wire_5712, wire_3921, wire_1686, wire_1632};
    // CHNAXY TOTAL: 880
    assign wire_3641 = lut_tile_4_4_chanxy_out[0];
    assign wire_3649 = lut_tile_4_4_chanxy_out[1];
    assign wire_3657 = lut_tile_4_4_chanxy_out[2];
    assign wire_3665 = lut_tile_4_4_chanxy_out[3];
    assign wire_3673 = lut_tile_4_4_chanxy_out[4];
    assign wire_3681 = lut_tile_4_4_chanxy_out[5];
    assign wire_3689 = lut_tile_4_4_chanxy_out[6];
    assign wire_3697 = lut_tile_4_4_chanxy_out[7];
    assign wire_3705 = lut_tile_4_4_chanxy_out[8];
    assign wire_3713 = lut_tile_4_4_chanxy_out[9];
    assign wire_3721 = lut_tile_4_4_chanxy_out[10];
    assign wire_3729 = lut_tile_4_4_chanxy_out[11];
    assign wire_3737 = lut_tile_4_4_chanxy_out[12];
    assign wire_3745 = lut_tile_4_4_chanxy_out[13];
    assign wire_3753 = lut_tile_4_4_chanxy_out[14];
    assign wire_3761 = lut_tile_4_4_chanxy_out[15];
    assign wire_3769 = lut_tile_4_4_chanxy_out[16];
    assign wire_3777 = lut_tile_4_4_chanxy_out[17];
    assign wire_3785 = lut_tile_4_4_chanxy_out[18];
    assign wire_3793 = lut_tile_4_4_chanxy_out[19];
    assign wire_3880 = lut_tile_4_4_chanxy_out[20];
    assign wire_3882 = lut_tile_4_4_chanxy_out[21];
    assign wire_3884 = lut_tile_4_4_chanxy_out[22];
    assign wire_3886 = lut_tile_4_4_chanxy_out[23];
    assign wire_3888 = lut_tile_4_4_chanxy_out[24];
    assign wire_3890 = lut_tile_4_4_chanxy_out[25];
    assign wire_3892 = lut_tile_4_4_chanxy_out[26];
    assign wire_3894 = lut_tile_4_4_chanxy_out[27];
    assign wire_3896 = lut_tile_4_4_chanxy_out[28];
    assign wire_3898 = lut_tile_4_4_chanxy_out[29];
    assign wire_3900 = lut_tile_4_4_chanxy_out[30];
    assign wire_3902 = lut_tile_4_4_chanxy_out[31];
    assign wire_3904 = lut_tile_4_4_chanxy_out[32];
    assign wire_3906 = lut_tile_4_4_chanxy_out[33];
    assign wire_3908 = lut_tile_4_4_chanxy_out[34];
    assign wire_3910 = lut_tile_4_4_chanxy_out[35];
    assign wire_3912 = lut_tile_4_4_chanxy_out[36];
    assign wire_3914 = lut_tile_4_4_chanxy_out[37];
    assign wire_3916 = lut_tile_4_4_chanxy_out[38];
    assign wire_3918 = lut_tile_4_4_chanxy_out[39];
    assign wire_5561 = lut_tile_4_4_chanxy_out[40];
    assign wire_5569 = lut_tile_4_4_chanxy_out[41];
    assign wire_5577 = lut_tile_4_4_chanxy_out[42];
    assign wire_5585 = lut_tile_4_4_chanxy_out[43];
    assign wire_5593 = lut_tile_4_4_chanxy_out[44];
    assign wire_5601 = lut_tile_4_4_chanxy_out[45];
    assign wire_5609 = lut_tile_4_4_chanxy_out[46];
    assign wire_5617 = lut_tile_4_4_chanxy_out[47];
    assign wire_5625 = lut_tile_4_4_chanxy_out[48];
    assign wire_5633 = lut_tile_4_4_chanxy_out[49];
    assign wire_5641 = lut_tile_4_4_chanxy_out[50];
    assign wire_5649 = lut_tile_4_4_chanxy_out[51];
    assign wire_5657 = lut_tile_4_4_chanxy_out[52];
    assign wire_5665 = lut_tile_4_4_chanxy_out[53];
    assign wire_5673 = lut_tile_4_4_chanxy_out[54];
    assign wire_5681 = lut_tile_4_4_chanxy_out[55];
    assign wire_5689 = lut_tile_4_4_chanxy_out[56];
    assign wire_5697 = lut_tile_4_4_chanxy_out[57];
    assign wire_5705 = lut_tile_4_4_chanxy_out[58];
    assign wire_5713 = lut_tile_4_4_chanxy_out[59];
    assign wire_5800 = lut_tile_4_4_chanxy_out[60];
    assign wire_5802 = lut_tile_4_4_chanxy_out[61];
    assign wire_5804 = lut_tile_4_4_chanxy_out[62];
    assign wire_5806 = lut_tile_4_4_chanxy_out[63];
    assign wire_5808 = lut_tile_4_4_chanxy_out[64];
    assign wire_5810 = lut_tile_4_4_chanxy_out[65];
    assign wire_5812 = lut_tile_4_4_chanxy_out[66];
    assign wire_5814 = lut_tile_4_4_chanxy_out[67];
    assign wire_5816 = lut_tile_4_4_chanxy_out[68];
    assign wire_5818 = lut_tile_4_4_chanxy_out[69];
    assign wire_5820 = lut_tile_4_4_chanxy_out[70];
    assign wire_5822 = lut_tile_4_4_chanxy_out[71];
    assign wire_5824 = lut_tile_4_4_chanxy_out[72];
    assign wire_5826 = lut_tile_4_4_chanxy_out[73];
    assign wire_5828 = lut_tile_4_4_chanxy_out[74];
    assign wire_5830 = lut_tile_4_4_chanxy_out[75];
    assign wire_5832 = lut_tile_4_4_chanxy_out[76];
    assign wire_5834 = lut_tile_4_4_chanxy_out[77];
    assign wire_5836 = lut_tile_4_4_chanxy_out[78];
    assign wire_5838 = lut_tile_4_4_chanxy_out[79];
   // CHANXY OUT
    assign lut_tile_4_5_chanxy_in = {wire_6032, wire_3638, wire_3628, wire_3618, wire_3608, wire_2307, wire_2301, wire_2292, wire_2013, wire_6024, wire_3598, wire_3588, wire_3578, wire_3568, wire_2307, wire_2301, wire_2292, wire_2013, wire_6016, wire_3558, wire_3548, wire_3538, wire_3528, wire_2307, wire_2301, wire_2292, wire_2013, wire_6008, wire_3518, wire_3508, wire_3498, wire_3488, wire_2307, wire_2301, wire_2292, wire_2013, wire_6000, wire_3636, wire_3626, wire_3616, wire_3606, wire_2307, wire_2298, wire_2292, wire_2009, wire_5992, wire_3596, wire_3586, wire_3576, wire_3566, wire_2307, wire_2298, wire_2292, wire_2009, wire_5984, wire_3556, wire_3546, wire_3536, wire_3526, wire_2307, wire_2298, wire_2292, wire_2009, wire_5976, wire_3516, wire_3506, wire_3496, wire_3486, wire_2307, wire_2298, wire_2292, wire_2009, wire_5968, wire_3634, wire_3624, wire_3614, wire_3604, wire_2304, wire_2298, wire_2289, wire_2009, wire_5960, wire_3594, wire_3584, wire_3574, wire_3564, wire_2304, wire_2298, wire_2289, wire_2009, wire_5952, wire_3554, wire_3544, wire_3534, wire_3524, wire_2304, wire_2298, wire_2289, wire_2009, wire_5944, wire_3514, wire_3504, wire_3494, wire_3484, wire_2304, wire_2298, wire_2289, wire_2009, wire_5936, wire_3632, wire_3622, wire_3612, wire_3602, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_5928, wire_3592, wire_3582, wire_3572, wire_3562, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_5920, wire_3552, wire_3542, wire_3532, wire_3522, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_5912, wire_3512, wire_3502, wire_3492, wire_3482, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_5904, wire_3630, wire_3620, wire_3610, wire_3600, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_5896, wire_3590, wire_3580, wire_3570, wire_3560, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_5888, wire_3550, wire_3540, wire_3530, wire_3520, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_5880, wire_3510, wire_3500, wire_3490, wire_3480, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_6199, wire_3918, wire_3908, wire_3898, wire_3888, wire_2307, wire_2301, wire_2292, wire_2013, wire_6197, wire_3878, wire_3868, wire_3858, wire_3848, wire_2307, wire_2301, wire_2292, wire_2013, wire_6195, wire_3838, wire_3828, wire_3818, wire_3808, wire_2307, wire_2301, wire_2292, wire_2013, wire_6193, wire_3958, wire_3948, wire_3938, wire_3928, wire_2307, wire_2301, wire_2292, wire_2013, wire_6191, wire_3916, wire_3906, wire_3896, wire_3886, wire_2307, wire_2298, wire_2292, wire_2009, wire_6189, wire_3876, wire_3866, wire_3856, wire_3846, wire_2307, wire_2298, wire_2292, wire_2009, wire_6187, wire_3836, wire_3826, wire_3816, wire_3806, wire_2307, wire_2298, wire_2292, wire_2009, wire_6185, wire_3956, wire_3946, wire_3936, wire_3926, wire_2307, wire_2298, wire_2292, wire_2009, wire_6183, wire_3914, wire_3904, wire_3894, wire_3884, wire_2304, wire_2298, wire_2289, wire_2009, wire_6181, wire_3874, wire_3864, wire_3854, wire_3844, wire_2304, wire_2298, wire_2289, wire_2009, wire_6179, wire_3834, wire_3824, wire_3814, wire_3804, wire_2304, wire_2298, wire_2289, wire_2009, wire_6177, wire_3954, wire_3944, wire_3934, wire_3924, wire_2304, wire_2298, wire_2289, wire_2009, wire_6175, wire_3912, wire_3902, wire_3892, wire_3882, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_6173, wire_3872, wire_3862, wire_3852, wire_3842, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_6171, wire_3832, wire_3822, wire_3812, wire_3802, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_6169, wire_3952, wire_3942, wire_3932, wire_3922, wire_2310, wire_2304, wire_2295, wire_2289, wire_2005, wire_6167, wire_3910, wire_3900, wire_3890, wire_3880, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_6165, wire_3870, wire_3860, wire_3850, wire_3840, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_6163, wire_3830, wire_3820, wire_3810, wire_3800, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_6161, wire_3950, wire_3940, wire_3930, wire_3920, wire_2310, wire_2301, wire_2295, wire_2013, wire_2005, wire_6199, wire_6034, wire_5877, wire_5839, wire_5838, wire_5773, wire_5772, wire_5747, wire_5746, wire_5712, wire_3792, wire_2070, wire_2062, wire_6139, wire_6138, wire_5875, wire_5825, wire_5824, wire_5799, wire_5798, wire_5733, wire_5732, wire_5560, wire_3784, wire_2070, wire_2062, wire_6177, wire_5946, wire_5873, wire_5811, wire_5810, wire_5785, wire_5784, wire_5759, wire_5758, wire_5568, wire_3776, wire_2070, wire_2062, wire_6055, wire_6054, wire_5871, wire_5837, wire_5836, wire_5771, wire_5770, wire_5745, wire_5744, wire_5576, wire_3768, wire_2070, wire_2062, wire_6115, wire_6114, wire_5869, wire_5823, wire_5822, wire_5797, wire_5796, wire_5731, wire_5730, wire_5584, wire_3760, wire_2070, wire_2012, wire_6155, wire_6154, wire_5867, wire_5809, wire_5808, wire_5783, wire_5782, wire_5757, wire_5756, wire_5592, wire_3752, wire_2070, wire_2012, wire_6193, wire_6010, wire_5865, wire_5835, wire_5834, wire_5769, wire_5768, wire_5743, wire_5742, wire_5600, wire_3744, wire_2070, wire_2012, wire_6133, wire_6132, wire_5863, wire_5821, wire_5820, wire_5795, wire_5794, wire_5729, wire_5728, wire_5608, wire_3736, wire_2070, wire_2012, wire_6171, wire_5922, wire_5861, wire_5807, wire_5806, wire_5781, wire_5780, wire_5755, wire_5754, wire_5616, wire_3728, wire_2066, wire_2012, wire_6049, wire_6048, wire_5859, wire_5833, wire_5832, wire_5767, wire_5766, wire_5741, wire_5740, wire_5624, wire_3720, wire_2066, wire_2012, wire_6109, wire_6108, wire_2070, wire_5857, wire_5819, wire_5818, wire_5793, wire_5792, wire_5727, wire_5726, wire_5632, wire_3712, wire_2066, wire_2012, wire_6149, wire_6148, wire_2070, wire_5855, wire_5805, wire_5804, wire_5779, wire_5778, wire_5753, wire_5752, wire_5640, wire_3704, wire_2066, wire_2012, wire_6187, wire_5986, wire_2066, wire_5853, wire_5831, wire_5830, wire_5765, wire_5764, wire_5739, wire_5738, wire_5648, wire_3696, wire_2066, wire_2008, wire_6127, wire_6126, wire_2066, wire_5851, wire_5817, wire_5816, wire_5791, wire_5790, wire_5725, wire_5724, wire_5656, wire_3688, wire_2066, wire_2008, wire_6165, wire_5898, wire_2062, wire_5849, wire_5803, wire_5802, wire_5777, wire_5776, wire_5751, wire_5750, wire_5664, wire_3680, wire_2066, wire_2008, wire_6043, wire_6042, wire_2062, wire_5847, wire_5829, wire_5828, wire_5763, wire_5762, wire_5737, wire_5736, wire_5672, wire_3672, wire_2066, wire_2008, wire_6103, wire_6102, wire_2012, wire_5845, wire_5815, wire_5814, wire_5789, wire_5788, wire_5723, wire_5722, wire_5680, wire_3664, wire_2062, wire_2008, wire_6143, wire_6142, wire_2012, wire_5843, wire_5801, wire_5800, wire_5775, wire_5774, wire_5749, wire_5748, wire_5688, wire_3656, wire_2062, wire_2008, wire_6181, wire_5962, wire_2008, wire_5841, wire_5827, wire_5826, wire_5761, wire_5760, wire_5735, wire_5734, wire_5696, wire_3648, wire_2062, wire_2008, wire_6121, wire_6120, wire_2008, wire_5879, wire_5813, wire_5812, wire_5787, wire_5786, wire_5721, wire_5720, wire_5704, wire_3640, wire_2062, wire_2008, wire_6119, wire_6118, wire_6179, wire_5954, wire_6097, wire_6096, wire_6137, wire_6136, wire_6157, wire_6156, wire_6075, wire_6074, wire_6113, wire_6112, wire_6173, wire_5930, wire_6091, wire_6090, wire_6131, wire_6130, wire_6151, wire_6150, wire_2070, wire_6069, wire_6068, wire_2070, wire_6107, wire_6106, wire_2066, wire_6167, wire_5906, wire_2066, wire_6085, wire_6084, wire_2062, wire_6125, wire_6124, wire_2062, wire_6145, wire_6144, wire_2012, wire_6063, wire_6062, wire_2012, wire_6101, wire_6100, wire_2008, wire_6161, wire_5882, wire_2008, wire_6059, wire_6058, wire_6159, wire_6158, wire_6057, wire_6056, wire_6197, wire_6026, wire_6175, wire_5938, wire_6195, wire_6018, wire_6053, wire_6052, wire_6153, wire_6152, wire_6051, wire_6050, wire_6191, wire_6002, wire_6169, wire_5914, wire_2070, wire_6189, wire_5994, wire_2070, wire_6047, wire_6046, wire_2066, wire_6147, wire_6146, wire_2066, wire_6045, wire_6044, wire_2062, wire_6185, wire_5978, wire_2062, wire_6163, wire_5890, wire_2012, wire_6183, wire_5970, wire_2012, wire_6041, wire_6040, wire_2008, wire_6141, wire_6140, wire_2008, wire_6079, wire_6078, wire_6117, wire_6116, wire_6077, wire_6076, wire_6095, wire_6094, wire_6135, wire_6134, wire_6093, wire_6092, wire_6073, wire_6072, wire_6111, wire_6110, wire_6071, wire_6070, wire_6089, wire_6088, wire_6129, wire_6128, wire_2070, wire_6087, wire_6086, wire_2070, wire_6067, wire_6066, wire_2066, wire_6105, wire_6104, wire_2066, wire_6065, wire_6064, wire_2062, wire_6083, wire_6082, wire_2062, wire_6123, wire_6122, wire_2012, wire_6081, wire_6080, wire_2012, wire_6061, wire_6060, wire_2008, wire_6099, wire_6098, wire_2008};
    // CHNAXY TOTAL: 796
    assign wire_3801 = lut_tile_4_5_chanxy_out[0];
    assign wire_3803 = lut_tile_4_5_chanxy_out[1];
    assign wire_3805 = lut_tile_4_5_chanxy_out[2];
    assign wire_3807 = lut_tile_4_5_chanxy_out[3];
    assign wire_3809 = lut_tile_4_5_chanxy_out[4];
    assign wire_3811 = lut_tile_4_5_chanxy_out[5];
    assign wire_3813 = lut_tile_4_5_chanxy_out[6];
    assign wire_3815 = lut_tile_4_5_chanxy_out[7];
    assign wire_3817 = lut_tile_4_5_chanxy_out[8];
    assign wire_3819 = lut_tile_4_5_chanxy_out[9];
    assign wire_3821 = lut_tile_4_5_chanxy_out[10];
    assign wire_3823 = lut_tile_4_5_chanxy_out[11];
    assign wire_3825 = lut_tile_4_5_chanxy_out[12];
    assign wire_3827 = lut_tile_4_5_chanxy_out[13];
    assign wire_3829 = lut_tile_4_5_chanxy_out[14];
    assign wire_3831 = lut_tile_4_5_chanxy_out[15];
    assign wire_3833 = lut_tile_4_5_chanxy_out[16];
    assign wire_3835 = lut_tile_4_5_chanxy_out[17];
    assign wire_3837 = lut_tile_4_5_chanxy_out[18];
    assign wire_3839 = lut_tile_4_5_chanxy_out[19];
    assign wire_3841 = lut_tile_4_5_chanxy_out[20];
    assign wire_3843 = lut_tile_4_5_chanxy_out[21];
    assign wire_3845 = lut_tile_4_5_chanxy_out[22];
    assign wire_3847 = lut_tile_4_5_chanxy_out[23];
    assign wire_3849 = lut_tile_4_5_chanxy_out[24];
    assign wire_3851 = lut_tile_4_5_chanxy_out[25];
    assign wire_3853 = lut_tile_4_5_chanxy_out[26];
    assign wire_3855 = lut_tile_4_5_chanxy_out[27];
    assign wire_3857 = lut_tile_4_5_chanxy_out[28];
    assign wire_3859 = lut_tile_4_5_chanxy_out[29];
    assign wire_3861 = lut_tile_4_5_chanxy_out[30];
    assign wire_3863 = lut_tile_4_5_chanxy_out[31];
    assign wire_3865 = lut_tile_4_5_chanxy_out[32];
    assign wire_3867 = lut_tile_4_5_chanxy_out[33];
    assign wire_3869 = lut_tile_4_5_chanxy_out[34];
    assign wire_3871 = lut_tile_4_5_chanxy_out[35];
    assign wire_3873 = lut_tile_4_5_chanxy_out[36];
    assign wire_3875 = lut_tile_4_5_chanxy_out[37];
    assign wire_3877 = lut_tile_4_5_chanxy_out[38];
    assign wire_3879 = lut_tile_4_5_chanxy_out[39];
    assign wire_3881 = lut_tile_4_5_chanxy_out[40];
    assign wire_3883 = lut_tile_4_5_chanxy_out[41];
    assign wire_3885 = lut_tile_4_5_chanxy_out[42];
    assign wire_3887 = lut_tile_4_5_chanxy_out[43];
    assign wire_3889 = lut_tile_4_5_chanxy_out[44];
    assign wire_3891 = lut_tile_4_5_chanxy_out[45];
    assign wire_3893 = lut_tile_4_5_chanxy_out[46];
    assign wire_3895 = lut_tile_4_5_chanxy_out[47];
    assign wire_3897 = lut_tile_4_5_chanxy_out[48];
    assign wire_3899 = lut_tile_4_5_chanxy_out[49];
    assign wire_3901 = lut_tile_4_5_chanxy_out[50];
    assign wire_3903 = lut_tile_4_5_chanxy_out[51];
    assign wire_3905 = lut_tile_4_5_chanxy_out[52];
    assign wire_3907 = lut_tile_4_5_chanxy_out[53];
    assign wire_3909 = lut_tile_4_5_chanxy_out[54];
    assign wire_3911 = lut_tile_4_5_chanxy_out[55];
    assign wire_3913 = lut_tile_4_5_chanxy_out[56];
    assign wire_3915 = lut_tile_4_5_chanxy_out[57];
    assign wire_3917 = lut_tile_4_5_chanxy_out[58];
    assign wire_3919 = lut_tile_4_5_chanxy_out[59];
    assign wire_3920 = lut_tile_4_5_chanxy_out[60];
    assign wire_3921 = lut_tile_4_5_chanxy_out[61];
    assign wire_3922 = lut_tile_4_5_chanxy_out[62];
    assign wire_3923 = lut_tile_4_5_chanxy_out[63];
    assign wire_3924 = lut_tile_4_5_chanxy_out[64];
    assign wire_3925 = lut_tile_4_5_chanxy_out[65];
    assign wire_3926 = lut_tile_4_5_chanxy_out[66];
    assign wire_3927 = lut_tile_4_5_chanxy_out[67];
    assign wire_3928 = lut_tile_4_5_chanxy_out[68];
    assign wire_3929 = lut_tile_4_5_chanxy_out[69];
    assign wire_3930 = lut_tile_4_5_chanxy_out[70];
    assign wire_3931 = lut_tile_4_5_chanxy_out[71];
    assign wire_3932 = lut_tile_4_5_chanxy_out[72];
    assign wire_3933 = lut_tile_4_5_chanxy_out[73];
    assign wire_3934 = lut_tile_4_5_chanxy_out[74];
    assign wire_3935 = lut_tile_4_5_chanxy_out[75];
    assign wire_3936 = lut_tile_4_5_chanxy_out[76];
    assign wire_3937 = lut_tile_4_5_chanxy_out[77];
    assign wire_3938 = lut_tile_4_5_chanxy_out[78];
    assign wire_3939 = lut_tile_4_5_chanxy_out[79];
    assign wire_3940 = lut_tile_4_5_chanxy_out[80];
    assign wire_3941 = lut_tile_4_5_chanxy_out[81];
    assign wire_3942 = lut_tile_4_5_chanxy_out[82];
    assign wire_3943 = lut_tile_4_5_chanxy_out[83];
    assign wire_3944 = lut_tile_4_5_chanxy_out[84];
    assign wire_3945 = lut_tile_4_5_chanxy_out[85];
    assign wire_3946 = lut_tile_4_5_chanxy_out[86];
    assign wire_3947 = lut_tile_4_5_chanxy_out[87];
    assign wire_3948 = lut_tile_4_5_chanxy_out[88];
    assign wire_3949 = lut_tile_4_5_chanxy_out[89];
    assign wire_3950 = lut_tile_4_5_chanxy_out[90];
    assign wire_3951 = lut_tile_4_5_chanxy_out[91];
    assign wire_3952 = lut_tile_4_5_chanxy_out[92];
    assign wire_3953 = lut_tile_4_5_chanxy_out[93];
    assign wire_3954 = lut_tile_4_5_chanxy_out[94];
    assign wire_3955 = lut_tile_4_5_chanxy_out[95];
    assign wire_3956 = lut_tile_4_5_chanxy_out[96];
    assign wire_3957 = lut_tile_4_5_chanxy_out[97];
    assign wire_3958 = lut_tile_4_5_chanxy_out[98];
    assign wire_3959 = lut_tile_4_5_chanxy_out[99];
    assign wire_5883 = lut_tile_4_5_chanxy_out[100];
    assign wire_5891 = lut_tile_4_5_chanxy_out[101];
    assign wire_5899 = lut_tile_4_5_chanxy_out[102];
    assign wire_5907 = lut_tile_4_5_chanxy_out[103];
    assign wire_5915 = lut_tile_4_5_chanxy_out[104];
    assign wire_5923 = lut_tile_4_5_chanxy_out[105];
    assign wire_5931 = lut_tile_4_5_chanxy_out[106];
    assign wire_5939 = lut_tile_4_5_chanxy_out[107];
    assign wire_5947 = lut_tile_4_5_chanxy_out[108];
    assign wire_5955 = lut_tile_4_5_chanxy_out[109];
    assign wire_5963 = lut_tile_4_5_chanxy_out[110];
    assign wire_5971 = lut_tile_4_5_chanxy_out[111];
    assign wire_5979 = lut_tile_4_5_chanxy_out[112];
    assign wire_5987 = lut_tile_4_5_chanxy_out[113];
    assign wire_5995 = lut_tile_4_5_chanxy_out[114];
    assign wire_6003 = lut_tile_4_5_chanxy_out[115];
    assign wire_6011 = lut_tile_4_5_chanxy_out[116];
    assign wire_6019 = lut_tile_4_5_chanxy_out[117];
    assign wire_6027 = lut_tile_4_5_chanxy_out[118];
    assign wire_6035 = lut_tile_4_5_chanxy_out[119];
    assign wire_6120 = lut_tile_4_5_chanxy_out[120];
    assign wire_6122 = lut_tile_4_5_chanxy_out[121];
    assign wire_6124 = lut_tile_4_5_chanxy_out[122];
    assign wire_6126 = lut_tile_4_5_chanxy_out[123];
    assign wire_6128 = lut_tile_4_5_chanxy_out[124];
    assign wire_6130 = lut_tile_4_5_chanxy_out[125];
    assign wire_6132 = lut_tile_4_5_chanxy_out[126];
    assign wire_6134 = lut_tile_4_5_chanxy_out[127];
    assign wire_6136 = lut_tile_4_5_chanxy_out[128];
    assign wire_6138 = lut_tile_4_5_chanxy_out[129];
    assign wire_6140 = lut_tile_4_5_chanxy_out[130];
    assign wire_6142 = lut_tile_4_5_chanxy_out[131];
    assign wire_6144 = lut_tile_4_5_chanxy_out[132];
    assign wire_6146 = lut_tile_4_5_chanxy_out[133];
    assign wire_6148 = lut_tile_4_5_chanxy_out[134];
    assign wire_6150 = lut_tile_4_5_chanxy_out[135];
    assign wire_6152 = lut_tile_4_5_chanxy_out[136];
    assign wire_6154 = lut_tile_4_5_chanxy_out[137];
    assign wire_6156 = lut_tile_4_5_chanxy_out[138];
    assign wire_6158 = lut_tile_4_5_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_5_1_chanxy_in = {wire_4159, wire_4116, wire_4754, wire_3801, wire_3799, wire_3798, wire_3745, wire_3744, wire_3693, wire_3692, wire_3650, wire_939, wire_565, wire_4111, wire_4110, wire_4746, wire_3839, wire_3797, wire_3796, wire_3743, wire_3742, wire_3689, wire_3688, wire_3658, wire_939, wire_565, wire_4157, wire_4108, wire_4738, wire_3837, wire_3793, wire_3792, wire_3741, wire_3740, wire_3687, wire_3686, wire_3666, wire_939, wire_565, wire_4023, wire_4022, wire_4730, wire_3835, wire_3791, wire_3790, wire_3737, wire_3736, wire_3685, wire_3684, wire_3674, wire_939, wire_565, wire_4017, wire_4016, wire_4722, wire_3833, wire_3789, wire_3788, wire_3735, wire_3734, wire_3682, wire_3681, wire_3680, wire_939, wire_561, wire_4015, wire_4014, wire_4714, wire_3831, wire_3785, wire_3784, wire_3733, wire_3732, wire_3690, wire_3679, wire_3678, wire_939, wire_561, wire_4153, wire_4092, wire_4706, wire_3829, wire_3783, wire_3782, wire_3729, wire_3728, wire_3698, wire_3677, wire_3676, wire_939, wire_561, wire_4087, wire_4086, wire_4698, wire_3827, wire_3781, wire_3780, wire_3727, wire_3726, wire_3706, wire_3673, wire_3672, wire_939, wire_561, wire_4151, wire_4084, wire_4690, wire_3825, wire_3777, wire_3776, wire_3725, wire_3724, wire_3714, wire_3671, wire_3670, wire_935, wire_561, wire_3999, wire_3998, wire_4682, wire_3823, wire_3775, wire_3774, wire_3722, wire_3721, wire_3720, wire_3669, wire_3668, wire_935, wire_561, wire_3993, wire_3992, wire_939, wire_4674, wire_3821, wire_3773, wire_3772, wire_3730, wire_3719, wire_3718, wire_3665, wire_3664, wire_935, wire_561, wire_3991, wire_3990, wire_939, wire_4666, wire_3819, wire_3769, wire_3768, wire_3738, wire_3717, wire_3716, wire_3663, wire_3662, wire_935, wire_561, wire_4147, wire_4068, wire_935, wire_4658, wire_3817, wire_3767, wire_3766, wire_3746, wire_3713, wire_3712, wire_3661, wire_3660, wire_935, wire_557, wire_4063, wire_4062, wire_935, wire_4650, wire_3815, wire_3765, wire_3764, wire_3754, wire_3711, wire_3710, wire_3657, wire_3656, wire_935, wire_557, wire_4145, wire_4060, wire_565, wire_4642, wire_3813, wire_3762, wire_3761, wire_3760, wire_3709, wire_3708, wire_3655, wire_3654, wire_935, wire_557, wire_3975, wire_3974, wire_565, wire_4634, wire_3811, wire_3770, wire_3759, wire_3758, wire_3705, wire_3704, wire_3653, wire_3652, wire_935, wire_557, wire_3969, wire_3968, wire_561, wire_4626, wire_3809, wire_3778, wire_3757, wire_3756, wire_3703, wire_3702, wire_3649, wire_3648, wire_565, wire_557, wire_3967, wire_3966, wire_561, wire_4618, wire_3807, wire_3786, wire_3753, wire_3752, wire_3701, wire_3700, wire_3647, wire_3646, wire_565, wire_557, wire_4141, wire_4044, wire_557, wire_4610, wire_3805, wire_3794, wire_3751, wire_3750, wire_3697, wire_3696, wire_3645, wire_3644, wire_565, wire_557, wire_4039, wire_4038, wire_557, wire_4602, wire_3803, wire_3749, wire_3748, wire_3695, wire_3694, wire_3642, wire_3641, wire_3640, wire_565, wire_557, wire_4115, wire_4114, wire_4033, wire_4032, wire_4027, wire_4026, wire_4135, wire_4020, wire_4103, wire_4102, wire_4097, wire_4096, wire_4091, wire_4090, wire_4009, wire_4008, wire_4003, wire_4002, wire_4129, wire_3996, wire_4079, wire_4078, wire_939, wire_4073, wire_4072, wire_939, wire_4067, wire_4066, wire_935, wire_3985, wire_3984, wire_935, wire_3979, wire_3978, wire_565, wire_4123, wire_3972, wire_565, wire_4055, wire_4054, wire_561, wire_4049, wire_4048, wire_561, wire_4043, wire_4042, wire_557, wire_3961, wire_3960, wire_557, wire_4119, wire_4118, wire_4035, wire_4034, wire_4031, wire_4030, wire_4025, wire_4024, wire_4105, wire_4104, wire_4155, wire_4100, wire_4095, wire_4094, wire_4011, wire_4010, wire_4007, wire_4006, wire_4001, wire_4000, wire_4081, wire_4080, wire_939, wire_4149, wire_4076, wire_939, wire_4071, wire_4070, wire_935, wire_3987, wire_3986, wire_935, wire_3983, wire_3982, wire_565, wire_3977, wire_3976, wire_565, wire_4057, wire_4056, wire_561, wire_4143, wire_4052, wire_561, wire_4047, wire_4046, wire_557, wire_3963, wire_3962, wire_557, wire_4139, wire_4036, wire_4113, wire_4112, wire_4137, wire_4028, wire_4107, wire_4106, wire_4019, wire_4018, wire_4099, wire_4098, wire_4133, wire_4012, wire_4089, wire_4088, wire_4131, wire_4004, wire_4083, wire_4082, wire_3995, wire_3994, wire_939, wire_4075, wire_4074, wire_939, wire_4127, wire_3988, wire_935, wire_4065, wire_4064, wire_935, wire_4125, wire_3980, wire_565, wire_4059, wire_4058, wire_565, wire_3971, wire_3970, wire_561, wire_4051, wire_4050, wire_561, wire_4121, wire_3964, wire_557, wire_4041, wire_4040, wire_557, wire_4558, wire_614, wire_4838, wire_4828, wire_4818, wire_4808, wire_4159, wire_614, wire_608, wire_599, wire_593, wire_4560, wire_614, wire_4440, wire_614, wire_4480, wire_614, wire_4520, wire_614, wire_4798, wire_4788, wire_4778, wire_4768, wire_4157, wire_614, wire_608, wire_599, wire_593, wire_4562, wire_614, wire_4442, wire_614, wire_4482, wire_614, wire_4522, wire_611, wire_4918, wire_4908, wire_4898, wire_4888, wire_4155, wire_614, wire_608, wire_599, wire_593, wire_4564, wire_611, wire_4444, wire_611, wire_4484, wire_611, wire_4524, wire_611, wire_4878, wire_4868, wire_4858, wire_4848, wire_4153, wire_614, wire_608, wire_599, wire_593, wire_4566, wire_611, wire_4446, wire_611, wire_4486, wire_611, wire_4526, wire_608, wire_4836, wire_4826, wire_4816, wire_4806, wire_4151, wire_614, wire_605, wire_599, wire_564, wire_4568, wire_608, wire_4448, wire_608, wire_4488, wire_608, wire_4528, wire_608, wire_4796, wire_4786, wire_4776, wire_4766, wire_4149, wire_614, wire_605, wire_599, wire_564, wire_4570, wire_608, wire_4450, wire_608, wire_4490, wire_608, wire_4530, wire_605, wire_4916, wire_4906, wire_4896, wire_4886, wire_4147, wire_614, wire_605, wire_599, wire_564, wire_4572, wire_605, wire_4452, wire_605, wire_4492, wire_605, wire_4532, wire_605, wire_4876, wire_4866, wire_4856, wire_4846, wire_4145, wire_614, wire_605, wire_599, wire_564, wire_4574, wire_605, wire_4454, wire_605, wire_4494, wire_605, wire_4534, wire_602, wire_4834, wire_4824, wire_4814, wire_4804, wire_4143, wire_611, wire_605, wire_596, wire_564, wire_4576, wire_602, wire_4456, wire_602, wire_4496, wire_602, wire_4536, wire_602, wire_4794, wire_4784, wire_4774, wire_4764, wire_4141, wire_611, wire_605, wire_596, wire_564, wire_4578, wire_602, wire_4458, wire_602, wire_4498, wire_602, wire_4538, wire_599, wire_4914, wire_4904, wire_4894, wire_4884, wire_4139, wire_611, wire_605, wire_596, wire_564, wire_4580, wire_599, wire_4460, wire_599, wire_4500, wire_599, wire_4540, wire_599, wire_4874, wire_4864, wire_4854, wire_4844, wire_4137, wire_611, wire_605, wire_596, wire_564, wire_4582, wire_599, wire_4462, wire_599, wire_4502, wire_599, wire_4542, wire_596, wire_4832, wire_4822, wire_4812, wire_4802, wire_4135, wire_611, wire_602, wire_596, wire_560, wire_4584, wire_596, wire_4464, wire_596, wire_4504, wire_596, wire_4544, wire_596, wire_4792, wire_4782, wire_4772, wire_4762, wire_4133, wire_611, wire_602, wire_596, wire_560, wire_4586, wire_596, wire_4466, wire_596, wire_4506, wire_596, wire_4546, wire_593, wire_4912, wire_4902, wire_4892, wire_4882, wire_4131, wire_611, wire_602, wire_596, wire_560, wire_4588, wire_593, wire_4468, wire_593, wire_4508, wire_593, wire_4548, wire_593, wire_4872, wire_4862, wire_4852, wire_4842, wire_4129, wire_611, wire_602, wire_596, wire_560, wire_4590, wire_593, wire_4470, wire_593, wire_4510, wire_593, wire_4550, wire_564, wire_4830, wire_4820, wire_4810, wire_4800, wire_4127, wire_608, wire_602, wire_593, wire_560, wire_4592, wire_564, wire_4472, wire_564, wire_4512, wire_564, wire_4552, wire_564, wire_4790, wire_4780, wire_4770, wire_4760, wire_4125, wire_608, wire_602, wire_593, wire_560, wire_4594, wire_564, wire_4474, wire_564, wire_4514, wire_564, wire_4554, wire_560, wire_4910, wire_4900, wire_4890, wire_4880, wire_4123, wire_608, wire_602, wire_593, wire_560, wire_4596, wire_560, wire_4476, wire_560, wire_4516, wire_560, wire_4556, wire_560, wire_4870, wire_4860, wire_4850, wire_4840, wire_4121, wire_608, wire_602, wire_593, wire_560, wire_4598, wire_560, wire_4478, wire_560, wire_4518, wire_560};
    // CHNAXY TOTAL: 760
    assign wire_3960 = lut_tile_5_1_chanxy_out[0];
    assign wire_3962 = lut_tile_5_1_chanxy_out[1];
    assign wire_3964 = lut_tile_5_1_chanxy_out[2];
    assign wire_3965 = lut_tile_5_1_chanxy_out[3];
    assign wire_3966 = lut_tile_5_1_chanxy_out[4];
    assign wire_3968 = lut_tile_5_1_chanxy_out[5];
    assign wire_3970 = lut_tile_5_1_chanxy_out[6];
    assign wire_3972 = lut_tile_5_1_chanxy_out[7];
    assign wire_3973 = lut_tile_5_1_chanxy_out[8];
    assign wire_3974 = lut_tile_5_1_chanxy_out[9];
    assign wire_3976 = lut_tile_5_1_chanxy_out[10];
    assign wire_3978 = lut_tile_5_1_chanxy_out[11];
    assign wire_3980 = lut_tile_5_1_chanxy_out[12];
    assign wire_3981 = lut_tile_5_1_chanxy_out[13];
    assign wire_3982 = lut_tile_5_1_chanxy_out[14];
    assign wire_3984 = lut_tile_5_1_chanxy_out[15];
    assign wire_3986 = lut_tile_5_1_chanxy_out[16];
    assign wire_3988 = lut_tile_5_1_chanxy_out[17];
    assign wire_3989 = lut_tile_5_1_chanxy_out[18];
    assign wire_3990 = lut_tile_5_1_chanxy_out[19];
    assign wire_3992 = lut_tile_5_1_chanxy_out[20];
    assign wire_3994 = lut_tile_5_1_chanxy_out[21];
    assign wire_3996 = lut_tile_5_1_chanxy_out[22];
    assign wire_3997 = lut_tile_5_1_chanxy_out[23];
    assign wire_3998 = lut_tile_5_1_chanxy_out[24];
    assign wire_4000 = lut_tile_5_1_chanxy_out[25];
    assign wire_4002 = lut_tile_5_1_chanxy_out[26];
    assign wire_4004 = lut_tile_5_1_chanxy_out[27];
    assign wire_4005 = lut_tile_5_1_chanxy_out[28];
    assign wire_4006 = lut_tile_5_1_chanxy_out[29];
    assign wire_4008 = lut_tile_5_1_chanxy_out[30];
    assign wire_4010 = lut_tile_5_1_chanxy_out[31];
    assign wire_4012 = lut_tile_5_1_chanxy_out[32];
    assign wire_4013 = lut_tile_5_1_chanxy_out[33];
    assign wire_4014 = lut_tile_5_1_chanxy_out[34];
    assign wire_4016 = lut_tile_5_1_chanxy_out[35];
    assign wire_4018 = lut_tile_5_1_chanxy_out[36];
    assign wire_4020 = lut_tile_5_1_chanxy_out[37];
    assign wire_4021 = lut_tile_5_1_chanxy_out[38];
    assign wire_4022 = lut_tile_5_1_chanxy_out[39];
    assign wire_4024 = lut_tile_5_1_chanxy_out[40];
    assign wire_4026 = lut_tile_5_1_chanxy_out[41];
    assign wire_4028 = lut_tile_5_1_chanxy_out[42];
    assign wire_4029 = lut_tile_5_1_chanxy_out[43];
    assign wire_4030 = lut_tile_5_1_chanxy_out[44];
    assign wire_4032 = lut_tile_5_1_chanxy_out[45];
    assign wire_4034 = lut_tile_5_1_chanxy_out[46];
    assign wire_4036 = lut_tile_5_1_chanxy_out[47];
    assign wire_4037 = lut_tile_5_1_chanxy_out[48];
    assign wire_4038 = lut_tile_5_1_chanxy_out[49];
    assign wire_4040 = lut_tile_5_1_chanxy_out[50];
    assign wire_4042 = lut_tile_5_1_chanxy_out[51];
    assign wire_4044 = lut_tile_5_1_chanxy_out[52];
    assign wire_4045 = lut_tile_5_1_chanxy_out[53];
    assign wire_4046 = lut_tile_5_1_chanxy_out[54];
    assign wire_4048 = lut_tile_5_1_chanxy_out[55];
    assign wire_4050 = lut_tile_5_1_chanxy_out[56];
    assign wire_4052 = lut_tile_5_1_chanxy_out[57];
    assign wire_4053 = lut_tile_5_1_chanxy_out[58];
    assign wire_4054 = lut_tile_5_1_chanxy_out[59];
    assign wire_4056 = lut_tile_5_1_chanxy_out[60];
    assign wire_4058 = lut_tile_5_1_chanxy_out[61];
    assign wire_4060 = lut_tile_5_1_chanxy_out[62];
    assign wire_4061 = lut_tile_5_1_chanxy_out[63];
    assign wire_4062 = lut_tile_5_1_chanxy_out[64];
    assign wire_4064 = lut_tile_5_1_chanxy_out[65];
    assign wire_4066 = lut_tile_5_1_chanxy_out[66];
    assign wire_4068 = lut_tile_5_1_chanxy_out[67];
    assign wire_4069 = lut_tile_5_1_chanxy_out[68];
    assign wire_4070 = lut_tile_5_1_chanxy_out[69];
    assign wire_4072 = lut_tile_5_1_chanxy_out[70];
    assign wire_4074 = lut_tile_5_1_chanxy_out[71];
    assign wire_4076 = lut_tile_5_1_chanxy_out[72];
    assign wire_4077 = lut_tile_5_1_chanxy_out[73];
    assign wire_4078 = lut_tile_5_1_chanxy_out[74];
    assign wire_4080 = lut_tile_5_1_chanxy_out[75];
    assign wire_4082 = lut_tile_5_1_chanxy_out[76];
    assign wire_4084 = lut_tile_5_1_chanxy_out[77];
    assign wire_4085 = lut_tile_5_1_chanxy_out[78];
    assign wire_4086 = lut_tile_5_1_chanxy_out[79];
    assign wire_4088 = lut_tile_5_1_chanxy_out[80];
    assign wire_4090 = lut_tile_5_1_chanxy_out[81];
    assign wire_4092 = lut_tile_5_1_chanxy_out[82];
    assign wire_4093 = lut_tile_5_1_chanxy_out[83];
    assign wire_4094 = lut_tile_5_1_chanxy_out[84];
    assign wire_4096 = lut_tile_5_1_chanxy_out[85];
    assign wire_4098 = lut_tile_5_1_chanxy_out[86];
    assign wire_4100 = lut_tile_5_1_chanxy_out[87];
    assign wire_4101 = lut_tile_5_1_chanxy_out[88];
    assign wire_4102 = lut_tile_5_1_chanxy_out[89];
    assign wire_4104 = lut_tile_5_1_chanxy_out[90];
    assign wire_4106 = lut_tile_5_1_chanxy_out[91];
    assign wire_4108 = lut_tile_5_1_chanxy_out[92];
    assign wire_4109 = lut_tile_5_1_chanxy_out[93];
    assign wire_4110 = lut_tile_5_1_chanxy_out[94];
    assign wire_4112 = lut_tile_5_1_chanxy_out[95];
    assign wire_4114 = lut_tile_5_1_chanxy_out[96];
    assign wire_4116 = lut_tile_5_1_chanxy_out[97];
    assign wire_4117 = lut_tile_5_1_chanxy_out[98];
    assign wire_4118 = lut_tile_5_1_chanxy_out[99];
    assign wire_4761 = lut_tile_5_1_chanxy_out[100];
    assign wire_4763 = lut_tile_5_1_chanxy_out[101];
    assign wire_4765 = lut_tile_5_1_chanxy_out[102];
    assign wire_4767 = lut_tile_5_1_chanxy_out[103];
    assign wire_4769 = lut_tile_5_1_chanxy_out[104];
    assign wire_4771 = lut_tile_5_1_chanxy_out[105];
    assign wire_4773 = lut_tile_5_1_chanxy_out[106];
    assign wire_4775 = lut_tile_5_1_chanxy_out[107];
    assign wire_4777 = lut_tile_5_1_chanxy_out[108];
    assign wire_4779 = lut_tile_5_1_chanxy_out[109];
    assign wire_4781 = lut_tile_5_1_chanxy_out[110];
    assign wire_4783 = lut_tile_5_1_chanxy_out[111];
    assign wire_4785 = lut_tile_5_1_chanxy_out[112];
    assign wire_4787 = lut_tile_5_1_chanxy_out[113];
    assign wire_4789 = lut_tile_5_1_chanxy_out[114];
    assign wire_4791 = lut_tile_5_1_chanxy_out[115];
    assign wire_4793 = lut_tile_5_1_chanxy_out[116];
    assign wire_4795 = lut_tile_5_1_chanxy_out[117];
    assign wire_4797 = lut_tile_5_1_chanxy_out[118];
    assign wire_4799 = lut_tile_5_1_chanxy_out[119];
    assign wire_4801 = lut_tile_5_1_chanxy_out[120];
    assign wire_4803 = lut_tile_5_1_chanxy_out[121];
    assign wire_4805 = lut_tile_5_1_chanxy_out[122];
    assign wire_4807 = lut_tile_5_1_chanxy_out[123];
    assign wire_4809 = lut_tile_5_1_chanxy_out[124];
    assign wire_4811 = lut_tile_5_1_chanxy_out[125];
    assign wire_4813 = lut_tile_5_1_chanxy_out[126];
    assign wire_4815 = lut_tile_5_1_chanxy_out[127];
    assign wire_4817 = lut_tile_5_1_chanxy_out[128];
    assign wire_4819 = lut_tile_5_1_chanxy_out[129];
    assign wire_4821 = lut_tile_5_1_chanxy_out[130];
    assign wire_4823 = lut_tile_5_1_chanxy_out[131];
    assign wire_4825 = lut_tile_5_1_chanxy_out[132];
    assign wire_4827 = lut_tile_5_1_chanxy_out[133];
    assign wire_4829 = lut_tile_5_1_chanxy_out[134];
    assign wire_4831 = lut_tile_5_1_chanxy_out[135];
    assign wire_4833 = lut_tile_5_1_chanxy_out[136];
    assign wire_4835 = lut_tile_5_1_chanxy_out[137];
    assign wire_4837 = lut_tile_5_1_chanxy_out[138];
    assign wire_4839 = lut_tile_5_1_chanxy_out[139];
    assign wire_4841 = lut_tile_5_1_chanxy_out[140];
    assign wire_4843 = lut_tile_5_1_chanxy_out[141];
    assign wire_4845 = lut_tile_5_1_chanxy_out[142];
    assign wire_4847 = lut_tile_5_1_chanxy_out[143];
    assign wire_4849 = lut_tile_5_1_chanxy_out[144];
    assign wire_4851 = lut_tile_5_1_chanxy_out[145];
    assign wire_4853 = lut_tile_5_1_chanxy_out[146];
    assign wire_4855 = lut_tile_5_1_chanxy_out[147];
    assign wire_4857 = lut_tile_5_1_chanxy_out[148];
    assign wire_4859 = lut_tile_5_1_chanxy_out[149];
    assign wire_4861 = lut_tile_5_1_chanxy_out[150];
    assign wire_4863 = lut_tile_5_1_chanxy_out[151];
    assign wire_4865 = lut_tile_5_1_chanxy_out[152];
    assign wire_4867 = lut_tile_5_1_chanxy_out[153];
    assign wire_4869 = lut_tile_5_1_chanxy_out[154];
    assign wire_4871 = lut_tile_5_1_chanxy_out[155];
    assign wire_4873 = lut_tile_5_1_chanxy_out[156];
    assign wire_4875 = lut_tile_5_1_chanxy_out[157];
    assign wire_4877 = lut_tile_5_1_chanxy_out[158];
    assign wire_4879 = lut_tile_5_1_chanxy_out[159];
    assign wire_4880 = lut_tile_5_1_chanxy_out[160];
    assign wire_4881 = lut_tile_5_1_chanxy_out[161];
    assign wire_4882 = lut_tile_5_1_chanxy_out[162];
    assign wire_4883 = lut_tile_5_1_chanxy_out[163];
    assign wire_4884 = lut_tile_5_1_chanxy_out[164];
    assign wire_4885 = lut_tile_5_1_chanxy_out[165];
    assign wire_4886 = lut_tile_5_1_chanxy_out[166];
    assign wire_4887 = lut_tile_5_1_chanxy_out[167];
    assign wire_4888 = lut_tile_5_1_chanxy_out[168];
    assign wire_4889 = lut_tile_5_1_chanxy_out[169];
    assign wire_4890 = lut_tile_5_1_chanxy_out[170];
    assign wire_4891 = lut_tile_5_1_chanxy_out[171];
    assign wire_4892 = lut_tile_5_1_chanxy_out[172];
    assign wire_4893 = lut_tile_5_1_chanxy_out[173];
    assign wire_4894 = lut_tile_5_1_chanxy_out[174];
    assign wire_4895 = lut_tile_5_1_chanxy_out[175];
    assign wire_4896 = lut_tile_5_1_chanxy_out[176];
    assign wire_4897 = lut_tile_5_1_chanxy_out[177];
    assign wire_4898 = lut_tile_5_1_chanxy_out[178];
    assign wire_4899 = lut_tile_5_1_chanxy_out[179];
    assign wire_4900 = lut_tile_5_1_chanxy_out[180];
    assign wire_4901 = lut_tile_5_1_chanxy_out[181];
    assign wire_4902 = lut_tile_5_1_chanxy_out[182];
    assign wire_4903 = lut_tile_5_1_chanxy_out[183];
    assign wire_4904 = lut_tile_5_1_chanxy_out[184];
    assign wire_4905 = lut_tile_5_1_chanxy_out[185];
    assign wire_4906 = lut_tile_5_1_chanxy_out[186];
    assign wire_4907 = lut_tile_5_1_chanxy_out[187];
    assign wire_4908 = lut_tile_5_1_chanxy_out[188];
    assign wire_4909 = lut_tile_5_1_chanxy_out[189];
    assign wire_4910 = lut_tile_5_1_chanxy_out[190];
    assign wire_4911 = lut_tile_5_1_chanxy_out[191];
    assign wire_4912 = lut_tile_5_1_chanxy_out[192];
    assign wire_4913 = lut_tile_5_1_chanxy_out[193];
    assign wire_4914 = lut_tile_5_1_chanxy_out[194];
    assign wire_4915 = lut_tile_5_1_chanxy_out[195];
    assign wire_4916 = lut_tile_5_1_chanxy_out[196];
    assign wire_4917 = lut_tile_5_1_chanxy_out[197];
    assign wire_4918 = lut_tile_5_1_chanxy_out[198];
    assign wire_4919 = lut_tile_5_1_chanxy_out[199];
   // CHANXY OUT
    assign lut_tile_5_2_chanxy_in = {wire_4139, wire_4138, wire_5076, wire_3841, wire_3813, wire_3812, wire_3799, wire_3798, wire_3745, wire_3744, wire_3652, wire_1315, wire_941, wire_4113, wire_4112, wire_5068, wire_3879, wire_3839, wire_3838, wire_3743, wire_3742, wire_3689, wire_3688, wire_3660, wire_1315, wire_941, wire_4137, wire_4136, wire_5060, wire_3877, wire_3825, wire_3824, wire_3793, wire_3792, wire_3687, wire_3686, wire_3668, wire_1315, wire_941, wire_4107, wire_4106, wire_5052, wire_3875, wire_3811, wire_3810, wire_3791, wire_3790, wire_3737, wire_3736, wire_3676, wire_1315, wire_941, wire_4019, wire_4018, wire_5044, wire_3873, wire_3837, wire_3836, wire_3735, wire_3734, wire_3684, wire_3681, wire_3680, wire_1315, wire_937, wire_4099, wire_4098, wire_5036, wire_3871, wire_3823, wire_3822, wire_3785, wire_3784, wire_3692, wire_3679, wire_3678, wire_1315, wire_937, wire_4133, wire_4132, wire_5028, wire_3869, wire_3809, wire_3808, wire_3783, wire_3782, wire_3729, wire_3728, wire_3700, wire_1315, wire_937, wire_4089, wire_4088, wire_5020, wire_3867, wire_3835, wire_3834, wire_3727, wire_3726, wire_3708, wire_3673, wire_3672, wire_1315, wire_937, wire_4131, wire_4130, wire_5012, wire_3865, wire_3821, wire_3820, wire_3777, wire_3776, wire_3716, wire_3671, wire_3670, wire_1311, wire_937, wire_4083, wire_4082, wire_5004, wire_3863, wire_3807, wire_3806, wire_3775, wire_3774, wire_3724, wire_3721, wire_3720, wire_1311, wire_937, wire_3995, wire_3994, wire_1315, wire_4996, wire_3861, wire_3833, wire_3832, wire_3732, wire_3719, wire_3718, wire_3665, wire_3664, wire_1311, wire_937, wire_4075, wire_4074, wire_1315, wire_4988, wire_3859, wire_3819, wire_3818, wire_3769, wire_3768, wire_3740, wire_3663, wire_3662, wire_1311, wire_937, wire_4127, wire_4126, wire_1311, wire_4980, wire_3857, wire_3805, wire_3804, wire_3767, wire_3766, wire_3748, wire_3713, wire_3712, wire_1311, wire_933, wire_4065, wire_4064, wire_1311, wire_4972, wire_3855, wire_3831, wire_3830, wire_3756, wire_3711, wire_3710, wire_3657, wire_3656, wire_1311, wire_933, wire_4125, wire_4124, wire_941, wire_4964, wire_3853, wire_3817, wire_3816, wire_3764, wire_3761, wire_3760, wire_3655, wire_3654, wire_1311, wire_933, wire_4059, wire_4058, wire_941, wire_4956, wire_3851, wire_3803, wire_3802, wire_3772, wire_3759, wire_3758, wire_3705, wire_3704, wire_1311, wire_933, wire_3971, wire_3970, wire_937, wire_4948, wire_3849, wire_3829, wire_3828, wire_3780, wire_3703, wire_3702, wire_3649, wire_3648, wire_941, wire_933, wire_4051, wire_4050, wire_937, wire_4940, wire_3847, wire_3815, wire_3814, wire_3788, wire_3753, wire_3752, wire_3647, wire_3646, wire_941, wire_933, wire_4121, wire_4120, wire_933, wire_4932, wire_3845, wire_3801, wire_3800, wire_3796, wire_3751, wire_3750, wire_3697, wire_3696, wire_941, wire_933, wire_4041, wire_4040, wire_933, wire_4924, wire_3843, wire_3827, wire_3826, wire_3695, wire_3694, wire_3644, wire_3641, wire_3640, wire_941, wire_933, wire_4159, wire_4158, wire_4197, wire_4110, wire_4157, wire_4156, wire_4175, wire_4022, wire_4017, wire_4016, wire_4173, wire_4014, wire_4153, wire_4152, wire_4191, wire_4086, wire_4151, wire_4150, wire_4169, wire_3998, wire_3993, wire_3992, wire_1315, wire_4167, wire_3990, wire_1315, wire_4147, wire_4146, wire_1311, wire_4185, wire_4062, wire_1311, wire_4145, wire_4144, wire_941, wire_4163, wire_3974, wire_941, wire_3969, wire_3968, wire_937, wire_4161, wire_3966, wire_937, wire_4141, wire_4140, wire_933, wire_4179, wire_4038, wire_933, wire_4115, wire_4114, wire_4033, wire_4032, wire_4027, wire_4026, wire_4135, wire_4134, wire_4195, wire_4102, wire_4097, wire_4096, wire_4091, wire_4090, wire_4009, wire_4008, wire_4003, wire_4002, wire_4129, wire_4128, wire_4189, wire_4078, wire_1315, wire_4073, wire_4072, wire_1315, wire_4067, wire_4066, wire_1311, wire_3985, wire_3984, wire_1311, wire_3979, wire_3978, wire_941, wire_4123, wire_4122, wire_941, wire_4183, wire_4054, wire_937, wire_4049, wire_4048, wire_937, wire_4043, wire_4042, wire_933, wire_3961, wire_3960, wire_933, wire_4199, wire_4118, wire_4035, wire_4034, wire_4177, wire_4030, wire_4025, wire_4024, wire_4105, wire_4104, wire_4155, wire_4154, wire_4193, wire_4094, wire_4011, wire_4010, wire_4171, wire_4006, wire_4001, wire_4000, wire_4081, wire_4080, wire_1315, wire_4149, wire_4148, wire_1315, wire_4187, wire_4070, wire_1311, wire_3987, wire_3986, wire_1311, wire_4165, wire_3982, wire_941, wire_3977, wire_3976, wire_941, wire_4057, wire_4056, wire_937, wire_4143, wire_4142, wire_937, wire_4181, wire_4046, wire_933, wire_3963, wire_3962, wire_933, wire_4838, wire_4828, wire_4818, wire_4808, wire_4116, wire_990, wire_984, wire_975, wire_969, wire_4798, wire_4788, wire_4778, wire_4768, wire_4108, wire_990, wire_984, wire_975, wire_969, wire_4918, wire_4908, wire_4898, wire_4888, wire_4100, wire_990, wire_984, wire_975, wire_969, wire_4878, wire_4868, wire_4858, wire_4848, wire_4092, wire_990, wire_984, wire_975, wire_969, wire_4836, wire_4826, wire_4816, wire_4806, wire_4084, wire_990, wire_981, wire_975, wire_940, wire_4796, wire_4786, wire_4776, wire_4766, wire_4076, wire_990, wire_981, wire_975, wire_940, wire_4916, wire_4906, wire_4896, wire_4886, wire_4068, wire_990, wire_981, wire_975, wire_940, wire_4876, wire_4866, wire_4856, wire_4846, wire_4060, wire_990, wire_981, wire_975, wire_940, wire_4834, wire_4824, wire_4814, wire_4804, wire_4052, wire_987, wire_981, wire_972, wire_940, wire_4794, wire_4784, wire_4774, wire_4764, wire_4044, wire_987, wire_981, wire_972, wire_940, wire_4914, wire_4904, wire_4894, wire_4884, wire_4036, wire_987, wire_981, wire_972, wire_940, wire_4874, wire_4864, wire_4854, wire_4844, wire_4028, wire_987, wire_981, wire_972, wire_940, wire_4832, wire_4822, wire_4812, wire_4802, wire_4020, wire_987, wire_978, wire_972, wire_936, wire_4792, wire_4782, wire_4772, wire_4762, wire_4012, wire_987, wire_978, wire_972, wire_936, wire_4912, wire_4902, wire_4892, wire_4882, wire_4004, wire_987, wire_978, wire_972, wire_936, wire_4872, wire_4862, wire_4852, wire_4842, wire_3996, wire_987, wire_978, wire_972, wire_936, wire_4830, wire_4820, wire_4810, wire_4800, wire_3988, wire_984, wire_978, wire_969, wire_936, wire_4790, wire_4780, wire_4770, wire_4760, wire_3980, wire_984, wire_978, wire_969, wire_936, wire_4910, wire_4900, wire_4890, wire_4880, wire_3972, wire_984, wire_978, wire_969, wire_936, wire_4870, wire_4860, wire_4850, wire_4840, wire_3964, wire_984, wire_978, wire_969, wire_936, wire_5118, wire_5108, wire_5098, wire_5088, wire_4199, wire_990, wire_984, wire_975, wire_969, wire_5238, wire_5228, wire_5218, wire_5208, wire_4197, wire_990, wire_984, wire_975, wire_969, wire_5198, wire_5188, wire_5178, wire_5168, wire_4195, wire_990, wire_984, wire_975, wire_969, wire_5158, wire_5148, wire_5138, wire_5128, wire_4193, wire_990, wire_984, wire_975, wire_969, wire_5116, wire_5106, wire_5096, wire_5086, wire_4191, wire_990, wire_981, wire_975, wire_940, wire_5236, wire_5226, wire_5216, wire_5206, wire_4189, wire_990, wire_981, wire_975, wire_940, wire_5196, wire_5186, wire_5176, wire_5166, wire_4187, wire_990, wire_981, wire_975, wire_940, wire_5156, wire_5146, wire_5136, wire_5126, wire_4185, wire_990, wire_981, wire_975, wire_940, wire_5114, wire_5104, wire_5094, wire_5084, wire_4183, wire_987, wire_981, wire_972, wire_940, wire_5234, wire_5224, wire_5214, wire_5204, wire_4181, wire_987, wire_981, wire_972, wire_940, wire_5194, wire_5184, wire_5174, wire_5164, wire_4179, wire_987, wire_981, wire_972, wire_940, wire_5154, wire_5144, wire_5134, wire_5124, wire_4177, wire_987, wire_981, wire_972, wire_940, wire_5112, wire_5102, wire_5092, wire_5082, wire_4175, wire_987, wire_978, wire_972, wire_936, wire_5232, wire_5222, wire_5212, wire_5202, wire_4173, wire_987, wire_978, wire_972, wire_936, wire_5192, wire_5182, wire_5172, wire_5162, wire_4171, wire_987, wire_978, wire_972, wire_936, wire_5152, wire_5142, wire_5132, wire_5122, wire_4169, wire_987, wire_978, wire_972, wire_936, wire_5110, wire_5100, wire_5090, wire_5080, wire_4167, wire_984, wire_978, wire_969, wire_936, wire_5230, wire_5220, wire_5210, wire_5200, wire_4165, wire_984, wire_978, wire_969, wire_936, wire_5190, wire_5180, wire_5170, wire_5160, wire_4163, wire_984, wire_978, wire_969, wire_936, wire_5150, wire_5140, wire_5130, wire_5120, wire_4161, wire_984, wire_978, wire_969, wire_936};
    // CHNAXY TOTAL: 780
    assign wire_3967 = lut_tile_5_2_chanxy_out[0];
    assign wire_3975 = lut_tile_5_2_chanxy_out[1];
    assign wire_3983 = lut_tile_5_2_chanxy_out[2];
    assign wire_3991 = lut_tile_5_2_chanxy_out[3];
    assign wire_3999 = lut_tile_5_2_chanxy_out[4];
    assign wire_4007 = lut_tile_5_2_chanxy_out[5];
    assign wire_4015 = lut_tile_5_2_chanxy_out[6];
    assign wire_4023 = lut_tile_5_2_chanxy_out[7];
    assign wire_4031 = lut_tile_5_2_chanxy_out[8];
    assign wire_4039 = lut_tile_5_2_chanxy_out[9];
    assign wire_4047 = lut_tile_5_2_chanxy_out[10];
    assign wire_4055 = lut_tile_5_2_chanxy_out[11];
    assign wire_4063 = lut_tile_5_2_chanxy_out[12];
    assign wire_4071 = lut_tile_5_2_chanxy_out[13];
    assign wire_4079 = lut_tile_5_2_chanxy_out[14];
    assign wire_4087 = lut_tile_5_2_chanxy_out[15];
    assign wire_4095 = lut_tile_5_2_chanxy_out[16];
    assign wire_4103 = lut_tile_5_2_chanxy_out[17];
    assign wire_4111 = lut_tile_5_2_chanxy_out[18];
    assign wire_4119 = lut_tile_5_2_chanxy_out[19];
    assign wire_4120 = lut_tile_5_2_chanxy_out[20];
    assign wire_4122 = lut_tile_5_2_chanxy_out[21];
    assign wire_4124 = lut_tile_5_2_chanxy_out[22];
    assign wire_4126 = lut_tile_5_2_chanxy_out[23];
    assign wire_4128 = lut_tile_5_2_chanxy_out[24];
    assign wire_4130 = lut_tile_5_2_chanxy_out[25];
    assign wire_4132 = lut_tile_5_2_chanxy_out[26];
    assign wire_4134 = lut_tile_5_2_chanxy_out[27];
    assign wire_4136 = lut_tile_5_2_chanxy_out[28];
    assign wire_4138 = lut_tile_5_2_chanxy_out[29];
    assign wire_4140 = lut_tile_5_2_chanxy_out[30];
    assign wire_4142 = lut_tile_5_2_chanxy_out[31];
    assign wire_4144 = lut_tile_5_2_chanxy_out[32];
    assign wire_4146 = lut_tile_5_2_chanxy_out[33];
    assign wire_4148 = lut_tile_5_2_chanxy_out[34];
    assign wire_4150 = lut_tile_5_2_chanxy_out[35];
    assign wire_4152 = lut_tile_5_2_chanxy_out[36];
    assign wire_4154 = lut_tile_5_2_chanxy_out[37];
    assign wire_4156 = lut_tile_5_2_chanxy_out[38];
    assign wire_4158 = lut_tile_5_2_chanxy_out[39];
    assign wire_5081 = lut_tile_5_2_chanxy_out[40];
    assign wire_5083 = lut_tile_5_2_chanxy_out[41];
    assign wire_5085 = lut_tile_5_2_chanxy_out[42];
    assign wire_5087 = lut_tile_5_2_chanxy_out[43];
    assign wire_5089 = lut_tile_5_2_chanxy_out[44];
    assign wire_5091 = lut_tile_5_2_chanxy_out[45];
    assign wire_5093 = lut_tile_5_2_chanxy_out[46];
    assign wire_5095 = lut_tile_5_2_chanxy_out[47];
    assign wire_5097 = lut_tile_5_2_chanxy_out[48];
    assign wire_5099 = lut_tile_5_2_chanxy_out[49];
    assign wire_5101 = lut_tile_5_2_chanxy_out[50];
    assign wire_5103 = lut_tile_5_2_chanxy_out[51];
    assign wire_5105 = lut_tile_5_2_chanxy_out[52];
    assign wire_5107 = lut_tile_5_2_chanxy_out[53];
    assign wire_5109 = lut_tile_5_2_chanxy_out[54];
    assign wire_5111 = lut_tile_5_2_chanxy_out[55];
    assign wire_5113 = lut_tile_5_2_chanxy_out[56];
    assign wire_5115 = lut_tile_5_2_chanxy_out[57];
    assign wire_5117 = lut_tile_5_2_chanxy_out[58];
    assign wire_5119 = lut_tile_5_2_chanxy_out[59];
    assign wire_5121 = lut_tile_5_2_chanxy_out[60];
    assign wire_5123 = lut_tile_5_2_chanxy_out[61];
    assign wire_5125 = lut_tile_5_2_chanxy_out[62];
    assign wire_5127 = lut_tile_5_2_chanxy_out[63];
    assign wire_5129 = lut_tile_5_2_chanxy_out[64];
    assign wire_5131 = lut_tile_5_2_chanxy_out[65];
    assign wire_5133 = lut_tile_5_2_chanxy_out[66];
    assign wire_5135 = lut_tile_5_2_chanxy_out[67];
    assign wire_5137 = lut_tile_5_2_chanxy_out[68];
    assign wire_5139 = lut_tile_5_2_chanxy_out[69];
    assign wire_5141 = lut_tile_5_2_chanxy_out[70];
    assign wire_5143 = lut_tile_5_2_chanxy_out[71];
    assign wire_5145 = lut_tile_5_2_chanxy_out[72];
    assign wire_5147 = lut_tile_5_2_chanxy_out[73];
    assign wire_5149 = lut_tile_5_2_chanxy_out[74];
    assign wire_5151 = lut_tile_5_2_chanxy_out[75];
    assign wire_5153 = lut_tile_5_2_chanxy_out[76];
    assign wire_5155 = lut_tile_5_2_chanxy_out[77];
    assign wire_5157 = lut_tile_5_2_chanxy_out[78];
    assign wire_5159 = lut_tile_5_2_chanxy_out[79];
    assign wire_5161 = lut_tile_5_2_chanxy_out[80];
    assign wire_5163 = lut_tile_5_2_chanxy_out[81];
    assign wire_5165 = lut_tile_5_2_chanxy_out[82];
    assign wire_5167 = lut_tile_5_2_chanxy_out[83];
    assign wire_5169 = lut_tile_5_2_chanxy_out[84];
    assign wire_5171 = lut_tile_5_2_chanxy_out[85];
    assign wire_5173 = lut_tile_5_2_chanxy_out[86];
    assign wire_5175 = lut_tile_5_2_chanxy_out[87];
    assign wire_5177 = lut_tile_5_2_chanxy_out[88];
    assign wire_5179 = lut_tile_5_2_chanxy_out[89];
    assign wire_5181 = lut_tile_5_2_chanxy_out[90];
    assign wire_5183 = lut_tile_5_2_chanxy_out[91];
    assign wire_5185 = lut_tile_5_2_chanxy_out[92];
    assign wire_5187 = lut_tile_5_2_chanxy_out[93];
    assign wire_5189 = lut_tile_5_2_chanxy_out[94];
    assign wire_5191 = lut_tile_5_2_chanxy_out[95];
    assign wire_5193 = lut_tile_5_2_chanxy_out[96];
    assign wire_5195 = lut_tile_5_2_chanxy_out[97];
    assign wire_5197 = lut_tile_5_2_chanxy_out[98];
    assign wire_5199 = lut_tile_5_2_chanxy_out[99];
    assign wire_5200 = lut_tile_5_2_chanxy_out[100];
    assign wire_5201 = lut_tile_5_2_chanxy_out[101];
    assign wire_5202 = lut_tile_5_2_chanxy_out[102];
    assign wire_5203 = lut_tile_5_2_chanxy_out[103];
    assign wire_5204 = lut_tile_5_2_chanxy_out[104];
    assign wire_5205 = lut_tile_5_2_chanxy_out[105];
    assign wire_5206 = lut_tile_5_2_chanxy_out[106];
    assign wire_5207 = lut_tile_5_2_chanxy_out[107];
    assign wire_5208 = lut_tile_5_2_chanxy_out[108];
    assign wire_5209 = lut_tile_5_2_chanxy_out[109];
    assign wire_5210 = lut_tile_5_2_chanxy_out[110];
    assign wire_5211 = lut_tile_5_2_chanxy_out[111];
    assign wire_5212 = lut_tile_5_2_chanxy_out[112];
    assign wire_5213 = lut_tile_5_2_chanxy_out[113];
    assign wire_5214 = lut_tile_5_2_chanxy_out[114];
    assign wire_5215 = lut_tile_5_2_chanxy_out[115];
    assign wire_5216 = lut_tile_5_2_chanxy_out[116];
    assign wire_5217 = lut_tile_5_2_chanxy_out[117];
    assign wire_5218 = lut_tile_5_2_chanxy_out[118];
    assign wire_5219 = lut_tile_5_2_chanxy_out[119];
    assign wire_5220 = lut_tile_5_2_chanxy_out[120];
    assign wire_5221 = lut_tile_5_2_chanxy_out[121];
    assign wire_5222 = lut_tile_5_2_chanxy_out[122];
    assign wire_5223 = lut_tile_5_2_chanxy_out[123];
    assign wire_5224 = lut_tile_5_2_chanxy_out[124];
    assign wire_5225 = lut_tile_5_2_chanxy_out[125];
    assign wire_5226 = lut_tile_5_2_chanxy_out[126];
    assign wire_5227 = lut_tile_5_2_chanxy_out[127];
    assign wire_5228 = lut_tile_5_2_chanxy_out[128];
    assign wire_5229 = lut_tile_5_2_chanxy_out[129];
    assign wire_5230 = lut_tile_5_2_chanxy_out[130];
    assign wire_5231 = lut_tile_5_2_chanxy_out[131];
    assign wire_5232 = lut_tile_5_2_chanxy_out[132];
    assign wire_5233 = lut_tile_5_2_chanxy_out[133];
    assign wire_5234 = lut_tile_5_2_chanxy_out[134];
    assign wire_5235 = lut_tile_5_2_chanxy_out[135];
    assign wire_5236 = lut_tile_5_2_chanxy_out[136];
    assign wire_5237 = lut_tile_5_2_chanxy_out[137];
    assign wire_5238 = lut_tile_5_2_chanxy_out[138];
    assign wire_5239 = lut_tile_5_2_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_5_3_chanxy_in = {wire_4199, wire_4198, wire_5398, wire_3881, wire_3879, wire_3878, wire_3813, wire_3812, wire_3745, wire_3744, wire_3654, wire_1691, wire_1317, wire_4035, wire_4034, wire_5390, wire_3919, wire_3865, wire_3864, wire_3839, wire_3838, wire_3689, wire_3688, wire_3662, wire_1691, wire_1317, wire_4177, wire_4176, wire_5382, wire_3917, wire_3851, wire_3850, wire_3825, wire_3824, wire_3793, wire_3792, wire_3670, wire_1691, wire_1317, wire_4217, wire_4024, wire_5374, wire_3915, wire_3877, wire_3876, wire_3811, wire_3810, wire_3737, wire_3736, wire_3678, wire_1691, wire_1317, wire_4237, wire_4104, wire_5366, wire_3913, wire_3863, wire_3862, wire_3837, wire_3836, wire_3686, wire_3681, wire_3680, wire_1691, wire_1313, wire_4155, wire_4154, wire_5358, wire_3911, wire_3849, wire_3848, wire_3823, wire_3822, wire_3785, wire_3784, wire_3694, wire_1691, wire_1313, wire_4193, wire_4192, wire_5350, wire_3909, wire_3875, wire_3874, wire_3809, wire_3808, wire_3729, wire_3728, wire_3702, wire_1691, wire_1313, wire_4011, wire_4010, wire_5342, wire_3907, wire_3861, wire_3860, wire_3835, wire_3834, wire_3710, wire_3673, wire_3672, wire_1691, wire_1313, wire_4171, wire_4170, wire_5334, wire_3905, wire_3847, wire_3846, wire_3821, wire_3820, wire_3777, wire_3776, wire_3718, wire_1687, wire_1313, wire_4211, wire_4000, wire_5326, wire_3903, wire_3873, wire_3872, wire_3807, wire_3806, wire_3726, wire_3721, wire_3720, wire_1687, wire_1313, wire_4231, wire_4080, wire_1691, wire_5318, wire_3901, wire_3859, wire_3858, wire_3833, wire_3832, wire_3734, wire_3665, wire_3664, wire_1687, wire_1313, wire_4149, wire_4148, wire_1691, wire_5310, wire_3899, wire_3845, wire_3844, wire_3819, wire_3818, wire_3769, wire_3768, wire_3742, wire_1687, wire_1313, wire_4187, wire_4186, wire_1687, wire_5302, wire_3897, wire_3871, wire_3870, wire_3805, wire_3804, wire_3750, wire_3713, wire_3712, wire_1687, wire_1309, wire_3987, wire_3986, wire_1687, wire_5294, wire_3895, wire_3857, wire_3856, wire_3831, wire_3830, wire_3758, wire_3657, wire_3656, wire_1687, wire_1309, wire_4165, wire_4164, wire_1317, wire_5286, wire_3893, wire_3843, wire_3842, wire_3817, wire_3816, wire_3766, wire_3761, wire_3760, wire_1687, wire_1309, wire_4205, wire_3976, wire_1317, wire_5278, wire_3891, wire_3869, wire_3868, wire_3803, wire_3802, wire_3774, wire_3705, wire_3704, wire_1687, wire_1309, wire_4225, wire_4056, wire_1313, wire_5270, wire_3889, wire_3855, wire_3854, wire_3829, wire_3828, wire_3782, wire_3649, wire_3648, wire_1317, wire_1309, wire_4143, wire_4142, wire_1313, wire_5262, wire_3887, wire_3841, wire_3840, wire_3815, wire_3814, wire_3790, wire_3753, wire_3752, wire_1317, wire_1309, wire_4181, wire_4180, wire_1309, wire_5254, wire_3885, wire_3867, wire_3866, wire_3801, wire_3800, wire_3798, wire_3697, wire_3696, wire_1317, wire_1309, wire_3963, wire_3962, wire_1309, wire_5246, wire_3883, wire_3853, wire_3852, wire_3827, wire_3826, wire_3646, wire_3641, wire_3640, wire_1317, wire_1309, wire_4139, wire_4138, wire_4239, wire_4112, wire_4137, wire_4136, wire_4107, wire_4106, wire_4019, wire_4018, wire_4099, wire_4098, wire_4133, wire_4132, wire_4233, wire_4088, wire_4131, wire_4130, wire_4083, wire_4082, wire_3995, wire_3994, wire_1691, wire_4075, wire_4074, wire_1691, wire_4127, wire_4126, wire_1687, wire_4227, wire_4064, wire_1687, wire_4125, wire_4124, wire_1317, wire_4059, wire_4058, wire_1317, wire_3971, wire_3970, wire_1313, wire_4051, wire_4050, wire_1313, wire_4121, wire_4120, wire_1309, wire_4221, wire_4040, wire_1309, wire_4159, wire_4158, wire_4197, wire_4196, wire_4157, wire_4156, wire_4175, wire_4174, wire_4215, wire_4016, wire_4173, wire_4172, wire_4153, wire_4152, wire_4191, wire_4190, wire_4151, wire_4150, wire_4169, wire_4168, wire_4209, wire_3992, wire_1691, wire_4167, wire_4166, wire_1691, wire_4147, wire_4146, wire_1687, wire_4185, wire_4184, wire_1687, wire_4145, wire_4144, wire_1317, wire_4163, wire_4162, wire_1317, wire_4203, wire_3968, wire_1313, wire_4161, wire_4160, wire_1313, wire_4141, wire_4140, wire_1309, wire_4179, wire_4178, wire_1309, wire_4115, wire_4114, wire_4219, wire_4032, wire_4027, wire_4026, wire_4135, wire_4134, wire_4195, wire_4194, wire_4235, wire_4096, wire_4091, wire_4090, wire_4213, wire_4008, wire_4003, wire_4002, wire_4129, wire_4128, wire_4189, wire_4188, wire_1691, wire_4229, wire_4072, wire_1691, wire_4067, wire_4066, wire_1687, wire_4207, wire_3984, wire_1687, wire_3979, wire_3978, wire_1317, wire_4123, wire_4122, wire_1317, wire_4183, wire_4182, wire_1313, wire_4223, wire_4048, wire_1313, wire_4043, wire_4042, wire_1309, wire_4201, wire_3960, wire_1309, wire_5118, wire_5108, wire_5098, wire_5088, wire_4118, wire_1366, wire_1360, wire_1351, wire_1345, wire_5238, wire_5228, wire_5218, wire_5208, wire_4110, wire_1366, wire_1360, wire_1351, wire_1345, wire_5198, wire_5188, wire_5178, wire_5168, wire_4102, wire_1366, wire_1360, wire_1351, wire_1345, wire_5158, wire_5148, wire_5138, wire_5128, wire_4094, wire_1366, wire_1360, wire_1351, wire_1345, wire_5116, wire_5106, wire_5096, wire_5086, wire_4086, wire_1366, wire_1357, wire_1351, wire_1316, wire_5236, wire_5226, wire_5216, wire_5206, wire_4078, wire_1366, wire_1357, wire_1351, wire_1316, wire_5196, wire_5186, wire_5176, wire_5166, wire_4070, wire_1366, wire_1357, wire_1351, wire_1316, wire_5156, wire_5146, wire_5136, wire_5126, wire_4062, wire_1366, wire_1357, wire_1351, wire_1316, wire_5114, wire_5104, wire_5094, wire_5084, wire_4054, wire_1363, wire_1357, wire_1348, wire_1316, wire_5234, wire_5224, wire_5214, wire_5204, wire_4046, wire_1363, wire_1357, wire_1348, wire_1316, wire_5194, wire_5184, wire_5174, wire_5164, wire_4038, wire_1363, wire_1357, wire_1348, wire_1316, wire_5154, wire_5144, wire_5134, wire_5124, wire_4030, wire_1363, wire_1357, wire_1348, wire_1316, wire_5112, wire_5102, wire_5092, wire_5082, wire_4022, wire_1363, wire_1354, wire_1348, wire_1312, wire_5232, wire_5222, wire_5212, wire_5202, wire_4014, wire_1363, wire_1354, wire_1348, wire_1312, wire_5192, wire_5182, wire_5172, wire_5162, wire_4006, wire_1363, wire_1354, wire_1348, wire_1312, wire_5152, wire_5142, wire_5132, wire_5122, wire_3998, wire_1363, wire_1354, wire_1348, wire_1312, wire_5110, wire_5100, wire_5090, wire_5080, wire_3990, wire_1360, wire_1354, wire_1345, wire_1312, wire_5230, wire_5220, wire_5210, wire_5200, wire_3982, wire_1360, wire_1354, wire_1345, wire_1312, wire_5190, wire_5180, wire_5170, wire_5160, wire_3974, wire_1360, wire_1354, wire_1345, wire_1312, wire_5150, wire_5140, wire_5130, wire_5120, wire_3966, wire_1360, wire_1354, wire_1345, wire_1312, wire_5558, wire_5548, wire_5538, wire_5528, wire_4239, wire_1366, wire_1360, wire_1351, wire_1345, wire_5518, wire_5508, wire_5498, wire_5488, wire_4237, wire_1366, wire_1360, wire_1351, wire_1345, wire_5478, wire_5468, wire_5458, wire_5448, wire_4235, wire_1366, wire_1360, wire_1351, wire_1345, wire_5438, wire_5428, wire_5418, wire_5408, wire_4233, wire_1366, wire_1360, wire_1351, wire_1345, wire_5556, wire_5546, wire_5536, wire_5526, wire_4231, wire_1366, wire_1357, wire_1351, wire_1316, wire_5516, wire_5506, wire_5496, wire_5486, wire_4229, wire_1366, wire_1357, wire_1351, wire_1316, wire_5476, wire_5466, wire_5456, wire_5446, wire_4227, wire_1366, wire_1357, wire_1351, wire_1316, wire_5436, wire_5426, wire_5416, wire_5406, wire_4225, wire_1366, wire_1357, wire_1351, wire_1316, wire_5554, wire_5544, wire_5534, wire_5524, wire_4223, wire_1363, wire_1357, wire_1348, wire_1316, wire_5514, wire_5504, wire_5494, wire_5484, wire_4221, wire_1363, wire_1357, wire_1348, wire_1316, wire_5474, wire_5464, wire_5454, wire_5444, wire_4219, wire_1363, wire_1357, wire_1348, wire_1316, wire_5434, wire_5424, wire_5414, wire_5404, wire_4217, wire_1363, wire_1357, wire_1348, wire_1316, wire_5552, wire_5542, wire_5532, wire_5522, wire_4215, wire_1363, wire_1354, wire_1348, wire_1312, wire_5512, wire_5502, wire_5492, wire_5482, wire_4213, wire_1363, wire_1354, wire_1348, wire_1312, wire_5472, wire_5462, wire_5452, wire_5442, wire_4211, wire_1363, wire_1354, wire_1348, wire_1312, wire_5432, wire_5422, wire_5412, wire_5402, wire_4209, wire_1363, wire_1354, wire_1348, wire_1312, wire_5550, wire_5540, wire_5530, wire_5520, wire_4207, wire_1360, wire_1354, wire_1345, wire_1312, wire_5510, wire_5500, wire_5490, wire_5480, wire_4205, wire_1360, wire_1354, wire_1345, wire_1312, wire_5470, wire_5460, wire_5450, wire_5440, wire_4203, wire_1360, wire_1354, wire_1345, wire_1312, wire_5430, wire_5420, wire_5410, wire_5400, wire_4201, wire_1360, wire_1354, wire_1345, wire_1312};
    // CHNAXY TOTAL: 780
    assign wire_3961 = lut_tile_5_3_chanxy_out[0];
    assign wire_3969 = lut_tile_5_3_chanxy_out[1];
    assign wire_3977 = lut_tile_5_3_chanxy_out[2];
    assign wire_3985 = lut_tile_5_3_chanxy_out[3];
    assign wire_3993 = lut_tile_5_3_chanxy_out[4];
    assign wire_4001 = lut_tile_5_3_chanxy_out[5];
    assign wire_4009 = lut_tile_5_3_chanxy_out[6];
    assign wire_4017 = lut_tile_5_3_chanxy_out[7];
    assign wire_4025 = lut_tile_5_3_chanxy_out[8];
    assign wire_4033 = lut_tile_5_3_chanxy_out[9];
    assign wire_4041 = lut_tile_5_3_chanxy_out[10];
    assign wire_4049 = lut_tile_5_3_chanxy_out[11];
    assign wire_4057 = lut_tile_5_3_chanxy_out[12];
    assign wire_4065 = lut_tile_5_3_chanxy_out[13];
    assign wire_4073 = lut_tile_5_3_chanxy_out[14];
    assign wire_4081 = lut_tile_5_3_chanxy_out[15];
    assign wire_4089 = lut_tile_5_3_chanxy_out[16];
    assign wire_4097 = lut_tile_5_3_chanxy_out[17];
    assign wire_4105 = lut_tile_5_3_chanxy_out[18];
    assign wire_4113 = lut_tile_5_3_chanxy_out[19];
    assign wire_4160 = lut_tile_5_3_chanxy_out[20];
    assign wire_4162 = lut_tile_5_3_chanxy_out[21];
    assign wire_4164 = lut_tile_5_3_chanxy_out[22];
    assign wire_4166 = lut_tile_5_3_chanxy_out[23];
    assign wire_4168 = lut_tile_5_3_chanxy_out[24];
    assign wire_4170 = lut_tile_5_3_chanxy_out[25];
    assign wire_4172 = lut_tile_5_3_chanxy_out[26];
    assign wire_4174 = lut_tile_5_3_chanxy_out[27];
    assign wire_4176 = lut_tile_5_3_chanxy_out[28];
    assign wire_4178 = lut_tile_5_3_chanxy_out[29];
    assign wire_4180 = lut_tile_5_3_chanxy_out[30];
    assign wire_4182 = lut_tile_5_3_chanxy_out[31];
    assign wire_4184 = lut_tile_5_3_chanxy_out[32];
    assign wire_4186 = lut_tile_5_3_chanxy_out[33];
    assign wire_4188 = lut_tile_5_3_chanxy_out[34];
    assign wire_4190 = lut_tile_5_3_chanxy_out[35];
    assign wire_4192 = lut_tile_5_3_chanxy_out[36];
    assign wire_4194 = lut_tile_5_3_chanxy_out[37];
    assign wire_4196 = lut_tile_5_3_chanxy_out[38];
    assign wire_4198 = lut_tile_5_3_chanxy_out[39];
    assign wire_5401 = lut_tile_5_3_chanxy_out[40];
    assign wire_5403 = lut_tile_5_3_chanxy_out[41];
    assign wire_5405 = lut_tile_5_3_chanxy_out[42];
    assign wire_5407 = lut_tile_5_3_chanxy_out[43];
    assign wire_5409 = lut_tile_5_3_chanxy_out[44];
    assign wire_5411 = lut_tile_5_3_chanxy_out[45];
    assign wire_5413 = lut_tile_5_3_chanxy_out[46];
    assign wire_5415 = lut_tile_5_3_chanxy_out[47];
    assign wire_5417 = lut_tile_5_3_chanxy_out[48];
    assign wire_5419 = lut_tile_5_3_chanxy_out[49];
    assign wire_5421 = lut_tile_5_3_chanxy_out[50];
    assign wire_5423 = lut_tile_5_3_chanxy_out[51];
    assign wire_5425 = lut_tile_5_3_chanxy_out[52];
    assign wire_5427 = lut_tile_5_3_chanxy_out[53];
    assign wire_5429 = lut_tile_5_3_chanxy_out[54];
    assign wire_5431 = lut_tile_5_3_chanxy_out[55];
    assign wire_5433 = lut_tile_5_3_chanxy_out[56];
    assign wire_5435 = lut_tile_5_3_chanxy_out[57];
    assign wire_5437 = lut_tile_5_3_chanxy_out[58];
    assign wire_5439 = lut_tile_5_3_chanxy_out[59];
    assign wire_5441 = lut_tile_5_3_chanxy_out[60];
    assign wire_5443 = lut_tile_5_3_chanxy_out[61];
    assign wire_5445 = lut_tile_5_3_chanxy_out[62];
    assign wire_5447 = lut_tile_5_3_chanxy_out[63];
    assign wire_5449 = lut_tile_5_3_chanxy_out[64];
    assign wire_5451 = lut_tile_5_3_chanxy_out[65];
    assign wire_5453 = lut_tile_5_3_chanxy_out[66];
    assign wire_5455 = lut_tile_5_3_chanxy_out[67];
    assign wire_5457 = lut_tile_5_3_chanxy_out[68];
    assign wire_5459 = lut_tile_5_3_chanxy_out[69];
    assign wire_5461 = lut_tile_5_3_chanxy_out[70];
    assign wire_5463 = lut_tile_5_3_chanxy_out[71];
    assign wire_5465 = lut_tile_5_3_chanxy_out[72];
    assign wire_5467 = lut_tile_5_3_chanxy_out[73];
    assign wire_5469 = lut_tile_5_3_chanxy_out[74];
    assign wire_5471 = lut_tile_5_3_chanxy_out[75];
    assign wire_5473 = lut_tile_5_3_chanxy_out[76];
    assign wire_5475 = lut_tile_5_3_chanxy_out[77];
    assign wire_5477 = lut_tile_5_3_chanxy_out[78];
    assign wire_5479 = lut_tile_5_3_chanxy_out[79];
    assign wire_5481 = lut_tile_5_3_chanxy_out[80];
    assign wire_5483 = lut_tile_5_3_chanxy_out[81];
    assign wire_5485 = lut_tile_5_3_chanxy_out[82];
    assign wire_5487 = lut_tile_5_3_chanxy_out[83];
    assign wire_5489 = lut_tile_5_3_chanxy_out[84];
    assign wire_5491 = lut_tile_5_3_chanxy_out[85];
    assign wire_5493 = lut_tile_5_3_chanxy_out[86];
    assign wire_5495 = lut_tile_5_3_chanxy_out[87];
    assign wire_5497 = lut_tile_5_3_chanxy_out[88];
    assign wire_5499 = lut_tile_5_3_chanxy_out[89];
    assign wire_5501 = lut_tile_5_3_chanxy_out[90];
    assign wire_5503 = lut_tile_5_3_chanxy_out[91];
    assign wire_5505 = lut_tile_5_3_chanxy_out[92];
    assign wire_5507 = lut_tile_5_3_chanxy_out[93];
    assign wire_5509 = lut_tile_5_3_chanxy_out[94];
    assign wire_5511 = lut_tile_5_3_chanxy_out[95];
    assign wire_5513 = lut_tile_5_3_chanxy_out[96];
    assign wire_5515 = lut_tile_5_3_chanxy_out[97];
    assign wire_5517 = lut_tile_5_3_chanxy_out[98];
    assign wire_5519 = lut_tile_5_3_chanxy_out[99];
    assign wire_5520 = lut_tile_5_3_chanxy_out[100];
    assign wire_5521 = lut_tile_5_3_chanxy_out[101];
    assign wire_5522 = lut_tile_5_3_chanxy_out[102];
    assign wire_5523 = lut_tile_5_3_chanxy_out[103];
    assign wire_5524 = lut_tile_5_3_chanxy_out[104];
    assign wire_5525 = lut_tile_5_3_chanxy_out[105];
    assign wire_5526 = lut_tile_5_3_chanxy_out[106];
    assign wire_5527 = lut_tile_5_3_chanxy_out[107];
    assign wire_5528 = lut_tile_5_3_chanxy_out[108];
    assign wire_5529 = lut_tile_5_3_chanxy_out[109];
    assign wire_5530 = lut_tile_5_3_chanxy_out[110];
    assign wire_5531 = lut_tile_5_3_chanxy_out[111];
    assign wire_5532 = lut_tile_5_3_chanxy_out[112];
    assign wire_5533 = lut_tile_5_3_chanxy_out[113];
    assign wire_5534 = lut_tile_5_3_chanxy_out[114];
    assign wire_5535 = lut_tile_5_3_chanxy_out[115];
    assign wire_5536 = lut_tile_5_3_chanxy_out[116];
    assign wire_5537 = lut_tile_5_3_chanxy_out[117];
    assign wire_5538 = lut_tile_5_3_chanxy_out[118];
    assign wire_5539 = lut_tile_5_3_chanxy_out[119];
    assign wire_5540 = lut_tile_5_3_chanxy_out[120];
    assign wire_5541 = lut_tile_5_3_chanxy_out[121];
    assign wire_5542 = lut_tile_5_3_chanxy_out[122];
    assign wire_5543 = lut_tile_5_3_chanxy_out[123];
    assign wire_5544 = lut_tile_5_3_chanxy_out[124];
    assign wire_5545 = lut_tile_5_3_chanxy_out[125];
    assign wire_5546 = lut_tile_5_3_chanxy_out[126];
    assign wire_5547 = lut_tile_5_3_chanxy_out[127];
    assign wire_5548 = lut_tile_5_3_chanxy_out[128];
    assign wire_5549 = lut_tile_5_3_chanxy_out[129];
    assign wire_5550 = lut_tile_5_3_chanxy_out[130];
    assign wire_5551 = lut_tile_5_3_chanxy_out[131];
    assign wire_5552 = lut_tile_5_3_chanxy_out[132];
    assign wire_5553 = lut_tile_5_3_chanxy_out[133];
    assign wire_5554 = lut_tile_5_3_chanxy_out[134];
    assign wire_5555 = lut_tile_5_3_chanxy_out[135];
    assign wire_5556 = lut_tile_5_3_chanxy_out[136];
    assign wire_5557 = lut_tile_5_3_chanxy_out[137];
    assign wire_5558 = lut_tile_5_3_chanxy_out[138];
    assign wire_5559 = lut_tile_5_3_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_5_4_chanxy_in = {wire_4279, wire_4114, wire_5712, wire_3921, wire_3919, wire_3918, wire_3853, wire_3852, wire_3827, wire_3826, wire_3648, wire_2067, wire_1693, wire_4219, wire_4218, wire_5704, wire_3959, wire_3905, wire_3904, wire_3879, wire_3878, wire_3813, wire_3812, wire_3656, wire_2067, wire_1693, wire_4257, wire_4026, wire_5696, wire_3957, wire_3891, wire_3890, wire_3865, wire_3864, wire_3839, wire_3838, wire_3664, wire_2067, wire_1693, wire_4135, wire_4134, wire_5688, wire_3955, wire_3917, wire_3916, wire_3851, wire_3850, wire_3825, wire_3824, wire_3672, wire_2067, wire_1693, wire_4195, wire_4194, wire_5680, wire_3953, wire_3903, wire_3902, wire_3877, wire_3876, wire_3811, wire_3810, wire_3680, wire_2067, wire_1689, wire_4235, wire_4234, wire_5672, wire_3951, wire_3889, wire_3888, wire_3863, wire_3862, wire_3837, wire_3836, wire_3688, wire_2067, wire_1689, wire_4273, wire_4090, wire_5664, wire_3949, wire_3915, wire_3914, wire_3849, wire_3848, wire_3823, wire_3822, wire_3696, wire_2067, wire_1689, wire_4213, wire_4212, wire_5656, wire_3947, wire_3901, wire_3900, wire_3875, wire_3874, wire_3809, wire_3808, wire_3704, wire_2067, wire_1689, wire_4251, wire_4002, wire_5648, wire_3945, wire_3887, wire_3886, wire_3861, wire_3860, wire_3835, wire_3834, wire_3712, wire_2063, wire_1689, wire_4129, wire_4128, wire_5640, wire_3943, wire_3913, wire_3912, wire_3847, wire_3846, wire_3821, wire_3820, wire_3720, wire_2063, wire_1689, wire_4189, wire_4188, wire_2067, wire_5632, wire_3941, wire_3899, wire_3898, wire_3873, wire_3872, wire_3807, wire_3806, wire_3728, wire_2063, wire_1689, wire_4229, wire_4228, wire_2067, wire_5624, wire_3939, wire_3885, wire_3884, wire_3859, wire_3858, wire_3833, wire_3832, wire_3736, wire_2063, wire_1689, wire_4267, wire_4066, wire_2063, wire_5616, wire_3937, wire_3911, wire_3910, wire_3845, wire_3844, wire_3819, wire_3818, wire_3744, wire_2063, wire_1685, wire_4207, wire_4206, wire_2063, wire_5608, wire_3935, wire_3897, wire_3896, wire_3871, wire_3870, wire_3805, wire_3804, wire_3752, wire_2063, wire_1685, wire_4245, wire_3978, wire_1693, wire_5600, wire_3933, wire_3883, wire_3882, wire_3857, wire_3856, wire_3831, wire_3830, wire_3760, wire_2063, wire_1685, wire_4123, wire_4122, wire_1693, wire_5592, wire_3931, wire_3909, wire_3908, wire_3843, wire_3842, wire_3817, wire_3816, wire_3768, wire_2063, wire_1685, wire_4183, wire_4182, wire_1689, wire_5584, wire_3929, wire_3895, wire_3894, wire_3869, wire_3868, wire_3803, wire_3802, wire_3776, wire_1693, wire_1685, wire_4223, wire_4222, wire_1689, wire_5576, wire_3927, wire_3881, wire_3880, wire_3855, wire_3854, wire_3829, wire_3828, wire_3784, wire_1693, wire_1685, wire_4261, wire_4042, wire_1685, wire_5568, wire_3925, wire_3907, wire_3906, wire_3841, wire_3840, wire_3815, wire_3814, wire_3792, wire_1693, wire_1685, wire_4201, wire_4200, wire_1685, wire_5560, wire_3923, wire_3893, wire_3892, wire_3867, wire_3866, wire_3801, wire_3800, wire_3640, wire_1693, wire_1685, wire_4199, wire_4198, wire_4259, wire_4034, wire_4177, wire_4176, wire_4217, wire_4216, wire_4237, wire_4236, wire_4155, wire_4154, wire_4193, wire_4192, wire_4253, wire_4010, wire_4171, wire_4170, wire_4211, wire_4210, wire_4231, wire_4230, wire_2067, wire_4149, wire_4148, wire_2067, wire_4187, wire_4186, wire_2063, wire_4247, wire_3986, wire_2063, wire_4165, wire_4164, wire_1693, wire_4205, wire_4204, wire_1693, wire_4225, wire_4224, wire_1689, wire_4143, wire_4142, wire_1689, wire_4181, wire_4180, wire_1685, wire_4241, wire_3962, wire_1685, wire_4139, wire_4138, wire_4239, wire_4238, wire_4137, wire_4136, wire_4277, wire_4106, wire_4255, wire_4018, wire_4275, wire_4098, wire_4133, wire_4132, wire_4233, wire_4232, wire_4131, wire_4130, wire_4271, wire_4082, wire_4249, wire_3994, wire_2067, wire_4269, wire_4074, wire_2067, wire_4127, wire_4126, wire_2063, wire_4227, wire_4226, wire_2063, wire_4125, wire_4124, wire_1693, wire_4265, wire_4058, wire_1693, wire_4243, wire_3970, wire_1689, wire_4263, wire_4050, wire_1689, wire_4121, wire_4120, wire_1685, wire_4221, wire_4220, wire_1685, wire_4159, wire_4158, wire_4197, wire_4196, wire_4157, wire_4156, wire_4175, wire_4174, wire_4215, wire_4214, wire_4173, wire_4172, wire_4153, wire_4152, wire_4191, wire_4190, wire_4151, wire_4150, wire_4169, wire_4168, wire_4209, wire_4208, wire_2067, wire_4167, wire_4166, wire_2067, wire_4147, wire_4146, wire_2063, wire_4185, wire_4184, wire_2063, wire_4145, wire_4144, wire_1693, wire_4163, wire_4162, wire_1693, wire_4203, wire_4202, wire_1689, wire_4161, wire_4160, wire_1689, wire_4141, wire_4140, wire_1685, wire_4179, wire_4178, wire_1685, wire_5558, wire_5548, wire_5538, wire_5528, wire_4112, wire_1742, wire_1736, wire_1727, wire_1721, wire_5518, wire_5508, wire_5498, wire_5488, wire_4104, wire_1742, wire_1736, wire_1727, wire_1721, wire_5478, wire_5468, wire_5458, wire_5448, wire_4096, wire_1742, wire_1736, wire_1727, wire_1721, wire_5438, wire_5428, wire_5418, wire_5408, wire_4088, wire_1742, wire_1736, wire_1727, wire_1721, wire_5556, wire_5546, wire_5536, wire_5526, wire_4080, wire_1742, wire_1733, wire_1727, wire_1692, wire_5516, wire_5506, wire_5496, wire_5486, wire_4072, wire_1742, wire_1733, wire_1727, wire_1692, wire_5476, wire_5466, wire_5456, wire_5446, wire_4064, wire_1742, wire_1733, wire_1727, wire_1692, wire_5436, wire_5426, wire_5416, wire_5406, wire_4056, wire_1742, wire_1733, wire_1727, wire_1692, wire_5554, wire_5544, wire_5534, wire_5524, wire_4048, wire_1739, wire_1733, wire_1724, wire_1692, wire_5514, wire_5504, wire_5494, wire_5484, wire_4040, wire_1739, wire_1733, wire_1724, wire_1692, wire_5474, wire_5464, wire_5454, wire_5444, wire_4032, wire_1739, wire_1733, wire_1724, wire_1692, wire_5434, wire_5424, wire_5414, wire_5404, wire_4024, wire_1739, wire_1733, wire_1724, wire_1692, wire_5552, wire_5542, wire_5532, wire_5522, wire_4016, wire_1739, wire_1730, wire_1724, wire_1688, wire_5512, wire_5502, wire_5492, wire_5482, wire_4008, wire_1739, wire_1730, wire_1724, wire_1688, wire_5472, wire_5462, wire_5452, wire_5442, wire_4000, wire_1739, wire_1730, wire_1724, wire_1688, wire_5432, wire_5422, wire_5412, wire_5402, wire_3992, wire_1739, wire_1730, wire_1724, wire_1688, wire_5550, wire_5540, wire_5530, wire_5520, wire_3984, wire_1736, wire_1730, wire_1721, wire_1688, wire_5510, wire_5500, wire_5490, wire_5480, wire_3976, wire_1736, wire_1730, wire_1721, wire_1688, wire_5470, wire_5460, wire_5450, wire_5440, wire_3968, wire_1736, wire_1730, wire_1721, wire_1688, wire_5430, wire_5420, wire_5410, wire_5400, wire_3960, wire_1736, wire_1730, wire_1721, wire_1688, wire_5838, wire_5828, wire_5818, wire_5808, wire_4279, wire_1742, wire_1736, wire_1727, wire_1721, wire_5798, wire_5788, wire_5778, wire_5768, wire_4277, wire_1742, wire_1736, wire_1727, wire_1721, wire_5758, wire_5748, wire_5738, wire_5728, wire_4275, wire_1742, wire_1736, wire_1727, wire_1721, wire_5878, wire_5868, wire_5858, wire_5848, wire_4273, wire_1742, wire_1736, wire_1727, wire_1721, wire_5836, wire_5826, wire_5816, wire_5806, wire_4271, wire_1742, wire_1733, wire_1727, wire_1692, wire_5796, wire_5786, wire_5776, wire_5766, wire_4269, wire_1742, wire_1733, wire_1727, wire_1692, wire_5756, wire_5746, wire_5736, wire_5726, wire_4267, wire_1742, wire_1733, wire_1727, wire_1692, wire_5876, wire_5866, wire_5856, wire_5846, wire_4265, wire_1742, wire_1733, wire_1727, wire_1692, wire_5834, wire_5824, wire_5814, wire_5804, wire_4263, wire_1739, wire_1733, wire_1724, wire_1692, wire_5794, wire_5784, wire_5774, wire_5764, wire_4261, wire_1739, wire_1733, wire_1724, wire_1692, wire_5754, wire_5744, wire_5734, wire_5724, wire_4259, wire_1739, wire_1733, wire_1724, wire_1692, wire_5874, wire_5864, wire_5854, wire_5844, wire_4257, wire_1739, wire_1733, wire_1724, wire_1692, wire_5832, wire_5822, wire_5812, wire_5802, wire_4255, wire_1739, wire_1730, wire_1724, wire_1688, wire_5792, wire_5782, wire_5772, wire_5762, wire_4253, wire_1739, wire_1730, wire_1724, wire_1688, wire_5752, wire_5742, wire_5732, wire_5722, wire_4251, wire_1739, wire_1730, wire_1724, wire_1688, wire_5872, wire_5862, wire_5852, wire_5842, wire_4249, wire_1739, wire_1730, wire_1724, wire_1688, wire_5830, wire_5820, wire_5810, wire_5800, wire_4247, wire_1736, wire_1730, wire_1721, wire_1688, wire_5790, wire_5780, wire_5770, wire_5760, wire_4245, wire_1736, wire_1730, wire_1721, wire_1688, wire_5750, wire_5740, wire_5730, wire_5720, wire_4243, wire_1736, wire_1730, wire_1721, wire_1688, wire_5870, wire_5860, wire_5850, wire_5840, wire_4241, wire_1736, wire_1730, wire_1721, wire_1688};
    // CHNAXY TOTAL: 780
    assign wire_3963 = lut_tile_5_4_chanxy_out[0];
    assign wire_3971 = lut_tile_5_4_chanxy_out[1];
    assign wire_3979 = lut_tile_5_4_chanxy_out[2];
    assign wire_3987 = lut_tile_5_4_chanxy_out[3];
    assign wire_3995 = lut_tile_5_4_chanxy_out[4];
    assign wire_4003 = lut_tile_5_4_chanxy_out[5];
    assign wire_4011 = lut_tile_5_4_chanxy_out[6];
    assign wire_4019 = lut_tile_5_4_chanxy_out[7];
    assign wire_4027 = lut_tile_5_4_chanxy_out[8];
    assign wire_4035 = lut_tile_5_4_chanxy_out[9];
    assign wire_4043 = lut_tile_5_4_chanxy_out[10];
    assign wire_4051 = lut_tile_5_4_chanxy_out[11];
    assign wire_4059 = lut_tile_5_4_chanxy_out[12];
    assign wire_4067 = lut_tile_5_4_chanxy_out[13];
    assign wire_4075 = lut_tile_5_4_chanxy_out[14];
    assign wire_4083 = lut_tile_5_4_chanxy_out[15];
    assign wire_4091 = lut_tile_5_4_chanxy_out[16];
    assign wire_4099 = lut_tile_5_4_chanxy_out[17];
    assign wire_4107 = lut_tile_5_4_chanxy_out[18];
    assign wire_4115 = lut_tile_5_4_chanxy_out[19];
    assign wire_4200 = lut_tile_5_4_chanxy_out[20];
    assign wire_4202 = lut_tile_5_4_chanxy_out[21];
    assign wire_4204 = lut_tile_5_4_chanxy_out[22];
    assign wire_4206 = lut_tile_5_4_chanxy_out[23];
    assign wire_4208 = lut_tile_5_4_chanxy_out[24];
    assign wire_4210 = lut_tile_5_4_chanxy_out[25];
    assign wire_4212 = lut_tile_5_4_chanxy_out[26];
    assign wire_4214 = lut_tile_5_4_chanxy_out[27];
    assign wire_4216 = lut_tile_5_4_chanxy_out[28];
    assign wire_4218 = lut_tile_5_4_chanxy_out[29];
    assign wire_4220 = lut_tile_5_4_chanxy_out[30];
    assign wire_4222 = lut_tile_5_4_chanxy_out[31];
    assign wire_4224 = lut_tile_5_4_chanxy_out[32];
    assign wire_4226 = lut_tile_5_4_chanxy_out[33];
    assign wire_4228 = lut_tile_5_4_chanxy_out[34];
    assign wire_4230 = lut_tile_5_4_chanxy_out[35];
    assign wire_4232 = lut_tile_5_4_chanxy_out[36];
    assign wire_4234 = lut_tile_5_4_chanxy_out[37];
    assign wire_4236 = lut_tile_5_4_chanxy_out[38];
    assign wire_4238 = lut_tile_5_4_chanxy_out[39];
    assign wire_5721 = lut_tile_5_4_chanxy_out[40];
    assign wire_5723 = lut_tile_5_4_chanxy_out[41];
    assign wire_5725 = lut_tile_5_4_chanxy_out[42];
    assign wire_5727 = lut_tile_5_4_chanxy_out[43];
    assign wire_5729 = lut_tile_5_4_chanxy_out[44];
    assign wire_5731 = lut_tile_5_4_chanxy_out[45];
    assign wire_5733 = lut_tile_5_4_chanxy_out[46];
    assign wire_5735 = lut_tile_5_4_chanxy_out[47];
    assign wire_5737 = lut_tile_5_4_chanxy_out[48];
    assign wire_5739 = lut_tile_5_4_chanxy_out[49];
    assign wire_5741 = lut_tile_5_4_chanxy_out[50];
    assign wire_5743 = lut_tile_5_4_chanxy_out[51];
    assign wire_5745 = lut_tile_5_4_chanxy_out[52];
    assign wire_5747 = lut_tile_5_4_chanxy_out[53];
    assign wire_5749 = lut_tile_5_4_chanxy_out[54];
    assign wire_5751 = lut_tile_5_4_chanxy_out[55];
    assign wire_5753 = lut_tile_5_4_chanxy_out[56];
    assign wire_5755 = lut_tile_5_4_chanxy_out[57];
    assign wire_5757 = lut_tile_5_4_chanxy_out[58];
    assign wire_5759 = lut_tile_5_4_chanxy_out[59];
    assign wire_5761 = lut_tile_5_4_chanxy_out[60];
    assign wire_5763 = lut_tile_5_4_chanxy_out[61];
    assign wire_5765 = lut_tile_5_4_chanxy_out[62];
    assign wire_5767 = lut_tile_5_4_chanxy_out[63];
    assign wire_5769 = lut_tile_5_4_chanxy_out[64];
    assign wire_5771 = lut_tile_5_4_chanxy_out[65];
    assign wire_5773 = lut_tile_5_4_chanxy_out[66];
    assign wire_5775 = lut_tile_5_4_chanxy_out[67];
    assign wire_5777 = lut_tile_5_4_chanxy_out[68];
    assign wire_5779 = lut_tile_5_4_chanxy_out[69];
    assign wire_5781 = lut_tile_5_4_chanxy_out[70];
    assign wire_5783 = lut_tile_5_4_chanxy_out[71];
    assign wire_5785 = lut_tile_5_4_chanxy_out[72];
    assign wire_5787 = lut_tile_5_4_chanxy_out[73];
    assign wire_5789 = lut_tile_5_4_chanxy_out[74];
    assign wire_5791 = lut_tile_5_4_chanxy_out[75];
    assign wire_5793 = lut_tile_5_4_chanxy_out[76];
    assign wire_5795 = lut_tile_5_4_chanxy_out[77];
    assign wire_5797 = lut_tile_5_4_chanxy_out[78];
    assign wire_5799 = lut_tile_5_4_chanxy_out[79];
    assign wire_5801 = lut_tile_5_4_chanxy_out[80];
    assign wire_5803 = lut_tile_5_4_chanxy_out[81];
    assign wire_5805 = lut_tile_5_4_chanxy_out[82];
    assign wire_5807 = lut_tile_5_4_chanxy_out[83];
    assign wire_5809 = lut_tile_5_4_chanxy_out[84];
    assign wire_5811 = lut_tile_5_4_chanxy_out[85];
    assign wire_5813 = lut_tile_5_4_chanxy_out[86];
    assign wire_5815 = lut_tile_5_4_chanxy_out[87];
    assign wire_5817 = lut_tile_5_4_chanxy_out[88];
    assign wire_5819 = lut_tile_5_4_chanxy_out[89];
    assign wire_5821 = lut_tile_5_4_chanxy_out[90];
    assign wire_5823 = lut_tile_5_4_chanxy_out[91];
    assign wire_5825 = lut_tile_5_4_chanxy_out[92];
    assign wire_5827 = lut_tile_5_4_chanxy_out[93];
    assign wire_5829 = lut_tile_5_4_chanxy_out[94];
    assign wire_5831 = lut_tile_5_4_chanxy_out[95];
    assign wire_5833 = lut_tile_5_4_chanxy_out[96];
    assign wire_5835 = lut_tile_5_4_chanxy_out[97];
    assign wire_5837 = lut_tile_5_4_chanxy_out[98];
    assign wire_5839 = lut_tile_5_4_chanxy_out[99];
    assign wire_5840 = lut_tile_5_4_chanxy_out[100];
    assign wire_5841 = lut_tile_5_4_chanxy_out[101];
    assign wire_5842 = lut_tile_5_4_chanxy_out[102];
    assign wire_5843 = lut_tile_5_4_chanxy_out[103];
    assign wire_5844 = lut_tile_5_4_chanxy_out[104];
    assign wire_5845 = lut_tile_5_4_chanxy_out[105];
    assign wire_5846 = lut_tile_5_4_chanxy_out[106];
    assign wire_5847 = lut_tile_5_4_chanxy_out[107];
    assign wire_5848 = lut_tile_5_4_chanxy_out[108];
    assign wire_5849 = lut_tile_5_4_chanxy_out[109];
    assign wire_5850 = lut_tile_5_4_chanxy_out[110];
    assign wire_5851 = lut_tile_5_4_chanxy_out[111];
    assign wire_5852 = lut_tile_5_4_chanxy_out[112];
    assign wire_5853 = lut_tile_5_4_chanxy_out[113];
    assign wire_5854 = lut_tile_5_4_chanxy_out[114];
    assign wire_5855 = lut_tile_5_4_chanxy_out[115];
    assign wire_5856 = lut_tile_5_4_chanxy_out[116];
    assign wire_5857 = lut_tile_5_4_chanxy_out[117];
    assign wire_5858 = lut_tile_5_4_chanxy_out[118];
    assign wire_5859 = lut_tile_5_4_chanxy_out[119];
    assign wire_5860 = lut_tile_5_4_chanxy_out[120];
    assign wire_5861 = lut_tile_5_4_chanxy_out[121];
    assign wire_5862 = lut_tile_5_4_chanxy_out[122];
    assign wire_5863 = lut_tile_5_4_chanxy_out[123];
    assign wire_5864 = lut_tile_5_4_chanxy_out[124];
    assign wire_5865 = lut_tile_5_4_chanxy_out[125];
    assign wire_5866 = lut_tile_5_4_chanxy_out[126];
    assign wire_5867 = lut_tile_5_4_chanxy_out[127];
    assign wire_5868 = lut_tile_5_4_chanxy_out[128];
    assign wire_5869 = lut_tile_5_4_chanxy_out[129];
    assign wire_5870 = lut_tile_5_4_chanxy_out[130];
    assign wire_5871 = lut_tile_5_4_chanxy_out[131];
    assign wire_5872 = lut_tile_5_4_chanxy_out[132];
    assign wire_5873 = lut_tile_5_4_chanxy_out[133];
    assign wire_5874 = lut_tile_5_4_chanxy_out[134];
    assign wire_5875 = lut_tile_5_4_chanxy_out[135];
    assign wire_5876 = lut_tile_5_4_chanxy_out[136];
    assign wire_5877 = lut_tile_5_4_chanxy_out[137];
    assign wire_5878 = lut_tile_5_4_chanxy_out[138];
    assign wire_5879 = lut_tile_5_4_chanxy_out[139];
   // CHANXY OUT
    assign lut_tile_5_5_chanxy_in = {wire_4158, wire_2355, wire_6034, wire_3918, wire_3908, wire_3898, wire_3888, wire_2355, wire_2349, wire_2340, wire_2069, wire_4156, wire_2355, wire_6026, wire_3878, wire_3868, wire_3858, wire_3848, wire_2355, wire_2349, wire_2340, wire_2069, wire_4154, wire_2352, wire_6018, wire_3838, wire_3828, wire_3818, wire_3808, wire_2355, wire_2349, wire_2340, wire_2069, wire_4152, wire_2352, wire_6010, wire_3958, wire_3948, wire_3938, wire_3928, wire_2355, wire_2349, wire_2340, wire_2069, wire_4150, wire_2349, wire_6002, wire_3916, wire_3906, wire_3896, wire_3886, wire_2355, wire_2346, wire_2340, wire_2065, wire_4148, wire_2349, wire_5994, wire_3876, wire_3866, wire_3856, wire_3846, wire_2355, wire_2346, wire_2340, wire_2065, wire_4146, wire_2346, wire_5986, wire_3836, wire_3826, wire_3816, wire_3806, wire_2355, wire_2346, wire_2340, wire_2065, wire_4144, wire_2346, wire_5978, wire_3956, wire_3946, wire_3936, wire_3926, wire_2355, wire_2346, wire_2340, wire_2065, wire_4142, wire_2343, wire_5970, wire_3914, wire_3904, wire_3894, wire_3884, wire_2352, wire_2346, wire_2337, wire_2065, wire_4140, wire_2343, wire_5962, wire_3874, wire_3864, wire_3854, wire_3844, wire_2352, wire_2346, wire_2337, wire_2065, wire_4138, wire_2340, wire_5954, wire_3834, wire_3824, wire_3814, wire_3804, wire_2352, wire_2346, wire_2337, wire_2065, wire_4136, wire_2340, wire_5946, wire_3954, wire_3944, wire_3934, wire_3924, wire_2352, wire_2346, wire_2337, wire_2065, wire_4134, wire_2337, wire_5938, wire_3912, wire_3902, wire_3892, wire_3882, wire_2358, wire_2352, wire_2343, wire_2337, wire_2061, wire_4132, wire_2337, wire_5930, wire_3872, wire_3862, wire_3852, wire_3842, wire_2358, wire_2352, wire_2343, wire_2337, wire_2061, wire_4130, wire_2069, wire_5922, wire_3832, wire_3822, wire_3812, wire_3802, wire_2358, wire_2352, wire_2343, wire_2337, wire_2061, wire_4128, wire_2069, wire_5914, wire_3952, wire_3942, wire_3932, wire_3922, wire_2358, wire_2352, wire_2343, wire_2337, wire_2061, wire_4126, wire_2065, wire_5906, wire_3910, wire_3900, wire_3890, wire_3880, wire_2358, wire_2349, wire_2343, wire_2069, wire_2061, wire_4124, wire_2065, wire_5898, wire_3870, wire_3860, wire_3850, wire_3840, wire_2358, wire_2349, wire_2343, wire_2069, wire_2061, wire_4122, wire_2358, wire_2061, wire_5890, wire_3830, wire_3820, wire_3810, wire_3800, wire_2358, wire_2349, wire_2343, wire_2069, wire_2061, wire_4120, wire_2358, wire_2061, wire_5882, wire_3950, wire_3940, wire_3930, wire_3920, wire_2358, wire_2349, wire_2343, wire_2069, wire_2061, wire_4278, wire_2355, wire_4276, wire_2355, wire_4274, wire_2352, wire_4272, wire_2352, wire_4270, wire_2349, wire_4268, wire_2349, wire_4266, wire_2346, wire_4264, wire_2346, wire_4262, wire_2343, wire_4260, wire_2343, wire_4258, wire_2340, wire_4256, wire_2340, wire_4254, wire_2337, wire_4252, wire_2337, wire_4250, wire_2069, wire_4248, wire_2069, wire_4246, wire_2065, wire_4244, wire_2065, wire_4242, wire_2358, wire_2061, wire_4240, wire_2358, wire_2061, wire_4200, wire_2355, wire_4238, wire_2355, wire_4236, wire_2352, wire_4234, wire_2352, wire_4232, wire_2349, wire_4230, wire_2349, wire_4228, wire_2346, wire_4226, wire_2346, wire_4224, wire_2343, wire_4222, wire_2343, wire_4220, wire_2340, wire_4218, wire_2340, wire_4216, wire_2337, wire_4214, wire_2337, wire_4212, wire_2069, wire_4210, wire_2069, wire_4208, wire_2065, wire_4206, wire_2065, wire_4204, wire_2358, wire_2061, wire_4202, wire_2358, wire_2061, wire_4198, wire_2355, wire_4196, wire_2355, wire_4194, wire_2352, wire_4192, wire_2352, wire_4190, wire_2349, wire_4188, wire_2349, wire_4186, wire_2346, wire_4184, wire_2346, wire_4182, wire_2343, wire_4180, wire_2343, wire_4178, wire_2340, wire_4176, wire_2340, wire_4174, wire_2337, wire_4172, wire_2337, wire_4170, wire_2069, wire_4168, wire_2069, wire_4166, wire_2065, wire_4164, wire_2065, wire_4162, wire_2358, wire_2061, wire_4160, wire_2358, wire_2061, wire_6158, wire_2118, wire_5838, wire_5828, wire_5818, wire_5808, wire_4114, wire_2118, wire_2112, wire_2103, wire_2097, wire_6156, wire_2118, wire_5798, wire_5788, wire_5778, wire_5768, wire_4106, wire_2118, wire_2112, wire_2103, wire_2097, wire_6154, wire_2115, wire_5758, wire_5748, wire_5738, wire_5728, wire_4098, wire_2118, wire_2112, wire_2103, wire_2097, wire_6152, wire_2115, wire_5878, wire_5868, wire_5858, wire_5848, wire_4090, wire_2118, wire_2112, wire_2103, wire_2097, wire_6150, wire_2112, wire_5836, wire_5826, wire_5816, wire_5806, wire_4082, wire_2118, wire_2109, wire_2103, wire_2068, wire_6148, wire_2112, wire_5796, wire_5786, wire_5776, wire_5766, wire_4074, wire_2118, wire_2109, wire_2103, wire_2068, wire_6146, wire_2109, wire_5756, wire_5746, wire_5736, wire_5726, wire_4066, wire_2118, wire_2109, wire_2103, wire_2068, wire_6144, wire_2109, wire_5876, wire_5866, wire_5856, wire_5846, wire_4058, wire_2118, wire_2109, wire_2103, wire_2068, wire_6142, wire_2106, wire_5834, wire_5824, wire_5814, wire_5804, wire_4050, wire_2115, wire_2109, wire_2100, wire_2068, wire_6140, wire_2106, wire_5794, wire_5784, wire_5774, wire_5764, wire_4042, wire_2115, wire_2109, wire_2100, wire_2068, wire_6138, wire_2103, wire_5754, wire_5744, wire_5734, wire_5724, wire_4034, wire_2115, wire_2109, wire_2100, wire_2068, wire_6136, wire_2103, wire_5874, wire_5864, wire_5854, wire_5844, wire_4026, wire_2115, wire_2109, wire_2100, wire_2068, wire_6134, wire_2100, wire_5832, wire_5822, wire_5812, wire_5802, wire_4018, wire_2115, wire_2106, wire_2100, wire_2064, wire_6132, wire_2100, wire_5792, wire_5782, wire_5772, wire_5762, wire_4010, wire_2115, wire_2106, wire_2100, wire_2064, wire_6130, wire_2097, wire_5752, wire_5742, wire_5732, wire_5722, wire_4002, wire_2115, wire_2106, wire_2100, wire_2064, wire_6128, wire_2097, wire_5872, wire_5862, wire_5852, wire_5842, wire_3994, wire_2115, wire_2106, wire_2100, wire_2064, wire_6126, wire_2068, wire_5830, wire_5820, wire_5810, wire_5800, wire_3986, wire_2112, wire_2106, wire_2097, wire_2064, wire_6124, wire_2068, wire_5790, wire_5780, wire_5770, wire_5760, wire_3978, wire_2112, wire_2106, wire_2097, wire_2064, wire_6122, wire_2064, wire_5750, wire_5740, wire_5730, wire_5720, wire_3970, wire_2112, wire_2106, wire_2097, wire_2064, wire_6120, wire_2064, wire_5870, wire_5860, wire_5850, wire_5840, wire_3962, wire_2112, wire_2106, wire_2097, wire_2064, wire_6116, wire_2118, wire_6114, wire_2118, wire_6112, wire_2115, wire_6110, wire_2115, wire_6108, wire_2112, wire_6106, wire_2112, wire_6104, wire_2109, wire_6102, wire_2109, wire_6100, wire_2106, wire_6098, wire_2106, wire_6096, wire_2103, wire_6094, wire_2103, wire_6092, wire_2100, wire_6090, wire_2100, wire_6088, wire_2097, wire_6086, wire_2097, wire_6084, wire_2068, wire_6082, wire_2068, wire_6080, wire_2064, wire_6118, wire_2064, wire_6078, wire_2118, wire_6076, wire_2118, wire_6074, wire_2115, wire_6072, wire_2115, wire_6070, wire_2112, wire_6068, wire_2112, wire_6066, wire_2109, wire_6064, wire_2109, wire_6062, wire_2106, wire_6060, wire_2106, wire_6058, wire_2103, wire_6056, wire_2103, wire_6054, wire_2100, wire_6052, wire_2100, wire_6050, wire_2097, wire_6048, wire_2097, wire_6046, wire_2068, wire_6044, wire_2068, wire_6042, wire_2064, wire_6040, wire_2064, wire_6198, wire_2118, wire_6196, wire_2118, wire_6194, wire_2115, wire_6192, wire_2115, wire_6190, wire_2112, wire_6188, wire_2112, wire_6186, wire_2109, wire_6184, wire_2109, wire_6182, wire_2106, wire_6180, wire_2106, wire_6178, wire_2103, wire_6176, wire_2103, wire_6174, wire_2100, wire_6172, wire_2100, wire_6170, wire_2097, wire_6168, wire_2097, wire_6166, wire_2068, wire_6164, wire_2068, wire_6162, wire_2064, wire_6160, wire_2064};
    // CHNAXY TOTAL: 696
    assign wire_4121 = lut_tile_5_5_chanxy_out[0];
    assign wire_4123 = lut_tile_5_5_chanxy_out[1];
    assign wire_4125 = lut_tile_5_5_chanxy_out[2];
    assign wire_4127 = lut_tile_5_5_chanxy_out[3];
    assign wire_4129 = lut_tile_5_5_chanxy_out[4];
    assign wire_4131 = lut_tile_5_5_chanxy_out[5];
    assign wire_4133 = lut_tile_5_5_chanxy_out[6];
    assign wire_4135 = lut_tile_5_5_chanxy_out[7];
    assign wire_4137 = lut_tile_5_5_chanxy_out[8];
    assign wire_4139 = lut_tile_5_5_chanxy_out[9];
    assign wire_4141 = lut_tile_5_5_chanxy_out[10];
    assign wire_4143 = lut_tile_5_5_chanxy_out[11];
    assign wire_4145 = lut_tile_5_5_chanxy_out[12];
    assign wire_4147 = lut_tile_5_5_chanxy_out[13];
    assign wire_4149 = lut_tile_5_5_chanxy_out[14];
    assign wire_4151 = lut_tile_5_5_chanxy_out[15];
    assign wire_4153 = lut_tile_5_5_chanxy_out[16];
    assign wire_4155 = lut_tile_5_5_chanxy_out[17];
    assign wire_4157 = lut_tile_5_5_chanxy_out[18];
    assign wire_4159 = lut_tile_5_5_chanxy_out[19];
    assign wire_4161 = lut_tile_5_5_chanxy_out[20];
    assign wire_4163 = lut_tile_5_5_chanxy_out[21];
    assign wire_4165 = lut_tile_5_5_chanxy_out[22];
    assign wire_4167 = lut_tile_5_5_chanxy_out[23];
    assign wire_4169 = lut_tile_5_5_chanxy_out[24];
    assign wire_4171 = lut_tile_5_5_chanxy_out[25];
    assign wire_4173 = lut_tile_5_5_chanxy_out[26];
    assign wire_4175 = lut_tile_5_5_chanxy_out[27];
    assign wire_4177 = lut_tile_5_5_chanxy_out[28];
    assign wire_4179 = lut_tile_5_5_chanxy_out[29];
    assign wire_4181 = lut_tile_5_5_chanxy_out[30];
    assign wire_4183 = lut_tile_5_5_chanxy_out[31];
    assign wire_4185 = lut_tile_5_5_chanxy_out[32];
    assign wire_4187 = lut_tile_5_5_chanxy_out[33];
    assign wire_4189 = lut_tile_5_5_chanxy_out[34];
    assign wire_4191 = lut_tile_5_5_chanxy_out[35];
    assign wire_4193 = lut_tile_5_5_chanxy_out[36];
    assign wire_4195 = lut_tile_5_5_chanxy_out[37];
    assign wire_4197 = lut_tile_5_5_chanxy_out[38];
    assign wire_4199 = lut_tile_5_5_chanxy_out[39];
    assign wire_4201 = lut_tile_5_5_chanxy_out[40];
    assign wire_4203 = lut_tile_5_5_chanxy_out[41];
    assign wire_4205 = lut_tile_5_5_chanxy_out[42];
    assign wire_4207 = lut_tile_5_5_chanxy_out[43];
    assign wire_4209 = lut_tile_5_5_chanxy_out[44];
    assign wire_4211 = lut_tile_5_5_chanxy_out[45];
    assign wire_4213 = lut_tile_5_5_chanxy_out[46];
    assign wire_4215 = lut_tile_5_5_chanxy_out[47];
    assign wire_4217 = lut_tile_5_5_chanxy_out[48];
    assign wire_4219 = lut_tile_5_5_chanxy_out[49];
    assign wire_4221 = lut_tile_5_5_chanxy_out[50];
    assign wire_4223 = lut_tile_5_5_chanxy_out[51];
    assign wire_4225 = lut_tile_5_5_chanxy_out[52];
    assign wire_4227 = lut_tile_5_5_chanxy_out[53];
    assign wire_4229 = lut_tile_5_5_chanxy_out[54];
    assign wire_4231 = lut_tile_5_5_chanxy_out[55];
    assign wire_4233 = lut_tile_5_5_chanxy_out[56];
    assign wire_4235 = lut_tile_5_5_chanxy_out[57];
    assign wire_4237 = lut_tile_5_5_chanxy_out[58];
    assign wire_4239 = lut_tile_5_5_chanxy_out[59];
    assign wire_4240 = lut_tile_5_5_chanxy_out[60];
    assign wire_4241 = lut_tile_5_5_chanxy_out[61];
    assign wire_4242 = lut_tile_5_5_chanxy_out[62];
    assign wire_4243 = lut_tile_5_5_chanxy_out[63];
    assign wire_4244 = lut_tile_5_5_chanxy_out[64];
    assign wire_4245 = lut_tile_5_5_chanxy_out[65];
    assign wire_4246 = lut_tile_5_5_chanxy_out[66];
    assign wire_4247 = lut_tile_5_5_chanxy_out[67];
    assign wire_4248 = lut_tile_5_5_chanxy_out[68];
    assign wire_4249 = lut_tile_5_5_chanxy_out[69];
    assign wire_4250 = lut_tile_5_5_chanxy_out[70];
    assign wire_4251 = lut_tile_5_5_chanxy_out[71];
    assign wire_4252 = lut_tile_5_5_chanxy_out[72];
    assign wire_4253 = lut_tile_5_5_chanxy_out[73];
    assign wire_4254 = lut_tile_5_5_chanxy_out[74];
    assign wire_4255 = lut_tile_5_5_chanxy_out[75];
    assign wire_4256 = lut_tile_5_5_chanxy_out[76];
    assign wire_4257 = lut_tile_5_5_chanxy_out[77];
    assign wire_4258 = lut_tile_5_5_chanxy_out[78];
    assign wire_4259 = lut_tile_5_5_chanxy_out[79];
    assign wire_4260 = lut_tile_5_5_chanxy_out[80];
    assign wire_4261 = lut_tile_5_5_chanxy_out[81];
    assign wire_4262 = lut_tile_5_5_chanxy_out[82];
    assign wire_4263 = lut_tile_5_5_chanxy_out[83];
    assign wire_4264 = lut_tile_5_5_chanxy_out[84];
    assign wire_4265 = lut_tile_5_5_chanxy_out[85];
    assign wire_4266 = lut_tile_5_5_chanxy_out[86];
    assign wire_4267 = lut_tile_5_5_chanxy_out[87];
    assign wire_4268 = lut_tile_5_5_chanxy_out[88];
    assign wire_4269 = lut_tile_5_5_chanxy_out[89];
    assign wire_4270 = lut_tile_5_5_chanxy_out[90];
    assign wire_4271 = lut_tile_5_5_chanxy_out[91];
    assign wire_4272 = lut_tile_5_5_chanxy_out[92];
    assign wire_4273 = lut_tile_5_5_chanxy_out[93];
    assign wire_4274 = lut_tile_5_5_chanxy_out[94];
    assign wire_4275 = lut_tile_5_5_chanxy_out[95];
    assign wire_4276 = lut_tile_5_5_chanxy_out[96];
    assign wire_4277 = lut_tile_5_5_chanxy_out[97];
    assign wire_4278 = lut_tile_5_5_chanxy_out[98];
    assign wire_4279 = lut_tile_5_5_chanxy_out[99];
    assign wire_6041 = lut_tile_5_5_chanxy_out[100];
    assign wire_6043 = lut_tile_5_5_chanxy_out[101];
    assign wire_6045 = lut_tile_5_5_chanxy_out[102];
    assign wire_6047 = lut_tile_5_5_chanxy_out[103];
    assign wire_6049 = lut_tile_5_5_chanxy_out[104];
    assign wire_6051 = lut_tile_5_5_chanxy_out[105];
    assign wire_6053 = lut_tile_5_5_chanxy_out[106];
    assign wire_6055 = lut_tile_5_5_chanxy_out[107];
    assign wire_6057 = lut_tile_5_5_chanxy_out[108];
    assign wire_6059 = lut_tile_5_5_chanxy_out[109];
    assign wire_6061 = lut_tile_5_5_chanxy_out[110];
    assign wire_6063 = lut_tile_5_5_chanxy_out[111];
    assign wire_6065 = lut_tile_5_5_chanxy_out[112];
    assign wire_6067 = lut_tile_5_5_chanxy_out[113];
    assign wire_6069 = lut_tile_5_5_chanxy_out[114];
    assign wire_6071 = lut_tile_5_5_chanxy_out[115];
    assign wire_6073 = lut_tile_5_5_chanxy_out[116];
    assign wire_6075 = lut_tile_5_5_chanxy_out[117];
    assign wire_6077 = lut_tile_5_5_chanxy_out[118];
    assign wire_6079 = lut_tile_5_5_chanxy_out[119];
    assign wire_6081 = lut_tile_5_5_chanxy_out[120];
    assign wire_6083 = lut_tile_5_5_chanxy_out[121];
    assign wire_6085 = lut_tile_5_5_chanxy_out[122];
    assign wire_6087 = lut_tile_5_5_chanxy_out[123];
    assign wire_6089 = lut_tile_5_5_chanxy_out[124];
    assign wire_6091 = lut_tile_5_5_chanxy_out[125];
    assign wire_6093 = lut_tile_5_5_chanxy_out[126];
    assign wire_6095 = lut_tile_5_5_chanxy_out[127];
    assign wire_6097 = lut_tile_5_5_chanxy_out[128];
    assign wire_6099 = lut_tile_5_5_chanxy_out[129];
    assign wire_6101 = lut_tile_5_5_chanxy_out[130];
    assign wire_6103 = lut_tile_5_5_chanxy_out[131];
    assign wire_6105 = lut_tile_5_5_chanxy_out[132];
    assign wire_6107 = lut_tile_5_5_chanxy_out[133];
    assign wire_6109 = lut_tile_5_5_chanxy_out[134];
    assign wire_6111 = lut_tile_5_5_chanxy_out[135];
    assign wire_6113 = lut_tile_5_5_chanxy_out[136];
    assign wire_6115 = lut_tile_5_5_chanxy_out[137];
    assign wire_6117 = lut_tile_5_5_chanxy_out[138];
    assign wire_6119 = lut_tile_5_5_chanxy_out[139];
    assign wire_6121 = lut_tile_5_5_chanxy_out[140];
    assign wire_6123 = lut_tile_5_5_chanxy_out[141];
    assign wire_6125 = lut_tile_5_5_chanxy_out[142];
    assign wire_6127 = lut_tile_5_5_chanxy_out[143];
    assign wire_6129 = lut_tile_5_5_chanxy_out[144];
    assign wire_6131 = lut_tile_5_5_chanxy_out[145];
    assign wire_6133 = lut_tile_5_5_chanxy_out[146];
    assign wire_6135 = lut_tile_5_5_chanxy_out[147];
    assign wire_6137 = lut_tile_5_5_chanxy_out[148];
    assign wire_6139 = lut_tile_5_5_chanxy_out[149];
    assign wire_6141 = lut_tile_5_5_chanxy_out[150];
    assign wire_6143 = lut_tile_5_5_chanxy_out[151];
    assign wire_6145 = lut_tile_5_5_chanxy_out[152];
    assign wire_6147 = lut_tile_5_5_chanxy_out[153];
    assign wire_6149 = lut_tile_5_5_chanxy_out[154];
    assign wire_6151 = lut_tile_5_5_chanxy_out[155];
    assign wire_6153 = lut_tile_5_5_chanxy_out[156];
    assign wire_6155 = lut_tile_5_5_chanxy_out[157];
    assign wire_6157 = lut_tile_5_5_chanxy_out[158];
    assign wire_6159 = lut_tile_5_5_chanxy_out[159];
    assign wire_6160 = lut_tile_5_5_chanxy_out[160];
    assign wire_6161 = lut_tile_5_5_chanxy_out[161];
    assign wire_6162 = lut_tile_5_5_chanxy_out[162];
    assign wire_6163 = lut_tile_5_5_chanxy_out[163];
    assign wire_6164 = lut_tile_5_5_chanxy_out[164];
    assign wire_6165 = lut_tile_5_5_chanxy_out[165];
    assign wire_6166 = lut_tile_5_5_chanxy_out[166];
    assign wire_6167 = lut_tile_5_5_chanxy_out[167];
    assign wire_6168 = lut_tile_5_5_chanxy_out[168];
    assign wire_6169 = lut_tile_5_5_chanxy_out[169];
    assign wire_6170 = lut_tile_5_5_chanxy_out[170];
    assign wire_6171 = lut_tile_5_5_chanxy_out[171];
    assign wire_6172 = lut_tile_5_5_chanxy_out[172];
    assign wire_6173 = lut_tile_5_5_chanxy_out[173];
    assign wire_6174 = lut_tile_5_5_chanxy_out[174];
    assign wire_6175 = lut_tile_5_5_chanxy_out[175];
    assign wire_6176 = lut_tile_5_5_chanxy_out[176];
    assign wire_6177 = lut_tile_5_5_chanxy_out[177];
    assign wire_6178 = lut_tile_5_5_chanxy_out[178];
    assign wire_6179 = lut_tile_5_5_chanxy_out[179];
    assign wire_6180 = lut_tile_5_5_chanxy_out[180];
    assign wire_6181 = lut_tile_5_5_chanxy_out[181];
    assign wire_6182 = lut_tile_5_5_chanxy_out[182];
    assign wire_6183 = lut_tile_5_5_chanxy_out[183];
    assign wire_6184 = lut_tile_5_5_chanxy_out[184];
    assign wire_6185 = lut_tile_5_5_chanxy_out[185];
    assign wire_6186 = lut_tile_5_5_chanxy_out[186];
    assign wire_6187 = lut_tile_5_5_chanxy_out[187];
    assign wire_6188 = lut_tile_5_5_chanxy_out[188];
    assign wire_6189 = lut_tile_5_5_chanxy_out[189];
    assign wire_6190 = lut_tile_5_5_chanxy_out[190];
    assign wire_6191 = lut_tile_5_5_chanxy_out[191];
    assign wire_6192 = lut_tile_5_5_chanxy_out[192];
    assign wire_6193 = lut_tile_5_5_chanxy_out[193];
    assign wire_6194 = lut_tile_5_5_chanxy_out[194];
    assign wire_6195 = lut_tile_5_5_chanxy_out[195];
    assign wire_6196 = lut_tile_5_5_chanxy_out[196];
    assign wire_6197 = lut_tile_5_5_chanxy_out[197];
    assign wire_6198 = lut_tile_5_5_chanxy_out[198];
    assign wire_6199 = lut_tile_5_5_chanxy_out[199];
   // CHANXY OUT
    // FPGA IO IPIN
    assign io_tile_1_0_ipin_in = {wire_4439, wire_4438, wire_4419, wire_4418, wire_4399, wire_4398, wire_4379, wire_4378, wire_4359, wire_4358, wire_4339, wire_4338, wire_4319, wire_4318, wire_4299, wire_4298, wire_4435, wire_4434, wire_4415, wire_4414, wire_4395, wire_4394, wire_4375, wire_4374, wire_4355, wire_4354, wire_4335, wire_4334, wire_4315, wire_4314, wire_4295, wire_4294, wire_4433, wire_4432, wire_4413, wire_4412, wire_4393, wire_4392, wire_4373, wire_4372, wire_4353, wire_4352, wire_4333, wire_4332, wire_4313, wire_4312, wire_4293, wire_4292, wire_4431, wire_4430, wire_4411, wire_4410, wire_4391, wire_4390, wire_4371, wire_4370, wire_4351, wire_4350, wire_4331, wire_4330, wire_4311, wire_4310, wire_4291, wire_4290, wire_4429, wire_4428, wire_4409, wire_4408, wire_4389, wire_4388, wire_4369, wire_4368, wire_4349, wire_4348, wire_4329, wire_4328, wire_4309, wire_4308, wire_4289, wire_4288, wire_4425, wire_4424, wire_4405, wire_4404, wire_4385, wire_4384, wire_4365, wire_4364, wire_4345, wire_4344, wire_4325, wire_4324, wire_4305, wire_4304, wire_4285, wire_4284, wire_4423, wire_4422, wire_4403, wire_4402, wire_4383, wire_4382, wire_4363, wire_4362, wire_4343, wire_4342, wire_4323, wire_4322, wire_4303, wire_4302, wire_4283, wire_4282, wire_4421, wire_4420, wire_4401, wire_4400, wire_4381, wire_4380, wire_4361, wire_4360, wire_4341, wire_4340, wire_4321, wire_4320, wire_4301, wire_4300, wire_4281, wire_4280};
    // FPGA IPIN IN
    assign io_tile_2_0_ipin_in = {wire_4437, wire_4436, wire_4417, wire_4416, wire_4397, wire_4396, wire_4377, wire_4376, wire_4357, wire_4356, wire_4337, wire_4336, wire_4317, wire_4316, wire_4297, wire_4296, wire_4433, wire_4432, wire_4413, wire_4412, wire_4393, wire_4392, wire_4373, wire_4372, wire_4353, wire_4352, wire_4333, wire_4332, wire_4313, wire_4312, wire_4293, wire_4292, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_4439, wire_4438, wire_4399, wire_4398, wire_4359, wire_4358, wire_4319, wire_4318, wire_4429, wire_4428, wire_4409, wire_4408, wire_4389, wire_4388, wire_4369, wire_4368, wire_4349, wire_4348, wire_4329, wire_4328, wire_4309, wire_4308, wire_4289, wire_4288, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_4415, wire_4414, wire_4375, wire_4374, wire_4335, wire_4334, wire_4295, wire_4294, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440, wire_4431, wire_4430, wire_4391, wire_4390, wire_4351, wire_4350, wire_4311, wire_4310, wire_4421, wire_4420, wire_4401, wire_4400, wire_4381, wire_4380, wire_4361, wire_4360, wire_4341, wire_4340, wire_4321, wire_4320, wire_4301, wire_4300, wire_4281, wire_4280, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_4407, wire_4406, wire_4367, wire_4366, wire_4327, wire_4326, wire_4287, wire_4286};
    // FPGA IPIN IN
    assign io_tile_3_0_ipin_in = {wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_4423, wire_4422, wire_4383, wire_4382, wire_4343, wire_4342, wire_4303, wire_4302, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_4439, wire_4438, wire_4399, wire_4398, wire_4359, wire_4358, wire_4319, wire_4318, wire_4519, wire_4518, wire_4509, wire_4508, wire_4499, wire_4498, wire_4489, wire_4488, wire_4409, wire_4408, wire_4369, wire_4368, wire_4329, wire_4328, wire_4289, wire_4288, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_4415, wire_4414, wire_4375, wire_4374, wire_4335, wire_4334, wire_4295, wire_4294, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_4425, wire_4424, wire_4385, wire_4384, wire_4345, wire_4344, wire_4305, wire_4304, wire_4517, wire_4516, wire_4507, wire_4506, wire_4497, wire_4496, wire_4487, wire_4486, wire_4401, wire_4400, wire_4361, wire_4360, wire_4321, wire_4320, wire_4281, wire_4280, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_4407, wire_4406, wire_4367, wire_4366, wire_4327, wire_4326, wire_4287, wire_4286, wire_4511, wire_4510, wire_4501, wire_4500, wire_4491, wire_4490, wire_4481, wire_4480, wire_4417, wire_4416, wire_4377, wire_4376, wire_4337, wire_4336, wire_4297, wire_4296};
    // FPGA IPIN IN
    assign io_tile_4_0_ipin_in = {wire_4515, wire_4514, wire_4505, wire_4504, wire_4495, wire_4494, wire_4485, wire_4484, wire_4433, wire_4432, wire_4393, wire_4392, wire_4353, wire_4352, wire_4313, wire_4312, wire_4519, wire_4518, wire_4509, wire_4508, wire_4499, wire_4498, wire_4489, wire_4488, wire_4409, wire_4408, wire_4369, wire_4368, wire_4329, wire_4328, wire_4289, wire_4288, wire_4553, wire_4552, wire_4543, wire_4542, wire_4533, wire_4532, wire_4523, wire_4522, wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_4425, wire_4424, wire_4385, wire_4384, wire_4345, wire_4344, wire_4305, wire_4304, wire_4557, wire_4556, wire_4547, wire_4546, wire_4537, wire_4536, wire_4527, wire_4526, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_4551, wire_4550, wire_4541, wire_4540, wire_4531, wire_4530, wire_4521, wire_4520, wire_4477, wire_4476, wire_4467, wire_4466, wire_4457, wire_4456, wire_4447, wire_4446, wire_4511, wire_4510, wire_4501, wire_4500, wire_4491, wire_4490, wire_4481, wire_4480, wire_4417, wire_4416, wire_4377, wire_4376, wire_4337, wire_4336, wire_4297, wire_4296, wire_4555, wire_4554, wire_4545, wire_4544, wire_4535, wire_4534, wire_4525, wire_4524, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440};
    // FPGA IPIN IN
    assign io_tile_5_0_ipin_in = {wire_4559, wire_4558, wire_4549, wire_4548, wire_4539, wire_4538, wire_4529, wire_4528, wire_4475, wire_4474, wire_4465, wire_4464, wire_4455, wire_4454, wire_4445, wire_4444, wire_4553, wire_4552, wire_4543, wire_4542, wire_4533, wire_4532, wire_4523, wire_4522, wire_4479, wire_4478, wire_4469, wire_4468, wire_4459, wire_4458, wire_4449, wire_4448, wire_4599, wire_4598, wire_4589, wire_4588, wire_4579, wire_4578, wire_4569, wire_4568, wire_4513, wire_4512, wire_4503, wire_4502, wire_4493, wire_4492, wire_4483, wire_4482, wire_4557, wire_4556, wire_4547, wire_4546, wire_4537, wire_4536, wire_4527, wire_4526, wire_4473, wire_4472, wire_4463, wire_4462, wire_4453, wire_4452, wire_4443, wire_4442, wire_4593, wire_4592, wire_4583, wire_4582, wire_4573, wire_4572, wire_4563, wire_4562, wire_4517, wire_4516, wire_4507, wire_4506, wire_4497, wire_4496, wire_4487, wire_4486, wire_4597, wire_4596, wire_4587, wire_4586, wire_4577, wire_4576, wire_4567, wire_4566, wire_4511, wire_4510, wire_4501, wire_4500, wire_4491, wire_4490, wire_4481, wire_4480, wire_4555, wire_4554, wire_4545, wire_4544, wire_4535, wire_4534, wire_4525, wire_4524, wire_4471, wire_4470, wire_4461, wire_4460, wire_4451, wire_4450, wire_4441, wire_4440, wire_4591, wire_4590, wire_4581, wire_4580, wire_4571, wire_4570, wire_4561, wire_4560, wire_4515, wire_4514, wire_4505, wire_4504, wire_4495, wire_4494, wire_4485, wire_4484};
    // FPGA IPIN IN
    assign io_tile_1_6_ipin_in = {wire_6037, wire_6036, wire_6017, wire_6016, wire_5997, wire_5996, wire_5977, wire_5976, wire_5957, wire_5956, wire_5937, wire_5936, wire_5917, wire_5916, wire_5897, wire_5896, wire_6035, wire_6034, wire_6023, wire_6022, wire_5995, wire_5994, wire_5983, wire_5982, wire_5955, wire_5954, wire_5943, wire_5942, wire_5915, wire_5914, wire_5903, wire_5902, wire_6033, wire_6032, wire_6013, wire_6012, wire_5993, wire_5992, wire_5973, wire_5972, wire_5953, wire_5952, wire_5933, wire_5932, wire_5913, wire_5912, wire_5893, wire_5892, wire_6029, wire_6028, wire_6009, wire_6008, wire_5989, wire_5988, wire_5969, wire_5968, wire_5949, wire_5948, wire_5929, wire_5928, wire_5909, wire_5908, wire_5889, wire_5888, wire_6027, wire_6026, wire_6015, wire_6014, wire_5987, wire_5986, wire_5975, wire_5974, wire_5947, wire_5946, wire_5935, wire_5934, wire_5907, wire_5906, wire_5895, wire_5894, wire_6025, wire_6024, wire_6005, wire_6004, wire_5985, wire_5984, wire_5965, wire_5964, wire_5945, wire_5944, wire_5925, wire_5924, wire_5905, wire_5904, wire_5885, wire_5884, wire_6031, wire_6030, wire_6003, wire_6002, wire_5991, wire_5990, wire_5963, wire_5962, wire_5951, wire_5950, wire_5923, wire_5922, wire_5911, wire_5910, wire_5883, wire_5882, wire_6019, wire_6018, wire_6007, wire_6006, wire_5979, wire_5978, wire_5967, wire_5966, wire_5939, wire_5938, wire_5927, wire_5926, wire_5899, wire_5898, wire_5887, wire_5886};
    // FPGA IPIN IN
    assign io_tile_2_6_ipin_in = {wire_6035, wire_6034, wire_6023, wire_6022, wire_5995, wire_5994, wire_5983, wire_5982, wire_5955, wire_5954, wire_5943, wire_5942, wire_5915, wire_5914, wire_5903, wire_5902, wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044, wire_6033, wire_6032, wire_5993, wire_5992, wire_5953, wire_5952, wire_5913, wire_5912, wire_6039, wire_6038, wire_6011, wire_6010, wire_5999, wire_5998, wire_5971, wire_5970, wire_5959, wire_5958, wire_5931, wire_5930, wire_5919, wire_5918, wire_5891, wire_5890, wire_6027, wire_6026, wire_6015, wire_6014, wire_5987, wire_5986, wire_5975, wire_5974, wire_5947, wire_5946, wire_5935, wire_5934, wire_5907, wire_5906, wire_5895, wire_5894, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_6025, wire_6024, wire_5985, wire_5984, wire_5945, wire_5944, wire_5905, wire_5904, wire_6031, wire_6030, wire_6003, wire_6002, wire_5991, wire_5990, wire_5963, wire_5962, wire_5951, wire_5950, wire_5923, wire_5922, wire_5911, wire_5910, wire_5883, wire_5882, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6001, wire_6000, wire_5961, wire_5960, wire_5921, wire_5920, wire_5881, wire_5880, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_6017, wire_6016, wire_5977, wire_5976, wire_5937, wire_5936, wire_5897, wire_5896};
    // FPGA IPIN IN
    assign io_tile_3_6_ipin_in = {wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044, wire_6033, wire_6032, wire_5993, wire_5992, wire_5953, wire_5952, wire_5913, wire_5912, wire_6119, wire_6118, wire_6109, wire_6108, wire_6099, wire_6098, wire_6089, wire_6088, wire_6019, wire_6018, wire_5979, wire_5978, wire_5939, wire_5938, wire_5899, wire_5898, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_6009, wire_6008, wire_5969, wire_5968, wire_5929, wire_5928, wire_5889, wire_5888, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_6025, wire_6024, wire_5985, wire_5984, wire_5945, wire_5944, wire_5905, wire_5904, wire_6117, wire_6116, wire_6107, wire_6106, wire_6097, wire_6096, wire_6087, wire_6086, wire_6011, wire_6010, wire_5971, wire_5970, wire_5931, wire_5930, wire_5891, wire_5890, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6001, wire_6000, wire_5961, wire_5960, wire_5921, wire_5920, wire_5881, wire_5880, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080, wire_6027, wire_6026, wire_5987, wire_5986, wire_5947, wire_5946, wire_5907, wire_5906, wire_6115, wire_6114, wire_6105, wire_6104, wire_6095, wire_6094, wire_6085, wire_6084, wire_6003, wire_6002, wire_5963, wire_5962, wire_5923, wire_5922, wire_5883, wire_5882};
    // FPGA IPIN IN
    assign io_tile_4_6_ipin_in = {wire_6119, wire_6118, wire_6109, wire_6108, wire_6099, wire_6098, wire_6089, wire_6088, wire_6019, wire_6018, wire_5979, wire_5978, wire_5939, wire_5938, wire_5899, wire_5898, wire_6155, wire_6154, wire_6145, wire_6144, wire_6135, wire_6134, wire_6125, wire_6124, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_6113, wire_6112, wire_6103, wire_6102, wire_6093, wire_6092, wire_6083, wire_6082, wire_6035, wire_6034, wire_5995, wire_5994, wire_5955, wire_5954, wire_5915, wire_5914, wire_6117, wire_6116, wire_6107, wire_6106, wire_6097, wire_6096, wire_6087, wire_6086, wire_6011, wire_6010, wire_5971, wire_5970, wire_5931, wire_5930, wire_5891, wire_5890, wire_6153, wire_6152, wire_6143, wire_6142, wire_6133, wire_6132, wire_6123, wire_6122, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080, wire_6027, wire_6026, wire_5987, wire_5986, wire_5947, wire_5946, wire_5907, wire_5906, wire_6157, wire_6156, wire_6147, wire_6146, wire_6137, wire_6136, wire_6127, wire_6126, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_6151, wire_6150, wire_6141, wire_6140, wire_6131, wire_6130, wire_6121, wire_6120, wire_6075, wire_6074, wire_6065, wire_6064, wire_6055, wire_6054, wire_6045, wire_6044};
    // FPGA IPIN IN
    assign io_tile_5_6_ipin_in = {wire_6155, wire_6154, wire_6145, wire_6144, wire_6135, wire_6134, wire_6125, wire_6124, wire_6079, wire_6078, wire_6069, wire_6068, wire_6059, wire_6058, wire_6049, wire_6048, wire_6199, wire_6198, wire_6189, wire_6188, wire_6179, wire_6178, wire_6169, wire_6168, wire_6115, wire_6114, wire_6105, wire_6104, wire_6095, wire_6094, wire_6085, wire_6084, wire_6159, wire_6158, wire_6149, wire_6148, wire_6139, wire_6138, wire_6129, wire_6128, wire_6073, wire_6072, wire_6063, wire_6062, wire_6053, wire_6052, wire_6043, wire_6042, wire_6153, wire_6152, wire_6143, wire_6142, wire_6133, wire_6132, wire_6123, wire_6122, wire_6077, wire_6076, wire_6067, wire_6066, wire_6057, wire_6056, wire_6047, wire_6046, wire_6197, wire_6196, wire_6187, wire_6186, wire_6177, wire_6176, wire_6167, wire_6166, wire_6113, wire_6112, wire_6103, wire_6102, wire_6093, wire_6092, wire_6083, wire_6082, wire_6157, wire_6156, wire_6147, wire_6146, wire_6137, wire_6136, wire_6127, wire_6126, wire_6071, wire_6070, wire_6061, wire_6060, wire_6051, wire_6050, wire_6041, wire_6040, wire_6191, wire_6190, wire_6181, wire_6180, wire_6171, wire_6170, wire_6161, wire_6160, wire_6117, wire_6116, wire_6107, wire_6106, wire_6097, wire_6096, wire_6087, wire_6086, wire_6195, wire_6194, wire_6185, wire_6184, wire_6175, wire_6174, wire_6165, wire_6164, wire_6111, wire_6110, wire_6101, wire_6100, wire_6091, wire_6090, wire_6081, wire_6080};
    // FPGA IPIN IN
    assign io_tile_0_1_ipin_in = {wire_2517, wire_2516, wire_2497, wire_2496, wire_2477, wire_2476, wire_2457, wire_2456, wire_2437, wire_2436, wire_2417, wire_2416, wire_2397, wire_2396, wire_2377, wire_2376, wire_2515, wire_2514, wire_2495, wire_2494, wire_2475, wire_2474, wire_2455, wire_2454, wire_2435, wire_2434, wire_2415, wire_2414, wire_2395, wire_2394, wire_2375, wire_2374, wire_2513, wire_2512, wire_2493, wire_2492, wire_2473, wire_2472, wire_2453, wire_2452, wire_2433, wire_2432, wire_2413, wire_2412, wire_2393, wire_2392, wire_2373, wire_2372, wire_2511, wire_2510, wire_2491, wire_2490, wire_2471, wire_2470, wire_2451, wire_2450, wire_2431, wire_2430, wire_2411, wire_2410, wire_2391, wire_2390, wire_2371, wire_2370, wire_2507, wire_2506, wire_2487, wire_2486, wire_2467, wire_2466, wire_2447, wire_2446, wire_2427, wire_2426, wire_2407, wire_2406, wire_2387, wire_2386, wire_2367, wire_2366, wire_2505, wire_2504, wire_2485, wire_2484, wire_2465, wire_2464, wire_2445, wire_2444, wire_2425, wire_2424, wire_2405, wire_2404, wire_2385, wire_2384, wire_2365, wire_2364, wire_2503, wire_2502, wire_2483, wire_2482, wire_2463, wire_2462, wire_2443, wire_2442, wire_2423, wire_2422, wire_2403, wire_2402, wire_2383, wire_2382, wire_2363, wire_2362, wire_2501, wire_2500, wire_2481, wire_2480, wire_2461, wire_2460, wire_2441, wire_2440, wire_2421, wire_2420, wire_2401, wire_2400, wire_2381, wire_2380, wire_2361, wire_2360};
    // FPGA IPIN IN
    assign io_tile_0_2_ipin_in = {wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_2503, wire_2502, wire_2463, wire_2462, wire_2423, wire_2422, wire_2383, wire_2382, wire_2513, wire_2512, wire_2493, wire_2492, wire_2473, wire_2472, wire_2453, wire_2452, wire_2433, wire_2432, wire_2413, wire_2412, wire_2393, wire_2392, wire_2373, wire_2372, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_2519, wire_2518, wire_2479, wire_2478, wire_2439, wire_2438, wire_2399, wire_2398, wire_2509, wire_2508, wire_2489, wire_2488, wire_2469, wire_2468, wire_2449, wire_2448, wire_2429, wire_2428, wire_2409, wire_2408, wire_2389, wire_2388, wire_2369, wire_2368, wire_2505, wire_2504, wire_2485, wire_2484, wire_2465, wire_2464, wire_2445, wire_2444, wire_2425, wire_2424, wire_2405, wire_2404, wire_2385, wire_2384, wire_2365, wire_2364, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_2511, wire_2510, wire_2471, wire_2470, wire_2431, wire_2430, wire_2391, wire_2390, wire_2501, wire_2500, wire_2481, wire_2480, wire_2461, wire_2460, wire_2441, wire_2440, wire_2421, wire_2420, wire_2401, wire_2400, wire_2381, wire_2380, wire_2361, wire_2360, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_2487, wire_2486, wire_2447, wire_2446, wire_2407, wire_2406, wire_2367, wire_2366};
    // FPGA IPIN IN
    assign io_tile_0_3_ipin_in = {wire_2595, wire_2594, wire_2585, wire_2584, wire_2575, wire_2574, wire_2565, wire_2564, wire_2513, wire_2512, wire_2473, wire_2472, wire_2433, wire_2432, wire_2393, wire_2392, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_2519, wire_2518, wire_2479, wire_2478, wire_2439, wire_2438, wire_2399, wire_2398, wire_2599, wire_2598, wire_2589, wire_2588, wire_2579, wire_2578, wire_2569, wire_2568, wire_2489, wire_2488, wire_2449, wire_2448, wire_2409, wire_2408, wire_2369, wire_2368, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_2495, wire_2494, wire_2455, wire_2454, wire_2415, wire_2414, wire_2375, wire_2374, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_2511, wire_2510, wire_2471, wire_2470, wire_2431, wire_2430, wire_2391, wire_2390, wire_2597, wire_2596, wire_2587, wire_2586, wire_2577, wire_2576, wire_2567, wire_2566, wire_2481, wire_2480, wire_2441, wire_2440, wire_2401, wire_2400, wire_2361, wire_2360, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_2487, wire_2486, wire_2447, wire_2446, wire_2407, wire_2406, wire_2367, wire_2366, wire_2591, wire_2590, wire_2581, wire_2580, wire_2571, wire_2570, wire_2561, wire_2560, wire_2497, wire_2496, wire_2457, wire_2456, wire_2417, wire_2416, wire_2377, wire_2376};
    // FPGA IPIN IN
    assign io_tile_0_4_ipin_in = {wire_2639, wire_2638, wire_2629, wire_2628, wire_2619, wire_2618, wire_2609, wire_2608, wire_2555, wire_2554, wire_2545, wire_2544, wire_2535, wire_2534, wire_2525, wire_2524, wire_2599, wire_2598, wire_2589, wire_2588, wire_2579, wire_2578, wire_2569, wire_2568, wire_2489, wire_2488, wire_2449, wire_2448, wire_2409, wire_2408, wire_2369, wire_2368, wire_2633, wire_2632, wire_2623, wire_2622, wire_2613, wire_2612, wire_2603, wire_2602, wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_2593, wire_2592, wire_2583, wire_2582, wire_2573, wire_2572, wire_2563, wire_2562, wire_2505, wire_2504, wire_2465, wire_2464, wire_2425, wire_2424, wire_2385, wire_2384, wire_2597, wire_2596, wire_2587, wire_2586, wire_2577, wire_2576, wire_2567, wire_2566, wire_2481, wire_2480, wire_2441, wire_2440, wire_2401, wire_2400, wire_2361, wire_2360, wire_2631, wire_2630, wire_2621, wire_2620, wire_2611, wire_2610, wire_2601, wire_2600, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_2591, wire_2590, wire_2581, wire_2580, wire_2571, wire_2570, wire_2561, wire_2560, wire_2497, wire_2496, wire_2457, wire_2456, wire_2417, wire_2416, wire_2377, wire_2376, wire_2635, wire_2634, wire_2625, wire_2624, wire_2615, wire_2614, wire_2605, wire_2604, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520};
    // FPGA IPIN IN
    assign io_tile_0_5_ipin_in = {wire_2675, wire_2674, wire_2665, wire_2664, wire_2655, wire_2654, wire_2645, wire_2644, wire_2599, wire_2598, wire_2589, wire_2588, wire_2579, wire_2578, wire_2569, wire_2568, wire_2633, wire_2632, wire_2623, wire_2622, wire_2613, wire_2612, wire_2603, wire_2602, wire_2559, wire_2558, wire_2549, wire_2548, wire_2539, wire_2538, wire_2529, wire_2528, wire_2679, wire_2678, wire_2669, wire_2668, wire_2659, wire_2658, wire_2649, wire_2648, wire_2593, wire_2592, wire_2583, wire_2582, wire_2573, wire_2572, wire_2563, wire_2562, wire_2637, wire_2636, wire_2627, wire_2626, wire_2617, wire_2616, wire_2607, wire_2606, wire_2553, wire_2552, wire_2543, wire_2542, wire_2533, wire_2532, wire_2523, wire_2522, wire_2631, wire_2630, wire_2621, wire_2620, wire_2611, wire_2610, wire_2601, wire_2600, wire_2557, wire_2556, wire_2547, wire_2546, wire_2537, wire_2536, wire_2527, wire_2526, wire_2677, wire_2676, wire_2667, wire_2666, wire_2657, wire_2656, wire_2647, wire_2646, wire_2591, wire_2590, wire_2581, wire_2580, wire_2571, wire_2570, wire_2561, wire_2560, wire_2635, wire_2634, wire_2625, wire_2624, wire_2615, wire_2614, wire_2605, wire_2604, wire_2551, wire_2550, wire_2541, wire_2540, wire_2531, wire_2530, wire_2521, wire_2520, wire_2671, wire_2670, wire_2661, wire_2660, wire_2651, wire_2650, wire_2641, wire_2640, wire_2595, wire_2594, wire_2585, wire_2584, wire_2575, wire_2574, wire_2565, wire_2564};
    // FPGA IPIN IN
    assign io_tile_6_1_ipin_in = {wire_4117, wire_4116, wire_4097, wire_4096, wire_4077, wire_4076, wire_4057, wire_4056, wire_4037, wire_4036, wire_4017, wire_4016, wire_3997, wire_3996, wire_3977, wire_3976, wire_4115, wire_4114, wire_4103, wire_4102, wire_4075, wire_4074, wire_4063, wire_4062, wire_4035, wire_4034, wire_4023, wire_4022, wire_3995, wire_3994, wire_3983, wire_3982, wire_4119, wire_4118, wire_4091, wire_4090, wire_4079, wire_4078, wire_4051, wire_4050, wire_4039, wire_4038, wire_4011, wire_4010, wire_3999, wire_3998, wire_3971, wire_3970, wire_4109, wire_4108, wire_4089, wire_4088, wire_4069, wire_4068, wire_4049, wire_4048, wire_4029, wire_4028, wire_4009, wire_4008, wire_3989, wire_3988, wire_3969, wire_3968, wire_4107, wire_4106, wire_4095, wire_4094, wire_4067, wire_4066, wire_4055, wire_4054, wire_4027, wire_4026, wire_4015, wire_4014, wire_3987, wire_3986, wire_3975, wire_3974, wire_4105, wire_4104, wire_4085, wire_4084, wire_4065, wire_4064, wire_4045, wire_4044, wire_4025, wire_4024, wire_4005, wire_4004, wire_3985, wire_3984, wire_3965, wire_3964, wire_4101, wire_4100, wire_4081, wire_4080, wire_4061, wire_4060, wire_4041, wire_4040, wire_4021, wire_4020, wire_4001, wire_4000, wire_3981, wire_3980, wire_3961, wire_3960, wire_4099, wire_4098, wire_4087, wire_4086, wire_4059, wire_4058, wire_4047, wire_4046, wire_4019, wire_4018, wire_4007, wire_4006, wire_3979, wire_3978, wire_3967, wire_3966};
    // FPGA IPIN IN
    assign io_tile_6_2_ipin_in = {wire_4115, wire_4114, wire_4103, wire_4102, wire_4075, wire_4074, wire_4063, wire_4062, wire_4035, wire_4034, wire_4023, wire_4022, wire_3995, wire_3994, wire_3983, wire_3982, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_4113, wire_4112, wire_4073, wire_4072, wire_4033, wire_4032, wire_3993, wire_3992, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_4089, wire_4088, wire_4049, wire_4048, wire_4009, wire_4008, wire_3969, wire_3968, wire_4107, wire_4106, wire_4095, wire_4094, wire_4067, wire_4066, wire_4055, wire_4054, wire_4027, wire_4026, wire_4015, wire_4014, wire_3987, wire_3986, wire_3975, wire_3974, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_4105, wire_4104, wire_4065, wire_4064, wire_4025, wire_4024, wire_3985, wire_3984, wire_4111, wire_4110, wire_4083, wire_4082, wire_4071, wire_4070, wire_4043, wire_4042, wire_4031, wire_4030, wire_4003, wire_4002, wire_3991, wire_3990, wire_3963, wire_3962, wire_4099, wire_4098, wire_4087, wire_4086, wire_4059, wire_4058, wire_4047, wire_4046, wire_4019, wire_4018, wire_4007, wire_4006, wire_3979, wire_3978, wire_3967, wire_3966, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_4097, wire_4096, wire_4057, wire_4056, wire_4017, wire_4016, wire_3977, wire_3976};
    // FPGA IPIN IN
    assign io_tile_6_3_ipin_in = {wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_4113, wire_4112, wire_4073, wire_4072, wire_4033, wire_4032, wire_3993, wire_3992, wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_4099, wire_4098, wire_4059, wire_4058, wire_4019, wire_4018, wire_3979, wire_3978, wire_4193, wire_4192, wire_4183, wire_4182, wire_4173, wire_4172, wire_4163, wire_4162, wire_4115, wire_4114, wire_4075, wire_4074, wire_4035, wire_4034, wire_3995, wire_3994, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_4105, wire_4104, wire_4065, wire_4064, wire_4025, wire_4024, wire_3985, wire_3984, wire_4197, wire_4196, wire_4187, wire_4186, wire_4177, wire_4176, wire_4167, wire_4166, wire_4091, wire_4090, wire_4051, wire_4050, wire_4011, wire_4010, wire_3971, wire_3970, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_4081, wire_4080, wire_4041, wire_4040, wire_4001, wire_4000, wire_3961, wire_3960, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_4097, wire_4096, wire_4057, wire_4056, wire_4017, wire_4016, wire_3977, wire_3976, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_4083, wire_4082, wire_4043, wire_4042, wire_4003, wire_4002, wire_3963, wire_3962};
    // FPGA IPIN IN
    assign io_tile_6_4_ipin_in = {wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_4099, wire_4098, wire_4059, wire_4058, wire_4019, wire_4018, wire_3979, wire_3978, wire_4235, wire_4234, wire_4225, wire_4224, wire_4215, wire_4214, wire_4205, wire_4204, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_4239, wire_4238, wire_4229, wire_4228, wire_4219, wire_4218, wire_4209, wire_4208, wire_4153, wire_4152, wire_4143, wire_4142, wire_4133, wire_4132, wire_4123, wire_4122, wire_4197, wire_4196, wire_4187, wire_4186, wire_4177, wire_4176, wire_4167, wire_4166, wire_4091, wire_4090, wire_4051, wire_4050, wire_4011, wire_4010, wire_3971, wire_3970, wire_4233, wire_4232, wire_4223, wire_4222, wire_4213, wire_4212, wire_4203, wire_4202, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_4191, wire_4190, wire_4181, wire_4180, wire_4171, wire_4170, wire_4161, wire_4160, wire_4107, wire_4106, wire_4067, wire_4066, wire_4027, wire_4026, wire_3987, wire_3986, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_4083, wire_4082, wire_4043, wire_4042, wire_4003, wire_4002, wire_3963, wire_3962, wire_4231, wire_4230, wire_4221, wire_4220, wire_4211, wire_4210, wire_4201, wire_4200, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124};
    // FPGA IPIN IN
    assign io_tile_6_5_ipin_in = {wire_4235, wire_4234, wire_4225, wire_4224, wire_4215, wire_4214, wire_4205, wire_4204, wire_4159, wire_4158, wire_4149, wire_4148, wire_4139, wire_4138, wire_4129, wire_4128, wire_4279, wire_4278, wire_4269, wire_4268, wire_4259, wire_4258, wire_4249, wire_4248, wire_4195, wire_4194, wire_4185, wire_4184, wire_4175, wire_4174, wire_4165, wire_4164, wire_4273, wire_4272, wire_4263, wire_4262, wire_4253, wire_4252, wire_4243, wire_4242, wire_4199, wire_4198, wire_4189, wire_4188, wire_4179, wire_4178, wire_4169, wire_4168, wire_4233, wire_4232, wire_4223, wire_4222, wire_4213, wire_4212, wire_4203, wire_4202, wire_4157, wire_4156, wire_4147, wire_4146, wire_4137, wire_4136, wire_4127, wire_4126, wire_4277, wire_4276, wire_4267, wire_4266, wire_4257, wire_4256, wire_4247, wire_4246, wire_4193, wire_4192, wire_4183, wire_4182, wire_4173, wire_4172, wire_4163, wire_4162, wire_4237, wire_4236, wire_4227, wire_4226, wire_4217, wire_4216, wire_4207, wire_4206, wire_4151, wire_4150, wire_4141, wire_4140, wire_4131, wire_4130, wire_4121, wire_4120, wire_4231, wire_4230, wire_4221, wire_4220, wire_4211, wire_4210, wire_4201, wire_4200, wire_4155, wire_4154, wire_4145, wire_4144, wire_4135, wire_4134, wire_4125, wire_4124, wire_4275, wire_4274, wire_4265, wire_4264, wire_4255, wire_4254, wire_4245, wire_4244, wire_4191, wire_4190, wire_4181, wire_4180, wire_4171, wire_4170, wire_4161, wire_4160};
    // FPGA IPIN IN


    // FPGA IO OPIN
    assign wire_25 = io_tile_1_0_opin_out[0];
    assign wire_28 = io_tile_1_0_opin_out[1];
    assign wire_31 = io_tile_1_0_opin_out[2];
    assign wire_34 = io_tile_1_0_opin_out[3];
    assign wire_37 = io_tile_1_0_opin_out[4];
    assign wire_40 = io_tile_1_0_opin_out[5];
    assign wire_43 = io_tile_1_0_opin_out[6];
    assign wire_46 = io_tile_1_0_opin_out[7];
    assign wire_73 = io_tile_2_0_opin_out[0];
    assign wire_76 = io_tile_2_0_opin_out[1];
    assign wire_79 = io_tile_2_0_opin_out[2];
    assign wire_82 = io_tile_2_0_opin_out[3];
    assign wire_85 = io_tile_2_0_opin_out[4];
    assign wire_88 = io_tile_2_0_opin_out[5];
    assign wire_91 = io_tile_2_0_opin_out[6];
    assign wire_94 = io_tile_2_0_opin_out[7];
    assign wire_121 = io_tile_3_0_opin_out[0];
    assign wire_124 = io_tile_3_0_opin_out[1];
    assign wire_127 = io_tile_3_0_opin_out[2];
    assign wire_130 = io_tile_3_0_opin_out[3];
    assign wire_133 = io_tile_3_0_opin_out[4];
    assign wire_136 = io_tile_3_0_opin_out[5];
    assign wire_139 = io_tile_3_0_opin_out[6];
    assign wire_142 = io_tile_3_0_opin_out[7];
    assign wire_169 = io_tile_4_0_opin_out[0];
    assign wire_172 = io_tile_4_0_opin_out[1];
    assign wire_175 = io_tile_4_0_opin_out[2];
    assign wire_178 = io_tile_4_0_opin_out[3];
    assign wire_181 = io_tile_4_0_opin_out[4];
    assign wire_184 = io_tile_4_0_opin_out[5];
    assign wire_187 = io_tile_4_0_opin_out[6];
    assign wire_190 = io_tile_4_0_opin_out[7];
    assign wire_217 = io_tile_5_0_opin_out[0];
    assign wire_220 = io_tile_5_0_opin_out[1];
    assign wire_223 = io_tile_5_0_opin_out[2];
    assign wire_226 = io_tile_5_0_opin_out[3];
    assign wire_229 = io_tile_5_0_opin_out[4];
    assign wire_232 = io_tile_5_0_opin_out[5];
    assign wire_235 = io_tile_5_0_opin_out[6];
    assign wire_238 = io_tile_5_0_opin_out[7];
    assign wire_2145 = io_tile_1_6_opin_out[0];
    assign wire_2148 = io_tile_1_6_opin_out[1];
    assign wire_2151 = io_tile_1_6_opin_out[2];
    assign wire_2154 = io_tile_1_6_opin_out[3];
    assign wire_2157 = io_tile_1_6_opin_out[4];
    assign wire_2160 = io_tile_1_6_opin_out[5];
    assign wire_2163 = io_tile_1_6_opin_out[6];
    assign wire_2166 = io_tile_1_6_opin_out[7];
    assign wire_2193 = io_tile_2_6_opin_out[0];
    assign wire_2196 = io_tile_2_6_opin_out[1];
    assign wire_2199 = io_tile_2_6_opin_out[2];
    assign wire_2202 = io_tile_2_6_opin_out[3];
    assign wire_2205 = io_tile_2_6_opin_out[4];
    assign wire_2208 = io_tile_2_6_opin_out[5];
    assign wire_2211 = io_tile_2_6_opin_out[6];
    assign wire_2214 = io_tile_2_6_opin_out[7];
    assign wire_2241 = io_tile_3_6_opin_out[0];
    assign wire_2244 = io_tile_3_6_opin_out[1];
    assign wire_2247 = io_tile_3_6_opin_out[2];
    assign wire_2250 = io_tile_3_6_opin_out[3];
    assign wire_2253 = io_tile_3_6_opin_out[4];
    assign wire_2256 = io_tile_3_6_opin_out[5];
    assign wire_2259 = io_tile_3_6_opin_out[6];
    assign wire_2262 = io_tile_3_6_opin_out[7];
    assign wire_2289 = io_tile_4_6_opin_out[0];
    assign wire_2292 = io_tile_4_6_opin_out[1];
    assign wire_2295 = io_tile_4_6_opin_out[2];
    assign wire_2298 = io_tile_4_6_opin_out[3];
    assign wire_2301 = io_tile_4_6_opin_out[4];
    assign wire_2304 = io_tile_4_6_opin_out[5];
    assign wire_2307 = io_tile_4_6_opin_out[6];
    assign wire_2310 = io_tile_4_6_opin_out[7];
    assign wire_2337 = io_tile_5_6_opin_out[0];
    assign wire_2340 = io_tile_5_6_opin_out[1];
    assign wire_2343 = io_tile_5_6_opin_out[2];
    assign wire_2346 = io_tile_5_6_opin_out[3];
    assign wire_2349 = io_tile_5_6_opin_out[4];
    assign wire_2352 = io_tile_5_6_opin_out[5];
    assign wire_2355 = io_tile_5_6_opin_out[6];
    assign wire_2358 = io_tile_5_6_opin_out[7];
    assign wire_265 = io_tile_0_1_opin_out[0];
    assign wire_268 = io_tile_0_1_opin_out[1];
    assign wire_271 = io_tile_0_1_opin_out[2];
    assign wire_274 = io_tile_0_1_opin_out[3];
    assign wire_277 = io_tile_0_1_opin_out[4];
    assign wire_280 = io_tile_0_1_opin_out[5];
    assign wire_283 = io_tile_0_1_opin_out[6];
    assign wire_286 = io_tile_0_1_opin_out[7];
    assign wire_641 = io_tile_0_2_opin_out[0];
    assign wire_644 = io_tile_0_2_opin_out[1];
    assign wire_647 = io_tile_0_2_opin_out[2];
    assign wire_650 = io_tile_0_2_opin_out[3];
    assign wire_653 = io_tile_0_2_opin_out[4];
    assign wire_656 = io_tile_0_2_opin_out[5];
    assign wire_659 = io_tile_0_2_opin_out[6];
    assign wire_662 = io_tile_0_2_opin_out[7];
    assign wire_1017 = io_tile_0_3_opin_out[0];
    assign wire_1020 = io_tile_0_3_opin_out[1];
    assign wire_1023 = io_tile_0_3_opin_out[2];
    assign wire_1026 = io_tile_0_3_opin_out[3];
    assign wire_1029 = io_tile_0_3_opin_out[4];
    assign wire_1032 = io_tile_0_3_opin_out[5];
    assign wire_1035 = io_tile_0_3_opin_out[6];
    assign wire_1038 = io_tile_0_3_opin_out[7];
    assign wire_1393 = io_tile_0_4_opin_out[0];
    assign wire_1396 = io_tile_0_4_opin_out[1];
    assign wire_1399 = io_tile_0_4_opin_out[2];
    assign wire_1402 = io_tile_0_4_opin_out[3];
    assign wire_1405 = io_tile_0_4_opin_out[4];
    assign wire_1408 = io_tile_0_4_opin_out[5];
    assign wire_1411 = io_tile_0_4_opin_out[6];
    assign wire_1414 = io_tile_0_4_opin_out[7];
    assign wire_1769 = io_tile_0_5_opin_out[0];
    assign wire_1772 = io_tile_0_5_opin_out[1];
    assign wire_1775 = io_tile_0_5_opin_out[2];
    assign wire_1778 = io_tile_0_5_opin_out[3];
    assign wire_1781 = io_tile_0_5_opin_out[4];
    assign wire_1784 = io_tile_0_5_opin_out[5];
    assign wire_1787 = io_tile_0_5_opin_out[6];
    assign wire_1790 = io_tile_0_5_opin_out[7];
    assign wire_593 = io_tile_6_1_opin_out[0];
    assign wire_596 = io_tile_6_1_opin_out[1];
    assign wire_599 = io_tile_6_1_opin_out[2];
    assign wire_602 = io_tile_6_1_opin_out[3];
    assign wire_605 = io_tile_6_1_opin_out[4];
    assign wire_608 = io_tile_6_1_opin_out[5];
    assign wire_611 = io_tile_6_1_opin_out[6];
    assign wire_614 = io_tile_6_1_opin_out[7];
    assign wire_969 = io_tile_6_2_opin_out[0];
    assign wire_972 = io_tile_6_2_opin_out[1];
    assign wire_975 = io_tile_6_2_opin_out[2];
    assign wire_978 = io_tile_6_2_opin_out[3];
    assign wire_981 = io_tile_6_2_opin_out[4];
    assign wire_984 = io_tile_6_2_opin_out[5];
    assign wire_987 = io_tile_6_2_opin_out[6];
    assign wire_990 = io_tile_6_2_opin_out[7];
    assign wire_1345 = io_tile_6_3_opin_out[0];
    assign wire_1348 = io_tile_6_3_opin_out[1];
    assign wire_1351 = io_tile_6_3_opin_out[2];
    assign wire_1354 = io_tile_6_3_opin_out[3];
    assign wire_1357 = io_tile_6_3_opin_out[4];
    assign wire_1360 = io_tile_6_3_opin_out[5];
    assign wire_1363 = io_tile_6_3_opin_out[6];
    assign wire_1366 = io_tile_6_3_opin_out[7];
    assign wire_1721 = io_tile_6_4_opin_out[0];
    assign wire_1724 = io_tile_6_4_opin_out[1];
    assign wire_1727 = io_tile_6_4_opin_out[2];
    assign wire_1730 = io_tile_6_4_opin_out[3];
    assign wire_1733 = io_tile_6_4_opin_out[4];
    assign wire_1736 = io_tile_6_4_opin_out[5];
    assign wire_1739 = io_tile_6_4_opin_out[6];
    assign wire_1742 = io_tile_6_4_opin_out[7];
    assign wire_2097 = io_tile_6_5_opin_out[0];
    assign wire_2100 = io_tile_6_5_opin_out[1];
    assign wire_2103 = io_tile_6_5_opin_out[2];
    assign wire_2106 = io_tile_6_5_opin_out[3];
    assign wire_2109 = io_tile_6_5_opin_out[4];
    assign wire_2112 = io_tile_6_5_opin_out[5];
    assign wire_2115 = io_tile_6_5_opin_out[6];
    assign wire_2118 = io_tile_6_5_opin_out[7];
    // FPGA IO CHANXY
    assign io_tile_1_0_chanxy_in = {wire_2361, wire_339, wire_2519, wire_339, wire_4479, wire_2839, wire_2799, wire_2759, wire_2719, wire_339, wire_46, wire_37, wire_31, wire_2517, wire_339, wire_2515, wire_339, wire_2513, wire_339, wire_2511, wire_339, wire_4477, wire_2837, wire_2797, wire_2757, wire_2717, wire_339, wire_46, wire_37, wire_31, wire_2509, wire_339, wire_2507, wire_339, wire_2505, wire_335, wire_2503, wire_335, wire_4475, wire_2835, wire_2795, wire_2755, wire_2715, wire_339, wire_46, wire_37, wire_31, wire_2501, wire_335, wire_2499, wire_335, wire_2497, wire_335, wire_2495, wire_335, wire_4473, wire_2833, wire_2793, wire_2753, wire_2713, wire_339, wire_46, wire_37, wire_31, wire_2493, wire_335, wire_2491, wire_335, wire_2489, wire_46, wire_2487, wire_46, wire_4471, wire_2831, wire_2791, wire_2751, wire_2711, wire_339, wire_43, wire_37, wire_28, wire_2485, wire_46, wire_2483, wire_46, wire_2481, wire_46, wire_2479, wire_46, wire_4469, wire_2829, wire_2789, wire_2749, wire_2709, wire_339, wire_43, wire_37, wire_28, wire_2477, wire_46, wire_2475, wire_46, wire_2473, wire_43, wire_2471, wire_43, wire_4467, wire_2827, wire_2787, wire_2747, wire_2707, wire_339, wire_43, wire_37, wire_28, wire_2469, wire_43, wire_2467, wire_43, wire_2465, wire_43, wire_2463, wire_43, wire_4465, wire_2825, wire_2785, wire_2745, wire_2705, wire_339, wire_43, wire_37, wire_28, wire_2461, wire_43, wire_2459, wire_43, wire_2457, wire_40, wire_2455, wire_40, wire_4463, wire_2823, wire_2783, wire_2743, wire_2703, wire_335, wire_43, wire_34, wire_28, wire_2453, wire_40, wire_2451, wire_40, wire_2449, wire_40, wire_2447, wire_40, wire_4461, wire_2821, wire_2781, wire_2741, wire_2701, wire_335, wire_43, wire_34, wire_28, wire_2445, wire_40, wire_2443, wire_40, wire_2441, wire_37, wire_2439, wire_37, wire_4459, wire_2819, wire_2779, wire_2739, wire_2699, wire_335, wire_43, wire_34, wire_28, wire_2437, wire_37, wire_2435, wire_37, wire_2433, wire_37, wire_2431, wire_37, wire_4457, wire_2817, wire_2777, wire_2737, wire_2697, wire_335, wire_43, wire_34, wire_28, wire_2429, wire_37, wire_2427, wire_37, wire_2425, wire_34, wire_2423, wire_34, wire_4455, wire_2815, wire_2775, wire_2735, wire_2695, wire_335, wire_40, wire_34, wire_25, wire_2421, wire_34, wire_2419, wire_34, wire_2417, wire_34, wire_2415, wire_34, wire_4453, wire_2813, wire_2773, wire_2733, wire_2693, wire_335, wire_40, wire_34, wire_25, wire_2413, wire_34, wire_2411, wire_34, wire_2409, wire_31, wire_2407, wire_31, wire_4451, wire_2811, wire_2771, wire_2731, wire_2691, wire_335, wire_40, wire_34, wire_25, wire_2405, wire_31, wire_2403, wire_31, wire_2401, wire_31, wire_2399, wire_31, wire_4449, wire_2809, wire_2769, wire_2729, wire_2689, wire_335, wire_40, wire_34, wire_25, wire_2397, wire_31, wire_2395, wire_31, wire_2393, wire_28, wire_2391, wire_28, wire_4447, wire_2807, wire_2767, wire_2727, wire_2687, wire_46, wire_40, wire_31, wire_25, wire_2389, wire_28, wire_2387, wire_28, wire_2385, wire_28, wire_2383, wire_28, wire_4445, wire_2805, wire_2765, wire_2725, wire_2685, wire_46, wire_40, wire_31, wire_25, wire_2381, wire_28, wire_2379, wire_28, wire_2377, wire_25, wire_2375, wire_25, wire_4443, wire_2803, wire_2763, wire_2723, wire_2683, wire_46, wire_40, wire_31, wire_25, wire_2373, wire_25, wire_2371, wire_25, wire_2369, wire_25, wire_2367, wire_25, wire_4441, wire_2801, wire_2761, wire_2721, wire_2681, wire_46, wire_40, wire_31, wire_25, wire_2365, wire_25, wire_2363, wire_25};
    // CHNAXY TOTAL: 100
    assign wire_4280 = io_tile_1_0_chanxy_out[0];
    assign wire_4282 = io_tile_1_0_chanxy_out[1];
    assign wire_4283 = io_tile_1_0_chanxy_out[2];
    assign wire_4284 = io_tile_1_0_chanxy_out[3];
    assign wire_4286 = io_tile_1_0_chanxy_out[4];
    assign wire_4288 = io_tile_1_0_chanxy_out[5];
    assign wire_4290 = io_tile_1_0_chanxy_out[6];
    assign wire_4291 = io_tile_1_0_chanxy_out[7];
    assign wire_4292 = io_tile_1_0_chanxy_out[8];
    assign wire_4294 = io_tile_1_0_chanxy_out[9];
    assign wire_4296 = io_tile_1_0_chanxy_out[10];
    assign wire_4298 = io_tile_1_0_chanxy_out[11];
    assign wire_4299 = io_tile_1_0_chanxy_out[12];
    assign wire_4300 = io_tile_1_0_chanxy_out[13];
    assign wire_4302 = io_tile_1_0_chanxy_out[14];
    assign wire_4304 = io_tile_1_0_chanxy_out[15];
    assign wire_4306 = io_tile_1_0_chanxy_out[16];
    assign wire_4307 = io_tile_1_0_chanxy_out[17];
    assign wire_4308 = io_tile_1_0_chanxy_out[18];
    assign wire_4310 = io_tile_1_0_chanxy_out[19];
    assign wire_4312 = io_tile_1_0_chanxy_out[20];
    assign wire_4314 = io_tile_1_0_chanxy_out[21];
    assign wire_4315 = io_tile_1_0_chanxy_out[22];
    assign wire_4316 = io_tile_1_0_chanxy_out[23];
    assign wire_4318 = io_tile_1_0_chanxy_out[24];
    assign wire_4320 = io_tile_1_0_chanxy_out[25];
    assign wire_4322 = io_tile_1_0_chanxy_out[26];
    assign wire_4323 = io_tile_1_0_chanxy_out[27];
    assign wire_4324 = io_tile_1_0_chanxy_out[28];
    assign wire_4326 = io_tile_1_0_chanxy_out[29];
    assign wire_4328 = io_tile_1_0_chanxy_out[30];
    assign wire_4330 = io_tile_1_0_chanxy_out[31];
    assign wire_4331 = io_tile_1_0_chanxy_out[32];
    assign wire_4332 = io_tile_1_0_chanxy_out[33];
    assign wire_4334 = io_tile_1_0_chanxy_out[34];
    assign wire_4336 = io_tile_1_0_chanxy_out[35];
    assign wire_4338 = io_tile_1_0_chanxy_out[36];
    assign wire_4339 = io_tile_1_0_chanxy_out[37];
    assign wire_4340 = io_tile_1_0_chanxy_out[38];
    assign wire_4342 = io_tile_1_0_chanxy_out[39];
    assign wire_4344 = io_tile_1_0_chanxy_out[40];
    assign wire_4346 = io_tile_1_0_chanxy_out[41];
    assign wire_4347 = io_tile_1_0_chanxy_out[42];
    assign wire_4348 = io_tile_1_0_chanxy_out[43];
    assign wire_4350 = io_tile_1_0_chanxy_out[44];
    assign wire_4352 = io_tile_1_0_chanxy_out[45];
    assign wire_4354 = io_tile_1_0_chanxy_out[46];
    assign wire_4355 = io_tile_1_0_chanxy_out[47];
    assign wire_4356 = io_tile_1_0_chanxy_out[48];
    assign wire_4358 = io_tile_1_0_chanxy_out[49];
    assign wire_4360 = io_tile_1_0_chanxy_out[50];
    assign wire_4362 = io_tile_1_0_chanxy_out[51];
    assign wire_4363 = io_tile_1_0_chanxy_out[52];
    assign wire_4364 = io_tile_1_0_chanxy_out[53];
    assign wire_4366 = io_tile_1_0_chanxy_out[54];
    assign wire_4368 = io_tile_1_0_chanxy_out[55];
    assign wire_4370 = io_tile_1_0_chanxy_out[56];
    assign wire_4371 = io_tile_1_0_chanxy_out[57];
    assign wire_4372 = io_tile_1_0_chanxy_out[58];
    assign wire_4374 = io_tile_1_0_chanxy_out[59];
    assign wire_4376 = io_tile_1_0_chanxy_out[60];
    assign wire_4378 = io_tile_1_0_chanxy_out[61];
    assign wire_4379 = io_tile_1_0_chanxy_out[62];
    assign wire_4380 = io_tile_1_0_chanxy_out[63];
    assign wire_4382 = io_tile_1_0_chanxy_out[64];
    assign wire_4384 = io_tile_1_0_chanxy_out[65];
    assign wire_4386 = io_tile_1_0_chanxy_out[66];
    assign wire_4387 = io_tile_1_0_chanxy_out[67];
    assign wire_4388 = io_tile_1_0_chanxy_out[68];
    assign wire_4390 = io_tile_1_0_chanxy_out[69];
    assign wire_4392 = io_tile_1_0_chanxy_out[70];
    assign wire_4394 = io_tile_1_0_chanxy_out[71];
    assign wire_4395 = io_tile_1_0_chanxy_out[72];
    assign wire_4396 = io_tile_1_0_chanxy_out[73];
    assign wire_4398 = io_tile_1_0_chanxy_out[74];
    assign wire_4400 = io_tile_1_0_chanxy_out[75];
    assign wire_4402 = io_tile_1_0_chanxy_out[76];
    assign wire_4403 = io_tile_1_0_chanxy_out[77];
    assign wire_4404 = io_tile_1_0_chanxy_out[78];
    assign wire_4406 = io_tile_1_0_chanxy_out[79];
    assign wire_4408 = io_tile_1_0_chanxy_out[80];
    assign wire_4410 = io_tile_1_0_chanxy_out[81];
    assign wire_4411 = io_tile_1_0_chanxy_out[82];
    assign wire_4412 = io_tile_1_0_chanxy_out[83];
    assign wire_4414 = io_tile_1_0_chanxy_out[84];
    assign wire_4416 = io_tile_1_0_chanxy_out[85];
    assign wire_4418 = io_tile_1_0_chanxy_out[86];
    assign wire_4419 = io_tile_1_0_chanxy_out[87];
    assign wire_4420 = io_tile_1_0_chanxy_out[88];
    assign wire_4422 = io_tile_1_0_chanxy_out[89];
    assign wire_4424 = io_tile_1_0_chanxy_out[90];
    assign wire_4426 = io_tile_1_0_chanxy_out[91];
    assign wire_4427 = io_tile_1_0_chanxy_out[92];
    assign wire_4428 = io_tile_1_0_chanxy_out[93];
    assign wire_4430 = io_tile_1_0_chanxy_out[94];
    assign wire_4432 = io_tile_1_0_chanxy_out[95];
    assign wire_4434 = io_tile_1_0_chanxy_out[96];
    assign wire_4435 = io_tile_1_0_chanxy_out[97];
    assign wire_4436 = io_tile_1_0_chanxy_out[98];
    assign wire_4438 = io_tile_1_0_chanxy_out[99];
    assign io_tile_2_0_chanxy_in = {wire_4434, wire_2839, wire_2799, wire_2759, wire_2719, wire_395, wire_94, wire_85, wire_79, wire_4426, wire_2837, wire_2797, wire_2757, wire_2717, wire_395, wire_94, wire_85, wire_79, wire_4418, wire_2835, wire_2795, wire_2755, wire_2715, wire_395, wire_94, wire_85, wire_79, wire_4410, wire_2833, wire_2793, wire_2753, wire_2713, wire_395, wire_94, wire_85, wire_79, wire_4402, wire_2831, wire_2791, wire_2751, wire_2711, wire_395, wire_91, wire_85, wire_76, wire_4394, wire_2829, wire_2789, wire_2749, wire_2709, wire_395, wire_91, wire_85, wire_76, wire_4386, wire_2827, wire_2787, wire_2747, wire_2707, wire_395, wire_91, wire_85, wire_76, wire_4378, wire_2825, wire_2785, wire_2745, wire_2705, wire_395, wire_91, wire_85, wire_76, wire_4370, wire_2823, wire_2783, wire_2743, wire_2703, wire_391, wire_91, wire_82, wire_76, wire_4362, wire_2821, wire_2781, wire_2741, wire_2701, wire_391, wire_91, wire_82, wire_76, wire_4354, wire_2819, wire_2779, wire_2739, wire_2699, wire_391, wire_91, wire_82, wire_76, wire_4346, wire_2817, wire_2777, wire_2737, wire_2697, wire_391, wire_91, wire_82, wire_76, wire_4338, wire_2815, wire_2775, wire_2735, wire_2695, wire_391, wire_88, wire_82, wire_73, wire_4330, wire_2813, wire_2773, wire_2733, wire_2693, wire_391, wire_88, wire_82, wire_73, wire_4322, wire_2811, wire_2771, wire_2731, wire_2691, wire_391, wire_88, wire_82, wire_73, wire_4314, wire_2809, wire_2769, wire_2729, wire_2689, wire_391, wire_88, wire_82, wire_73, wire_4306, wire_2807, wire_2767, wire_2727, wire_2687, wire_94, wire_88, wire_79, wire_73, wire_4298, wire_2805, wire_2765, wire_2725, wire_2685, wire_94, wire_88, wire_79, wire_73, wire_4290, wire_2803, wire_2763, wire_2723, wire_2683, wire_94, wire_88, wire_79, wire_73, wire_4282, wire_2801, wire_2761, wire_2721, wire_2681, wire_94, wire_88, wire_79, wire_73, wire_4519, wire_3159, wire_3119, wire_3079, wire_3039, wire_395, wire_94, wire_85, wire_79, wire_4517, wire_3157, wire_3117, wire_3077, wire_3037, wire_395, wire_94, wire_85, wire_79, wire_4515, wire_3155, wire_3115, wire_3075, wire_3035, wire_395, wire_94, wire_85, wire_79, wire_4513, wire_3153, wire_3113, wire_3073, wire_3033, wire_395, wire_94, wire_85, wire_79, wire_4511, wire_3151, wire_3111, wire_3071, wire_3031, wire_395, wire_91, wire_85, wire_76, wire_4509, wire_3149, wire_3109, wire_3069, wire_3029, wire_395, wire_91, wire_85, wire_76, wire_4507, wire_3147, wire_3107, wire_3067, wire_3027, wire_395, wire_91, wire_85, wire_76, wire_4505, wire_3145, wire_3105, wire_3065, wire_3025, wire_395, wire_91, wire_85, wire_76, wire_4503, wire_3143, wire_3103, wire_3063, wire_3023, wire_391, wire_91, wire_82, wire_76, wire_4501, wire_3141, wire_3101, wire_3061, wire_3021, wire_391, wire_91, wire_82, wire_76, wire_4499, wire_3139, wire_3099, wire_3059, wire_3019, wire_391, wire_91, wire_82, wire_76, wire_4497, wire_3137, wire_3097, wire_3057, wire_3017, wire_391, wire_91, wire_82, wire_76, wire_4495, wire_3135, wire_3095, wire_3055, wire_3015, wire_391, wire_88, wire_82, wire_73, wire_4493, wire_3133, wire_3093, wire_3053, wire_3013, wire_391, wire_88, wire_82, wire_73, wire_4491, wire_3131, wire_3091, wire_3051, wire_3011, wire_391, wire_88, wire_82, wire_73, wire_4489, wire_3129, wire_3089, wire_3049, wire_3009, wire_391, wire_88, wire_82, wire_73, wire_4487, wire_3127, wire_3087, wire_3047, wire_3007, wire_94, wire_88, wire_79, wire_73, wire_4485, wire_3125, wire_3085, wire_3045, wire_3005, wire_94, wire_88, wire_79, wire_73, wire_4483, wire_3123, wire_3083, wire_3043, wire_3003, wire_94, wire_88, wire_79, wire_73, wire_4481, wire_3121, wire_3081, wire_3041, wire_3001, wire_94, wire_88, wire_79, wire_73};
    // CHNAXY TOTAL: 40
    assign wire_4285 = io_tile_2_0_chanxy_out[0];
    assign wire_4293 = io_tile_2_0_chanxy_out[1];
    assign wire_4301 = io_tile_2_0_chanxy_out[2];
    assign wire_4309 = io_tile_2_0_chanxy_out[3];
    assign wire_4317 = io_tile_2_0_chanxy_out[4];
    assign wire_4325 = io_tile_2_0_chanxy_out[5];
    assign wire_4333 = io_tile_2_0_chanxy_out[6];
    assign wire_4341 = io_tile_2_0_chanxy_out[7];
    assign wire_4349 = io_tile_2_0_chanxy_out[8];
    assign wire_4357 = io_tile_2_0_chanxy_out[9];
    assign wire_4365 = io_tile_2_0_chanxy_out[10];
    assign wire_4373 = io_tile_2_0_chanxy_out[11];
    assign wire_4381 = io_tile_2_0_chanxy_out[12];
    assign wire_4389 = io_tile_2_0_chanxy_out[13];
    assign wire_4397 = io_tile_2_0_chanxy_out[14];
    assign wire_4405 = io_tile_2_0_chanxy_out[15];
    assign wire_4413 = io_tile_2_0_chanxy_out[16];
    assign wire_4421 = io_tile_2_0_chanxy_out[17];
    assign wire_4429 = io_tile_2_0_chanxy_out[18];
    assign wire_4437 = io_tile_2_0_chanxy_out[19];
    assign wire_4440 = io_tile_2_0_chanxy_out[20];
    assign wire_4442 = io_tile_2_0_chanxy_out[21];
    assign wire_4444 = io_tile_2_0_chanxy_out[22];
    assign wire_4446 = io_tile_2_0_chanxy_out[23];
    assign wire_4448 = io_tile_2_0_chanxy_out[24];
    assign wire_4450 = io_tile_2_0_chanxy_out[25];
    assign wire_4452 = io_tile_2_0_chanxy_out[26];
    assign wire_4454 = io_tile_2_0_chanxy_out[27];
    assign wire_4456 = io_tile_2_0_chanxy_out[28];
    assign wire_4458 = io_tile_2_0_chanxy_out[29];
    assign wire_4460 = io_tile_2_0_chanxy_out[30];
    assign wire_4462 = io_tile_2_0_chanxy_out[31];
    assign wire_4464 = io_tile_2_0_chanxy_out[32];
    assign wire_4466 = io_tile_2_0_chanxy_out[33];
    assign wire_4468 = io_tile_2_0_chanxy_out[34];
    assign wire_4470 = io_tile_2_0_chanxy_out[35];
    assign wire_4472 = io_tile_2_0_chanxy_out[36];
    assign wire_4474 = io_tile_2_0_chanxy_out[37];
    assign wire_4476 = io_tile_2_0_chanxy_out[38];
    assign wire_4478 = io_tile_2_0_chanxy_out[39];
    assign io_tile_3_0_chanxy_in = {wire_4436, wire_3159, wire_3119, wire_3079, wire_3039, wire_451, wire_142, wire_133, wire_127, wire_4428, wire_3157, wire_3117, wire_3077, wire_3037, wire_451, wire_142, wire_133, wire_127, wire_4420, wire_3155, wire_3115, wire_3075, wire_3035, wire_451, wire_142, wire_133, wire_127, wire_4412, wire_3153, wire_3113, wire_3073, wire_3033, wire_451, wire_142, wire_133, wire_127, wire_4404, wire_3151, wire_3111, wire_3071, wire_3031, wire_451, wire_139, wire_133, wire_124, wire_4396, wire_3149, wire_3109, wire_3069, wire_3029, wire_451, wire_139, wire_133, wire_124, wire_4388, wire_3147, wire_3107, wire_3067, wire_3027, wire_451, wire_139, wire_133, wire_124, wire_4380, wire_3145, wire_3105, wire_3065, wire_3025, wire_451, wire_139, wire_133, wire_124, wire_4372, wire_3143, wire_3103, wire_3063, wire_3023, wire_447, wire_139, wire_130, wire_124, wire_4364, wire_3141, wire_3101, wire_3061, wire_3021, wire_447, wire_139, wire_130, wire_124, wire_4356, wire_3139, wire_3099, wire_3059, wire_3019, wire_447, wire_139, wire_130, wire_124, wire_4348, wire_3137, wire_3097, wire_3057, wire_3017, wire_447, wire_139, wire_130, wire_124, wire_4340, wire_3135, wire_3095, wire_3055, wire_3015, wire_447, wire_136, wire_130, wire_121, wire_4332, wire_3133, wire_3093, wire_3053, wire_3013, wire_447, wire_136, wire_130, wire_121, wire_4324, wire_3131, wire_3091, wire_3051, wire_3011, wire_447, wire_136, wire_130, wire_121, wire_4316, wire_3129, wire_3089, wire_3049, wire_3009, wire_447, wire_136, wire_130, wire_121, wire_4308, wire_3127, wire_3087, wire_3047, wire_3007, wire_142, wire_136, wire_127, wire_121, wire_4300, wire_3125, wire_3085, wire_3045, wire_3005, wire_142, wire_136, wire_127, wire_121, wire_4292, wire_3123, wire_3083, wire_3043, wire_3003, wire_142, wire_136, wire_127, wire_121, wire_4284, wire_3121, wire_3081, wire_3041, wire_3001, wire_142, wire_136, wire_127, wire_121, wire_4559, wire_3479, wire_3439, wire_3399, wire_3359, wire_451, wire_142, wire_133, wire_127, wire_4557, wire_3477, wire_3437, wire_3397, wire_3357, wire_451, wire_142, wire_133, wire_127, wire_4555, wire_3475, wire_3435, wire_3395, wire_3355, wire_451, wire_142, wire_133, wire_127, wire_4553, wire_3473, wire_3433, wire_3393, wire_3353, wire_451, wire_142, wire_133, wire_127, wire_4551, wire_3471, wire_3431, wire_3391, wire_3351, wire_451, wire_139, wire_133, wire_124, wire_4549, wire_3469, wire_3429, wire_3389, wire_3349, wire_451, wire_139, wire_133, wire_124, wire_4547, wire_3467, wire_3427, wire_3387, wire_3347, wire_451, wire_139, wire_133, wire_124, wire_4545, wire_3465, wire_3425, wire_3385, wire_3345, wire_451, wire_139, wire_133, wire_124, wire_4543, wire_3463, wire_3423, wire_3383, wire_3343, wire_447, wire_139, wire_130, wire_124, wire_4541, wire_3461, wire_3421, wire_3381, wire_3341, wire_447, wire_139, wire_130, wire_124, wire_4539, wire_3459, wire_3419, wire_3379, wire_3339, wire_447, wire_139, wire_130, wire_124, wire_4537, wire_3457, wire_3417, wire_3377, wire_3337, wire_447, wire_139, wire_130, wire_124, wire_4535, wire_3455, wire_3415, wire_3375, wire_3335, wire_447, wire_136, wire_130, wire_121, wire_4533, wire_3453, wire_3413, wire_3373, wire_3333, wire_447, wire_136, wire_130, wire_121, wire_4531, wire_3451, wire_3411, wire_3371, wire_3331, wire_447, wire_136, wire_130, wire_121, wire_4529, wire_3449, wire_3409, wire_3369, wire_3329, wire_447, wire_136, wire_130, wire_121, wire_4527, wire_3447, wire_3407, wire_3367, wire_3327, wire_142, wire_136, wire_127, wire_121, wire_4525, wire_3445, wire_3405, wire_3365, wire_3325, wire_142, wire_136, wire_127, wire_121, wire_4523, wire_3443, wire_3403, wire_3363, wire_3323, wire_142, wire_136, wire_127, wire_121, wire_4521, wire_3441, wire_3401, wire_3361, wire_3321, wire_142, wire_136, wire_127, wire_121};
    // CHNAXY TOTAL: 40
    assign wire_4287 = io_tile_3_0_chanxy_out[0];
    assign wire_4295 = io_tile_3_0_chanxy_out[1];
    assign wire_4303 = io_tile_3_0_chanxy_out[2];
    assign wire_4311 = io_tile_3_0_chanxy_out[3];
    assign wire_4319 = io_tile_3_0_chanxy_out[4];
    assign wire_4327 = io_tile_3_0_chanxy_out[5];
    assign wire_4335 = io_tile_3_0_chanxy_out[6];
    assign wire_4343 = io_tile_3_0_chanxy_out[7];
    assign wire_4351 = io_tile_3_0_chanxy_out[8];
    assign wire_4359 = io_tile_3_0_chanxy_out[9];
    assign wire_4367 = io_tile_3_0_chanxy_out[10];
    assign wire_4375 = io_tile_3_0_chanxy_out[11];
    assign wire_4383 = io_tile_3_0_chanxy_out[12];
    assign wire_4391 = io_tile_3_0_chanxy_out[13];
    assign wire_4399 = io_tile_3_0_chanxy_out[14];
    assign wire_4407 = io_tile_3_0_chanxy_out[15];
    assign wire_4415 = io_tile_3_0_chanxy_out[16];
    assign wire_4423 = io_tile_3_0_chanxy_out[17];
    assign wire_4431 = io_tile_3_0_chanxy_out[18];
    assign wire_4439 = io_tile_3_0_chanxy_out[19];
    assign wire_4480 = io_tile_3_0_chanxy_out[20];
    assign wire_4482 = io_tile_3_0_chanxy_out[21];
    assign wire_4484 = io_tile_3_0_chanxy_out[22];
    assign wire_4486 = io_tile_3_0_chanxy_out[23];
    assign wire_4488 = io_tile_3_0_chanxy_out[24];
    assign wire_4490 = io_tile_3_0_chanxy_out[25];
    assign wire_4492 = io_tile_3_0_chanxy_out[26];
    assign wire_4494 = io_tile_3_0_chanxy_out[27];
    assign wire_4496 = io_tile_3_0_chanxy_out[28];
    assign wire_4498 = io_tile_3_0_chanxy_out[29];
    assign wire_4500 = io_tile_3_0_chanxy_out[30];
    assign wire_4502 = io_tile_3_0_chanxy_out[31];
    assign wire_4504 = io_tile_3_0_chanxy_out[32];
    assign wire_4506 = io_tile_3_0_chanxy_out[33];
    assign wire_4508 = io_tile_3_0_chanxy_out[34];
    assign wire_4510 = io_tile_3_0_chanxy_out[35];
    assign wire_4512 = io_tile_3_0_chanxy_out[36];
    assign wire_4514 = io_tile_3_0_chanxy_out[37];
    assign wire_4516 = io_tile_3_0_chanxy_out[38];
    assign wire_4518 = io_tile_3_0_chanxy_out[39];
    assign io_tile_4_0_chanxy_in = {wire_4438, wire_3479, wire_3439, wire_3399, wire_3359, wire_507, wire_190, wire_181, wire_175, wire_4430, wire_3477, wire_3437, wire_3397, wire_3357, wire_507, wire_190, wire_181, wire_175, wire_4422, wire_3475, wire_3435, wire_3395, wire_3355, wire_507, wire_190, wire_181, wire_175, wire_4414, wire_3473, wire_3433, wire_3393, wire_3353, wire_507, wire_190, wire_181, wire_175, wire_4406, wire_3471, wire_3431, wire_3391, wire_3351, wire_507, wire_187, wire_181, wire_172, wire_4398, wire_3469, wire_3429, wire_3389, wire_3349, wire_507, wire_187, wire_181, wire_172, wire_4390, wire_3467, wire_3427, wire_3387, wire_3347, wire_507, wire_187, wire_181, wire_172, wire_4382, wire_3465, wire_3425, wire_3385, wire_3345, wire_507, wire_187, wire_181, wire_172, wire_4374, wire_3463, wire_3423, wire_3383, wire_3343, wire_503, wire_187, wire_178, wire_172, wire_4366, wire_3461, wire_3421, wire_3381, wire_3341, wire_503, wire_187, wire_178, wire_172, wire_4358, wire_3459, wire_3419, wire_3379, wire_3339, wire_503, wire_187, wire_178, wire_172, wire_4350, wire_3457, wire_3417, wire_3377, wire_3337, wire_503, wire_187, wire_178, wire_172, wire_4342, wire_3455, wire_3415, wire_3375, wire_3335, wire_503, wire_184, wire_178, wire_169, wire_4334, wire_3453, wire_3413, wire_3373, wire_3333, wire_503, wire_184, wire_178, wire_169, wire_4326, wire_3451, wire_3411, wire_3371, wire_3331, wire_503, wire_184, wire_178, wire_169, wire_4318, wire_3449, wire_3409, wire_3369, wire_3329, wire_503, wire_184, wire_178, wire_169, wire_4310, wire_3447, wire_3407, wire_3367, wire_3327, wire_190, wire_184, wire_175, wire_169, wire_4302, wire_3445, wire_3405, wire_3365, wire_3325, wire_190, wire_184, wire_175, wire_169, wire_4294, wire_3443, wire_3403, wire_3363, wire_3323, wire_190, wire_184, wire_175, wire_169, wire_4286, wire_3441, wire_3401, wire_3361, wire_3321, wire_190, wire_184, wire_175, wire_169, wire_4599, wire_3799, wire_3759, wire_3719, wire_3679, wire_507, wire_190, wire_181, wire_175, wire_4597, wire_3797, wire_3757, wire_3717, wire_3677, wire_507, wire_190, wire_181, wire_175, wire_4595, wire_3795, wire_3755, wire_3715, wire_3675, wire_507, wire_190, wire_181, wire_175, wire_4593, wire_3793, wire_3753, wire_3713, wire_3673, wire_507, wire_190, wire_181, wire_175, wire_4591, wire_3791, wire_3751, wire_3711, wire_3671, wire_507, wire_187, wire_181, wire_172, wire_4589, wire_3789, wire_3749, wire_3709, wire_3669, wire_507, wire_187, wire_181, wire_172, wire_4587, wire_3787, wire_3747, wire_3707, wire_3667, wire_507, wire_187, wire_181, wire_172, wire_4585, wire_3785, wire_3745, wire_3705, wire_3665, wire_507, wire_187, wire_181, wire_172, wire_4583, wire_3783, wire_3743, wire_3703, wire_3663, wire_503, wire_187, wire_178, wire_172, wire_4581, wire_3781, wire_3741, wire_3701, wire_3661, wire_503, wire_187, wire_178, wire_172, wire_4579, wire_3779, wire_3739, wire_3699, wire_3659, wire_503, wire_187, wire_178, wire_172, wire_4577, wire_3777, wire_3737, wire_3697, wire_3657, wire_503, wire_187, wire_178, wire_172, wire_4575, wire_3775, wire_3735, wire_3695, wire_3655, wire_503, wire_184, wire_178, wire_169, wire_4573, wire_3773, wire_3733, wire_3693, wire_3653, wire_503, wire_184, wire_178, wire_169, wire_4571, wire_3771, wire_3731, wire_3691, wire_3651, wire_503, wire_184, wire_178, wire_169, wire_4569, wire_3769, wire_3729, wire_3689, wire_3649, wire_503, wire_184, wire_178, wire_169, wire_4567, wire_3767, wire_3727, wire_3687, wire_3647, wire_190, wire_184, wire_175, wire_169, wire_4565, wire_3765, wire_3725, wire_3685, wire_3645, wire_190, wire_184, wire_175, wire_169, wire_4563, wire_3763, wire_3723, wire_3683, wire_3643, wire_190, wire_184, wire_175, wire_169, wire_4561, wire_3761, wire_3721, wire_3681, wire_3641, wire_190, wire_184, wire_175, wire_169};
    // CHNAXY TOTAL: 40
    assign wire_4281 = io_tile_4_0_chanxy_out[0];
    assign wire_4289 = io_tile_4_0_chanxy_out[1];
    assign wire_4297 = io_tile_4_0_chanxy_out[2];
    assign wire_4305 = io_tile_4_0_chanxy_out[3];
    assign wire_4313 = io_tile_4_0_chanxy_out[4];
    assign wire_4321 = io_tile_4_0_chanxy_out[5];
    assign wire_4329 = io_tile_4_0_chanxy_out[6];
    assign wire_4337 = io_tile_4_0_chanxy_out[7];
    assign wire_4345 = io_tile_4_0_chanxy_out[8];
    assign wire_4353 = io_tile_4_0_chanxy_out[9];
    assign wire_4361 = io_tile_4_0_chanxy_out[10];
    assign wire_4369 = io_tile_4_0_chanxy_out[11];
    assign wire_4377 = io_tile_4_0_chanxy_out[12];
    assign wire_4385 = io_tile_4_0_chanxy_out[13];
    assign wire_4393 = io_tile_4_0_chanxy_out[14];
    assign wire_4401 = io_tile_4_0_chanxy_out[15];
    assign wire_4409 = io_tile_4_0_chanxy_out[16];
    assign wire_4417 = io_tile_4_0_chanxy_out[17];
    assign wire_4425 = io_tile_4_0_chanxy_out[18];
    assign wire_4433 = io_tile_4_0_chanxy_out[19];
    assign wire_4520 = io_tile_4_0_chanxy_out[20];
    assign wire_4522 = io_tile_4_0_chanxy_out[21];
    assign wire_4524 = io_tile_4_0_chanxy_out[22];
    assign wire_4526 = io_tile_4_0_chanxy_out[23];
    assign wire_4528 = io_tile_4_0_chanxy_out[24];
    assign wire_4530 = io_tile_4_0_chanxy_out[25];
    assign wire_4532 = io_tile_4_0_chanxy_out[26];
    assign wire_4534 = io_tile_4_0_chanxy_out[27];
    assign wire_4536 = io_tile_4_0_chanxy_out[28];
    assign wire_4538 = io_tile_4_0_chanxy_out[29];
    assign wire_4540 = io_tile_4_0_chanxy_out[30];
    assign wire_4542 = io_tile_4_0_chanxy_out[31];
    assign wire_4544 = io_tile_4_0_chanxy_out[32];
    assign wire_4546 = io_tile_4_0_chanxy_out[33];
    assign wire_4548 = io_tile_4_0_chanxy_out[34];
    assign wire_4550 = io_tile_4_0_chanxy_out[35];
    assign wire_4552 = io_tile_4_0_chanxy_out[36];
    assign wire_4554 = io_tile_4_0_chanxy_out[37];
    assign wire_4556 = io_tile_4_0_chanxy_out[38];
    assign wire_4558 = io_tile_4_0_chanxy_out[39];
    assign io_tile_5_0_chanxy_in = {wire_3965, wire_563, wire_4432, wire_3799, wire_3759, wire_3719, wire_3679, wire_563, wire_238, wire_229, wire_223, wire_3973, wire_563, wire_4424, wire_3797, wire_3757, wire_3717, wire_3677, wire_563, wire_238, wire_229, wire_223, wire_3981, wire_559, wire_4416, wire_3795, wire_3755, wire_3715, wire_3675, wire_563, wire_238, wire_229, wire_223, wire_3989, wire_559, wire_4408, wire_3793, wire_3753, wire_3713, wire_3673, wire_563, wire_238, wire_229, wire_223, wire_3997, wire_238, wire_4400, wire_3791, wire_3751, wire_3711, wire_3671, wire_563, wire_235, wire_229, wire_220, wire_4005, wire_238, wire_4392, wire_3789, wire_3749, wire_3709, wire_3669, wire_563, wire_235, wire_229, wire_220, wire_4013, wire_235, wire_4384, wire_3787, wire_3747, wire_3707, wire_3667, wire_563, wire_235, wire_229, wire_220, wire_4021, wire_235, wire_4376, wire_3785, wire_3745, wire_3705, wire_3665, wire_563, wire_235, wire_229, wire_220, wire_4029, wire_232, wire_4368, wire_3783, wire_3743, wire_3703, wire_3663, wire_559, wire_235, wire_226, wire_220, wire_4037, wire_232, wire_4360, wire_3781, wire_3741, wire_3701, wire_3661, wire_559, wire_235, wire_226, wire_220, wire_4045, wire_229, wire_4352, wire_3779, wire_3739, wire_3699, wire_3659, wire_559, wire_235, wire_226, wire_220, wire_4053, wire_229, wire_4344, wire_3777, wire_3737, wire_3697, wire_3657, wire_559, wire_235, wire_226, wire_220, wire_4061, wire_226, wire_4336, wire_3775, wire_3735, wire_3695, wire_3655, wire_559, wire_232, wire_226, wire_217, wire_4069, wire_226, wire_4328, wire_3773, wire_3733, wire_3693, wire_3653, wire_559, wire_232, wire_226, wire_217, wire_4077, wire_223, wire_4320, wire_3771, wire_3731, wire_3691, wire_3651, wire_559, wire_232, wire_226, wire_217, wire_4085, wire_223, wire_4312, wire_3769, wire_3729, wire_3689, wire_3649, wire_559, wire_232, wire_226, wire_217, wire_4093, wire_220, wire_4304, wire_3767, wire_3727, wire_3687, wire_3647, wire_238, wire_232, wire_223, wire_217, wire_4101, wire_220, wire_4296, wire_3765, wire_3725, wire_3685, wire_3645, wire_238, wire_232, wire_223, wire_217, wire_4109, wire_217, wire_4288, wire_3763, wire_3723, wire_3683, wire_3643, wire_238, wire_232, wire_223, wire_217, wire_4117, wire_217, wire_4280, wire_3761, wire_3721, wire_3681, wire_3641, wire_238, wire_232, wire_223, wire_217, wire_4119, wire_563, wire_3967, wire_563, wire_3975, wire_559, wire_3983, wire_559, wire_3991, wire_238, wire_3999, wire_238, wire_4007, wire_235, wire_4015, wire_235, wire_4023, wire_232, wire_4031, wire_232, wire_4039, wire_229, wire_4047, wire_229, wire_4055, wire_226, wire_4063, wire_226, wire_4071, wire_223, wire_4079, wire_223, wire_4087, wire_220, wire_4095, wire_220, wire_4103, wire_217, wire_4111, wire_217, wire_3961, wire_563, wire_3969, wire_563, wire_3977, wire_559, wire_3985, wire_559, wire_3993, wire_238, wire_4001, wire_238, wire_4009, wire_235, wire_4017, wire_235, wire_4025, wire_232, wire_4033, wire_232, wire_4041, wire_229, wire_4049, wire_229, wire_4057, wire_226, wire_4065, wire_226, wire_4073, wire_223, wire_4081, wire_223, wire_4089, wire_220, wire_4097, wire_220, wire_4105, wire_217, wire_4113, wire_217, wire_3963, wire_563, wire_3971, wire_563, wire_3979, wire_559, wire_3987, wire_559, wire_3995, wire_238, wire_4003, wire_238, wire_4011, wire_235, wire_4019, wire_235, wire_4027, wire_232, wire_4035, wire_232, wire_4043, wire_229, wire_4051, wire_229, wire_4059, wire_226, wire_4067, wire_226, wire_4075, wire_223, wire_4083, wire_223, wire_4091, wire_220, wire_4099, wire_220, wire_4107, wire_217, wire_4115, wire_217};
    // CHNAXY TOTAL: 100
    assign wire_4441 = io_tile_5_0_chanxy_out[0];
    assign wire_4443 = io_tile_5_0_chanxy_out[1];
    assign wire_4445 = io_tile_5_0_chanxy_out[2];
    assign wire_4447 = io_tile_5_0_chanxy_out[3];
    assign wire_4449 = io_tile_5_0_chanxy_out[4];
    assign wire_4451 = io_tile_5_0_chanxy_out[5];
    assign wire_4453 = io_tile_5_0_chanxy_out[6];
    assign wire_4455 = io_tile_5_0_chanxy_out[7];
    assign wire_4457 = io_tile_5_0_chanxy_out[8];
    assign wire_4459 = io_tile_5_0_chanxy_out[9];
    assign wire_4461 = io_tile_5_0_chanxy_out[10];
    assign wire_4463 = io_tile_5_0_chanxy_out[11];
    assign wire_4465 = io_tile_5_0_chanxy_out[12];
    assign wire_4467 = io_tile_5_0_chanxy_out[13];
    assign wire_4469 = io_tile_5_0_chanxy_out[14];
    assign wire_4471 = io_tile_5_0_chanxy_out[15];
    assign wire_4473 = io_tile_5_0_chanxy_out[16];
    assign wire_4475 = io_tile_5_0_chanxy_out[17];
    assign wire_4477 = io_tile_5_0_chanxy_out[18];
    assign wire_4479 = io_tile_5_0_chanxy_out[19];
    assign wire_4481 = io_tile_5_0_chanxy_out[20];
    assign wire_4483 = io_tile_5_0_chanxy_out[21];
    assign wire_4485 = io_tile_5_0_chanxy_out[22];
    assign wire_4487 = io_tile_5_0_chanxy_out[23];
    assign wire_4489 = io_tile_5_0_chanxy_out[24];
    assign wire_4491 = io_tile_5_0_chanxy_out[25];
    assign wire_4493 = io_tile_5_0_chanxy_out[26];
    assign wire_4495 = io_tile_5_0_chanxy_out[27];
    assign wire_4497 = io_tile_5_0_chanxy_out[28];
    assign wire_4499 = io_tile_5_0_chanxy_out[29];
    assign wire_4501 = io_tile_5_0_chanxy_out[30];
    assign wire_4503 = io_tile_5_0_chanxy_out[31];
    assign wire_4505 = io_tile_5_0_chanxy_out[32];
    assign wire_4507 = io_tile_5_0_chanxy_out[33];
    assign wire_4509 = io_tile_5_0_chanxy_out[34];
    assign wire_4511 = io_tile_5_0_chanxy_out[35];
    assign wire_4513 = io_tile_5_0_chanxy_out[36];
    assign wire_4515 = io_tile_5_0_chanxy_out[37];
    assign wire_4517 = io_tile_5_0_chanxy_out[38];
    assign wire_4519 = io_tile_5_0_chanxy_out[39];
    assign wire_4521 = io_tile_5_0_chanxy_out[40];
    assign wire_4523 = io_tile_5_0_chanxy_out[41];
    assign wire_4525 = io_tile_5_0_chanxy_out[42];
    assign wire_4527 = io_tile_5_0_chanxy_out[43];
    assign wire_4529 = io_tile_5_0_chanxy_out[44];
    assign wire_4531 = io_tile_5_0_chanxy_out[45];
    assign wire_4533 = io_tile_5_0_chanxy_out[46];
    assign wire_4535 = io_tile_5_0_chanxy_out[47];
    assign wire_4537 = io_tile_5_0_chanxy_out[48];
    assign wire_4539 = io_tile_5_0_chanxy_out[49];
    assign wire_4541 = io_tile_5_0_chanxy_out[50];
    assign wire_4543 = io_tile_5_0_chanxy_out[51];
    assign wire_4545 = io_tile_5_0_chanxy_out[52];
    assign wire_4547 = io_tile_5_0_chanxy_out[53];
    assign wire_4549 = io_tile_5_0_chanxy_out[54];
    assign wire_4551 = io_tile_5_0_chanxy_out[55];
    assign wire_4553 = io_tile_5_0_chanxy_out[56];
    assign wire_4555 = io_tile_5_0_chanxy_out[57];
    assign wire_4557 = io_tile_5_0_chanxy_out[58];
    assign wire_4559 = io_tile_5_0_chanxy_out[59];
    assign wire_4560 = io_tile_5_0_chanxy_out[60];
    assign wire_4561 = io_tile_5_0_chanxy_out[61];
    assign wire_4562 = io_tile_5_0_chanxy_out[62];
    assign wire_4563 = io_tile_5_0_chanxy_out[63];
    assign wire_4564 = io_tile_5_0_chanxy_out[64];
    assign wire_4565 = io_tile_5_0_chanxy_out[65];
    assign wire_4566 = io_tile_5_0_chanxy_out[66];
    assign wire_4567 = io_tile_5_0_chanxy_out[67];
    assign wire_4568 = io_tile_5_0_chanxy_out[68];
    assign wire_4569 = io_tile_5_0_chanxy_out[69];
    assign wire_4570 = io_tile_5_0_chanxy_out[70];
    assign wire_4571 = io_tile_5_0_chanxy_out[71];
    assign wire_4572 = io_tile_5_0_chanxy_out[72];
    assign wire_4573 = io_tile_5_0_chanxy_out[73];
    assign wire_4574 = io_tile_5_0_chanxy_out[74];
    assign wire_4575 = io_tile_5_0_chanxy_out[75];
    assign wire_4576 = io_tile_5_0_chanxy_out[76];
    assign wire_4577 = io_tile_5_0_chanxy_out[77];
    assign wire_4578 = io_tile_5_0_chanxy_out[78];
    assign wire_4579 = io_tile_5_0_chanxy_out[79];
    assign wire_4580 = io_tile_5_0_chanxy_out[80];
    assign wire_4581 = io_tile_5_0_chanxy_out[81];
    assign wire_4582 = io_tile_5_0_chanxy_out[82];
    assign wire_4583 = io_tile_5_0_chanxy_out[83];
    assign wire_4584 = io_tile_5_0_chanxy_out[84];
    assign wire_4585 = io_tile_5_0_chanxy_out[85];
    assign wire_4586 = io_tile_5_0_chanxy_out[86];
    assign wire_4587 = io_tile_5_0_chanxy_out[87];
    assign wire_4588 = io_tile_5_0_chanxy_out[88];
    assign wire_4589 = io_tile_5_0_chanxy_out[89];
    assign wire_4590 = io_tile_5_0_chanxy_out[90];
    assign wire_4591 = io_tile_5_0_chanxy_out[91];
    assign wire_4592 = io_tile_5_0_chanxy_out[92];
    assign wire_4593 = io_tile_5_0_chanxy_out[93];
    assign wire_4594 = io_tile_5_0_chanxy_out[94];
    assign wire_4595 = io_tile_5_0_chanxy_out[95];
    assign wire_4596 = io_tile_5_0_chanxy_out[96];
    assign wire_4597 = io_tile_5_0_chanxy_out[97];
    assign wire_4598 = io_tile_5_0_chanxy_out[98];
    assign wire_4599 = io_tile_5_0_chanxy_out[99];
    assign io_tile_0_1_chanxy_in = {wire_4437, wire_338, wire_4435, wire_338, wire_4759, wire_4719, wire_4679, wire_4639, wire_2559, wire_338, wire_286, wire_277, wire_271, wire_4433, wire_338, wire_4431, wire_338, wire_4429, wire_338, wire_4427, wire_338, wire_4757, wire_4717, wire_4677, wire_4637, wire_2557, wire_338, wire_286, wire_277, wire_271, wire_4425, wire_338, wire_4423, wire_338, wire_4421, wire_334, wire_4419, wire_334, wire_4755, wire_4715, wire_4675, wire_4635, wire_2555, wire_338, wire_286, wire_277, wire_271, wire_4417, wire_334, wire_4415, wire_334, wire_4413, wire_334, wire_4411, wire_334, wire_4753, wire_4713, wire_4673, wire_4633, wire_2553, wire_338, wire_286, wire_277, wire_271, wire_4409, wire_334, wire_4407, wire_334, wire_4405, wire_286, wire_4403, wire_286, wire_4751, wire_4711, wire_4671, wire_4631, wire_2551, wire_338, wire_283, wire_277, wire_268, wire_4401, wire_286, wire_4399, wire_286, wire_4397, wire_286, wire_4395, wire_286, wire_4749, wire_4709, wire_4669, wire_4629, wire_2549, wire_338, wire_283, wire_277, wire_268, wire_4393, wire_286, wire_4391, wire_286, wire_4389, wire_283, wire_4387, wire_283, wire_4747, wire_4707, wire_4667, wire_4627, wire_2547, wire_338, wire_283, wire_277, wire_268, wire_4385, wire_283, wire_4383, wire_283, wire_4381, wire_283, wire_4379, wire_283, wire_4745, wire_4705, wire_4665, wire_4625, wire_2545, wire_338, wire_283, wire_277, wire_268, wire_4377, wire_283, wire_4375, wire_283, wire_4373, wire_280, wire_4371, wire_280, wire_4743, wire_4703, wire_4663, wire_4623, wire_2543, wire_334, wire_283, wire_274, wire_268, wire_4369, wire_280, wire_4367, wire_280, wire_4365, wire_280, wire_4363, wire_280, wire_4741, wire_4701, wire_4661, wire_4621, wire_2541, wire_334, wire_283, wire_274, wire_268, wire_4361, wire_280, wire_4359, wire_280, wire_4357, wire_277, wire_4355, wire_277, wire_4739, wire_4699, wire_4659, wire_4619, wire_2539, wire_334, wire_283, wire_274, wire_268, wire_4353, wire_277, wire_4351, wire_277, wire_4349, wire_277, wire_4347, wire_277, wire_4737, wire_4697, wire_4657, wire_4617, wire_2537, wire_334, wire_283, wire_274, wire_268, wire_4345, wire_277, wire_4343, wire_277, wire_4341, wire_274, wire_4339, wire_274, wire_4735, wire_4695, wire_4655, wire_4615, wire_2535, wire_342, wire_334, wire_280, wire_274, wire_265, wire_4337, wire_274, wire_4335, wire_274, wire_4333, wire_274, wire_4331, wire_274, wire_4733, wire_4693, wire_4653, wire_4613, wire_2533, wire_342, wire_334, wire_280, wire_274, wire_265, wire_4329, wire_274, wire_4327, wire_274, wire_4325, wire_271, wire_4323, wire_271, wire_4731, wire_4691, wire_4651, wire_4611, wire_2531, wire_342, wire_334, wire_280, wire_274, wire_265, wire_4321, wire_271, wire_4319, wire_271, wire_4317, wire_271, wire_4315, wire_271, wire_4729, wire_4689, wire_4649, wire_4609, wire_2529, wire_342, wire_334, wire_280, wire_274, wire_265, wire_4313, wire_271, wire_4311, wire_271, wire_4309, wire_268, wire_4307, wire_268, wire_4727, wire_4687, wire_4647, wire_4607, wire_2527, wire_342, wire_286, wire_280, wire_271, wire_265, wire_4305, wire_268, wire_4303, wire_268, wire_4301, wire_268, wire_4299, wire_268, wire_4725, wire_4685, wire_4645, wire_4605, wire_2525, wire_342, wire_286, wire_280, wire_271, wire_265, wire_4297, wire_268, wire_4295, wire_268, wire_4293, wire_342, wire_265, wire_4291, wire_342, wire_265, wire_4723, wire_4683, wire_4643, wire_4603, wire_2523, wire_342, wire_286, wire_280, wire_271, wire_265, wire_4289, wire_342, wire_265, wire_4287, wire_342, wire_265, wire_4285, wire_342, wire_265, wire_4283, wire_342, wire_265, wire_4721, wire_4681, wire_4641, wire_4601, wire_2521, wire_342, wire_286, wire_280, wire_271, wire_265, wire_4281, wire_342, wire_265, wire_4439, wire_342, wire_265};
    // CHNAXY TOTAL: 100
    assign wire_2360 = io_tile_0_1_chanxy_out[0];
    assign wire_2362 = io_tile_0_1_chanxy_out[1];
    assign wire_2363 = io_tile_0_1_chanxy_out[2];
    assign wire_2364 = io_tile_0_1_chanxy_out[3];
    assign wire_2366 = io_tile_0_1_chanxy_out[4];
    assign wire_2368 = io_tile_0_1_chanxy_out[5];
    assign wire_2370 = io_tile_0_1_chanxy_out[6];
    assign wire_2371 = io_tile_0_1_chanxy_out[7];
    assign wire_2372 = io_tile_0_1_chanxy_out[8];
    assign wire_2374 = io_tile_0_1_chanxy_out[9];
    assign wire_2376 = io_tile_0_1_chanxy_out[10];
    assign wire_2378 = io_tile_0_1_chanxy_out[11];
    assign wire_2379 = io_tile_0_1_chanxy_out[12];
    assign wire_2380 = io_tile_0_1_chanxy_out[13];
    assign wire_2382 = io_tile_0_1_chanxy_out[14];
    assign wire_2384 = io_tile_0_1_chanxy_out[15];
    assign wire_2386 = io_tile_0_1_chanxy_out[16];
    assign wire_2387 = io_tile_0_1_chanxy_out[17];
    assign wire_2388 = io_tile_0_1_chanxy_out[18];
    assign wire_2390 = io_tile_0_1_chanxy_out[19];
    assign wire_2392 = io_tile_0_1_chanxy_out[20];
    assign wire_2394 = io_tile_0_1_chanxy_out[21];
    assign wire_2395 = io_tile_0_1_chanxy_out[22];
    assign wire_2396 = io_tile_0_1_chanxy_out[23];
    assign wire_2398 = io_tile_0_1_chanxy_out[24];
    assign wire_2400 = io_tile_0_1_chanxy_out[25];
    assign wire_2402 = io_tile_0_1_chanxy_out[26];
    assign wire_2403 = io_tile_0_1_chanxy_out[27];
    assign wire_2404 = io_tile_0_1_chanxy_out[28];
    assign wire_2406 = io_tile_0_1_chanxy_out[29];
    assign wire_2408 = io_tile_0_1_chanxy_out[30];
    assign wire_2410 = io_tile_0_1_chanxy_out[31];
    assign wire_2411 = io_tile_0_1_chanxy_out[32];
    assign wire_2412 = io_tile_0_1_chanxy_out[33];
    assign wire_2414 = io_tile_0_1_chanxy_out[34];
    assign wire_2416 = io_tile_0_1_chanxy_out[35];
    assign wire_2418 = io_tile_0_1_chanxy_out[36];
    assign wire_2419 = io_tile_0_1_chanxy_out[37];
    assign wire_2420 = io_tile_0_1_chanxy_out[38];
    assign wire_2422 = io_tile_0_1_chanxy_out[39];
    assign wire_2424 = io_tile_0_1_chanxy_out[40];
    assign wire_2426 = io_tile_0_1_chanxy_out[41];
    assign wire_2427 = io_tile_0_1_chanxy_out[42];
    assign wire_2428 = io_tile_0_1_chanxy_out[43];
    assign wire_2430 = io_tile_0_1_chanxy_out[44];
    assign wire_2432 = io_tile_0_1_chanxy_out[45];
    assign wire_2434 = io_tile_0_1_chanxy_out[46];
    assign wire_2435 = io_tile_0_1_chanxy_out[47];
    assign wire_2436 = io_tile_0_1_chanxy_out[48];
    assign wire_2438 = io_tile_0_1_chanxy_out[49];
    assign wire_2440 = io_tile_0_1_chanxy_out[50];
    assign wire_2442 = io_tile_0_1_chanxy_out[51];
    assign wire_2443 = io_tile_0_1_chanxy_out[52];
    assign wire_2444 = io_tile_0_1_chanxy_out[53];
    assign wire_2446 = io_tile_0_1_chanxy_out[54];
    assign wire_2448 = io_tile_0_1_chanxy_out[55];
    assign wire_2450 = io_tile_0_1_chanxy_out[56];
    assign wire_2451 = io_tile_0_1_chanxy_out[57];
    assign wire_2452 = io_tile_0_1_chanxy_out[58];
    assign wire_2454 = io_tile_0_1_chanxy_out[59];
    assign wire_2456 = io_tile_0_1_chanxy_out[60];
    assign wire_2458 = io_tile_0_1_chanxy_out[61];
    assign wire_2459 = io_tile_0_1_chanxy_out[62];
    assign wire_2460 = io_tile_0_1_chanxy_out[63];
    assign wire_2462 = io_tile_0_1_chanxy_out[64];
    assign wire_2464 = io_tile_0_1_chanxy_out[65];
    assign wire_2466 = io_tile_0_1_chanxy_out[66];
    assign wire_2467 = io_tile_0_1_chanxy_out[67];
    assign wire_2468 = io_tile_0_1_chanxy_out[68];
    assign wire_2470 = io_tile_0_1_chanxy_out[69];
    assign wire_2472 = io_tile_0_1_chanxy_out[70];
    assign wire_2474 = io_tile_0_1_chanxy_out[71];
    assign wire_2475 = io_tile_0_1_chanxy_out[72];
    assign wire_2476 = io_tile_0_1_chanxy_out[73];
    assign wire_2478 = io_tile_0_1_chanxy_out[74];
    assign wire_2480 = io_tile_0_1_chanxy_out[75];
    assign wire_2482 = io_tile_0_1_chanxy_out[76];
    assign wire_2483 = io_tile_0_1_chanxy_out[77];
    assign wire_2484 = io_tile_0_1_chanxy_out[78];
    assign wire_2486 = io_tile_0_1_chanxy_out[79];
    assign wire_2488 = io_tile_0_1_chanxy_out[80];
    assign wire_2490 = io_tile_0_1_chanxy_out[81];
    assign wire_2491 = io_tile_0_1_chanxy_out[82];
    assign wire_2492 = io_tile_0_1_chanxy_out[83];
    assign wire_2494 = io_tile_0_1_chanxy_out[84];
    assign wire_2496 = io_tile_0_1_chanxy_out[85];
    assign wire_2498 = io_tile_0_1_chanxy_out[86];
    assign wire_2499 = io_tile_0_1_chanxy_out[87];
    assign wire_2500 = io_tile_0_1_chanxy_out[88];
    assign wire_2502 = io_tile_0_1_chanxy_out[89];
    assign wire_2504 = io_tile_0_1_chanxy_out[90];
    assign wire_2506 = io_tile_0_1_chanxy_out[91];
    assign wire_2507 = io_tile_0_1_chanxy_out[92];
    assign wire_2508 = io_tile_0_1_chanxy_out[93];
    assign wire_2510 = io_tile_0_1_chanxy_out[94];
    assign wire_2512 = io_tile_0_1_chanxy_out[95];
    assign wire_2514 = io_tile_0_1_chanxy_out[96];
    assign wire_2515 = io_tile_0_1_chanxy_out[97];
    assign wire_2516 = io_tile_0_1_chanxy_out[98];
    assign wire_2518 = io_tile_0_1_chanxy_out[99];
    assign io_tile_0_2_chanxy_in = {wire_4759, wire_4719, wire_4679, wire_4639, wire_2514, wire_714, wire_662, wire_653, wire_647, wire_4757, wire_4717, wire_4677, wire_4637, wire_2506, wire_714, wire_662, wire_653, wire_647, wire_4755, wire_4715, wire_4675, wire_4635, wire_2498, wire_714, wire_662, wire_653, wire_647, wire_4753, wire_4713, wire_4673, wire_4633, wire_2490, wire_714, wire_662, wire_653, wire_647, wire_4751, wire_4711, wire_4671, wire_4631, wire_2482, wire_714, wire_659, wire_653, wire_644, wire_4749, wire_4709, wire_4669, wire_4629, wire_2474, wire_714, wire_659, wire_653, wire_644, wire_4747, wire_4707, wire_4667, wire_4627, wire_2466, wire_714, wire_659, wire_653, wire_644, wire_4745, wire_4705, wire_4665, wire_4625, wire_2458, wire_714, wire_659, wire_653, wire_644, wire_4743, wire_4703, wire_4663, wire_4623, wire_2450, wire_710, wire_659, wire_650, wire_644, wire_4741, wire_4701, wire_4661, wire_4621, wire_2442, wire_710, wire_659, wire_650, wire_644, wire_4739, wire_4699, wire_4659, wire_4619, wire_2434, wire_710, wire_659, wire_650, wire_644, wire_4737, wire_4697, wire_4657, wire_4617, wire_2426, wire_710, wire_659, wire_650, wire_644, wire_4735, wire_4695, wire_4655, wire_4615, wire_2418, wire_718, wire_710, wire_656, wire_650, wire_641, wire_4733, wire_4693, wire_4653, wire_4613, wire_2410, wire_718, wire_710, wire_656, wire_650, wire_641, wire_4731, wire_4691, wire_4651, wire_4611, wire_2402, wire_718, wire_710, wire_656, wire_650, wire_641, wire_4729, wire_4689, wire_4649, wire_4609, wire_2394, wire_718, wire_710, wire_656, wire_650, wire_641, wire_4727, wire_4687, wire_4647, wire_4607, wire_2386, wire_718, wire_662, wire_656, wire_647, wire_641, wire_4725, wire_4685, wire_4645, wire_4605, wire_2378, wire_718, wire_662, wire_656, wire_647, wire_641, wire_4723, wire_4683, wire_4643, wire_4603, wire_2370, wire_718, wire_662, wire_656, wire_647, wire_641, wire_4721, wire_4681, wire_4641, wire_4601, wire_2362, wire_718, wire_662, wire_656, wire_647, wire_641, wire_5079, wire_5039, wire_4999, wire_4959, wire_2599, wire_714, wire_662, wire_653, wire_647, wire_5077, wire_5037, wire_4997, wire_4957, wire_2597, wire_714, wire_662, wire_653, wire_647, wire_5075, wire_5035, wire_4995, wire_4955, wire_2595, wire_714, wire_662, wire_653, wire_647, wire_5073, wire_5033, wire_4993, wire_4953, wire_2593, wire_714, wire_662, wire_653, wire_647, wire_5071, wire_5031, wire_4991, wire_4951, wire_2591, wire_714, wire_659, wire_653, wire_644, wire_5069, wire_5029, wire_4989, wire_4949, wire_2589, wire_714, wire_659, wire_653, wire_644, wire_5067, wire_5027, wire_4987, wire_4947, wire_2587, wire_714, wire_659, wire_653, wire_644, wire_5065, wire_5025, wire_4985, wire_4945, wire_2585, wire_714, wire_659, wire_653, wire_644, wire_5063, wire_5023, wire_4983, wire_4943, wire_2583, wire_710, wire_659, wire_650, wire_644, wire_5061, wire_5021, wire_4981, wire_4941, wire_2581, wire_710, wire_659, wire_650, wire_644, wire_5059, wire_5019, wire_4979, wire_4939, wire_2579, wire_710, wire_659, wire_650, wire_644, wire_5057, wire_5017, wire_4977, wire_4937, wire_2577, wire_710, wire_659, wire_650, wire_644, wire_5055, wire_5015, wire_4975, wire_4935, wire_2575, wire_718, wire_710, wire_656, wire_650, wire_641, wire_5053, wire_5013, wire_4973, wire_4933, wire_2573, wire_718, wire_710, wire_656, wire_650, wire_641, wire_5051, wire_5011, wire_4971, wire_4931, wire_2571, wire_718, wire_710, wire_656, wire_650, wire_641, wire_5049, wire_5009, wire_4969, wire_4929, wire_2569, wire_718, wire_710, wire_656, wire_650, wire_641, wire_5047, wire_5007, wire_4967, wire_4927, wire_2567, wire_718, wire_662, wire_656, wire_647, wire_641, wire_5045, wire_5005, wire_4965, wire_4925, wire_2565, wire_718, wire_662, wire_656, wire_647, wire_641, wire_5043, wire_5003, wire_4963, wire_4923, wire_2563, wire_718, wire_662, wire_656, wire_647, wire_641, wire_5041, wire_5001, wire_4961, wire_4921, wire_2561, wire_718, wire_662, wire_656, wire_647, wire_641};
    // CHNAXY TOTAL: 40
    assign wire_2365 = io_tile_0_2_chanxy_out[0];
    assign wire_2373 = io_tile_0_2_chanxy_out[1];
    assign wire_2381 = io_tile_0_2_chanxy_out[2];
    assign wire_2389 = io_tile_0_2_chanxy_out[3];
    assign wire_2397 = io_tile_0_2_chanxy_out[4];
    assign wire_2405 = io_tile_0_2_chanxy_out[5];
    assign wire_2413 = io_tile_0_2_chanxy_out[6];
    assign wire_2421 = io_tile_0_2_chanxy_out[7];
    assign wire_2429 = io_tile_0_2_chanxy_out[8];
    assign wire_2437 = io_tile_0_2_chanxy_out[9];
    assign wire_2445 = io_tile_0_2_chanxy_out[10];
    assign wire_2453 = io_tile_0_2_chanxy_out[11];
    assign wire_2461 = io_tile_0_2_chanxy_out[12];
    assign wire_2469 = io_tile_0_2_chanxy_out[13];
    assign wire_2477 = io_tile_0_2_chanxy_out[14];
    assign wire_2485 = io_tile_0_2_chanxy_out[15];
    assign wire_2493 = io_tile_0_2_chanxy_out[16];
    assign wire_2501 = io_tile_0_2_chanxy_out[17];
    assign wire_2509 = io_tile_0_2_chanxy_out[18];
    assign wire_2517 = io_tile_0_2_chanxy_out[19];
    assign wire_2520 = io_tile_0_2_chanxy_out[20];
    assign wire_2522 = io_tile_0_2_chanxy_out[21];
    assign wire_2524 = io_tile_0_2_chanxy_out[22];
    assign wire_2526 = io_tile_0_2_chanxy_out[23];
    assign wire_2528 = io_tile_0_2_chanxy_out[24];
    assign wire_2530 = io_tile_0_2_chanxy_out[25];
    assign wire_2532 = io_tile_0_2_chanxy_out[26];
    assign wire_2534 = io_tile_0_2_chanxy_out[27];
    assign wire_2536 = io_tile_0_2_chanxy_out[28];
    assign wire_2538 = io_tile_0_2_chanxy_out[29];
    assign wire_2540 = io_tile_0_2_chanxy_out[30];
    assign wire_2542 = io_tile_0_2_chanxy_out[31];
    assign wire_2544 = io_tile_0_2_chanxy_out[32];
    assign wire_2546 = io_tile_0_2_chanxy_out[33];
    assign wire_2548 = io_tile_0_2_chanxy_out[34];
    assign wire_2550 = io_tile_0_2_chanxy_out[35];
    assign wire_2552 = io_tile_0_2_chanxy_out[36];
    assign wire_2554 = io_tile_0_2_chanxy_out[37];
    assign wire_2556 = io_tile_0_2_chanxy_out[38];
    assign wire_2558 = io_tile_0_2_chanxy_out[39];
    assign io_tile_0_3_chanxy_in = {wire_5079, wire_5039, wire_4999, wire_4959, wire_2516, wire_1090, wire_1038, wire_1029, wire_1023, wire_5077, wire_5037, wire_4997, wire_4957, wire_2508, wire_1090, wire_1038, wire_1029, wire_1023, wire_5075, wire_5035, wire_4995, wire_4955, wire_2500, wire_1090, wire_1038, wire_1029, wire_1023, wire_5073, wire_5033, wire_4993, wire_4953, wire_2492, wire_1090, wire_1038, wire_1029, wire_1023, wire_5071, wire_5031, wire_4991, wire_4951, wire_2484, wire_1090, wire_1035, wire_1029, wire_1020, wire_5069, wire_5029, wire_4989, wire_4949, wire_2476, wire_1090, wire_1035, wire_1029, wire_1020, wire_5067, wire_5027, wire_4987, wire_4947, wire_2468, wire_1090, wire_1035, wire_1029, wire_1020, wire_5065, wire_5025, wire_4985, wire_4945, wire_2460, wire_1090, wire_1035, wire_1029, wire_1020, wire_5063, wire_5023, wire_4983, wire_4943, wire_2452, wire_1086, wire_1035, wire_1026, wire_1020, wire_5061, wire_5021, wire_4981, wire_4941, wire_2444, wire_1086, wire_1035, wire_1026, wire_1020, wire_5059, wire_5019, wire_4979, wire_4939, wire_2436, wire_1086, wire_1035, wire_1026, wire_1020, wire_5057, wire_5017, wire_4977, wire_4937, wire_2428, wire_1086, wire_1035, wire_1026, wire_1020, wire_5055, wire_5015, wire_4975, wire_4935, wire_2420, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5053, wire_5013, wire_4973, wire_4933, wire_2412, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5051, wire_5011, wire_4971, wire_4931, wire_2404, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5049, wire_5009, wire_4969, wire_4929, wire_2396, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5047, wire_5007, wire_4967, wire_4927, wire_2388, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5045, wire_5005, wire_4965, wire_4925, wire_2380, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5043, wire_5003, wire_4963, wire_4923, wire_2372, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5041, wire_5001, wire_4961, wire_4921, wire_2364, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5399, wire_5359, wire_5319, wire_5279, wire_2639, wire_1090, wire_1038, wire_1029, wire_1023, wire_5397, wire_5357, wire_5317, wire_5277, wire_2637, wire_1090, wire_1038, wire_1029, wire_1023, wire_5395, wire_5355, wire_5315, wire_5275, wire_2635, wire_1090, wire_1038, wire_1029, wire_1023, wire_5393, wire_5353, wire_5313, wire_5273, wire_2633, wire_1090, wire_1038, wire_1029, wire_1023, wire_5391, wire_5351, wire_5311, wire_5271, wire_2631, wire_1090, wire_1035, wire_1029, wire_1020, wire_5389, wire_5349, wire_5309, wire_5269, wire_2629, wire_1090, wire_1035, wire_1029, wire_1020, wire_5387, wire_5347, wire_5307, wire_5267, wire_2627, wire_1090, wire_1035, wire_1029, wire_1020, wire_5385, wire_5345, wire_5305, wire_5265, wire_2625, wire_1090, wire_1035, wire_1029, wire_1020, wire_5383, wire_5343, wire_5303, wire_5263, wire_2623, wire_1086, wire_1035, wire_1026, wire_1020, wire_5381, wire_5341, wire_5301, wire_5261, wire_2621, wire_1086, wire_1035, wire_1026, wire_1020, wire_5379, wire_5339, wire_5299, wire_5259, wire_2619, wire_1086, wire_1035, wire_1026, wire_1020, wire_5377, wire_5337, wire_5297, wire_5257, wire_2617, wire_1086, wire_1035, wire_1026, wire_1020, wire_5375, wire_5335, wire_5295, wire_5255, wire_2615, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5373, wire_5333, wire_5293, wire_5253, wire_2613, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5371, wire_5331, wire_5291, wire_5251, wire_2611, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5369, wire_5329, wire_5289, wire_5249, wire_2609, wire_1094, wire_1086, wire_1032, wire_1026, wire_1017, wire_5367, wire_5327, wire_5287, wire_5247, wire_2607, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5365, wire_5325, wire_5285, wire_5245, wire_2605, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5363, wire_5323, wire_5283, wire_5243, wire_2603, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017, wire_5361, wire_5321, wire_5281, wire_5241, wire_2601, wire_1094, wire_1038, wire_1032, wire_1023, wire_1017};
    // CHNAXY TOTAL: 40
    assign wire_2367 = io_tile_0_3_chanxy_out[0];
    assign wire_2375 = io_tile_0_3_chanxy_out[1];
    assign wire_2383 = io_tile_0_3_chanxy_out[2];
    assign wire_2391 = io_tile_0_3_chanxy_out[3];
    assign wire_2399 = io_tile_0_3_chanxy_out[4];
    assign wire_2407 = io_tile_0_3_chanxy_out[5];
    assign wire_2415 = io_tile_0_3_chanxy_out[6];
    assign wire_2423 = io_tile_0_3_chanxy_out[7];
    assign wire_2431 = io_tile_0_3_chanxy_out[8];
    assign wire_2439 = io_tile_0_3_chanxy_out[9];
    assign wire_2447 = io_tile_0_3_chanxy_out[10];
    assign wire_2455 = io_tile_0_3_chanxy_out[11];
    assign wire_2463 = io_tile_0_3_chanxy_out[12];
    assign wire_2471 = io_tile_0_3_chanxy_out[13];
    assign wire_2479 = io_tile_0_3_chanxy_out[14];
    assign wire_2487 = io_tile_0_3_chanxy_out[15];
    assign wire_2495 = io_tile_0_3_chanxy_out[16];
    assign wire_2503 = io_tile_0_3_chanxy_out[17];
    assign wire_2511 = io_tile_0_3_chanxy_out[18];
    assign wire_2519 = io_tile_0_3_chanxy_out[19];
    assign wire_2560 = io_tile_0_3_chanxy_out[20];
    assign wire_2562 = io_tile_0_3_chanxy_out[21];
    assign wire_2564 = io_tile_0_3_chanxy_out[22];
    assign wire_2566 = io_tile_0_3_chanxy_out[23];
    assign wire_2568 = io_tile_0_3_chanxy_out[24];
    assign wire_2570 = io_tile_0_3_chanxy_out[25];
    assign wire_2572 = io_tile_0_3_chanxy_out[26];
    assign wire_2574 = io_tile_0_3_chanxy_out[27];
    assign wire_2576 = io_tile_0_3_chanxy_out[28];
    assign wire_2578 = io_tile_0_3_chanxy_out[29];
    assign wire_2580 = io_tile_0_3_chanxy_out[30];
    assign wire_2582 = io_tile_0_3_chanxy_out[31];
    assign wire_2584 = io_tile_0_3_chanxy_out[32];
    assign wire_2586 = io_tile_0_3_chanxy_out[33];
    assign wire_2588 = io_tile_0_3_chanxy_out[34];
    assign wire_2590 = io_tile_0_3_chanxy_out[35];
    assign wire_2592 = io_tile_0_3_chanxy_out[36];
    assign wire_2594 = io_tile_0_3_chanxy_out[37];
    assign wire_2596 = io_tile_0_3_chanxy_out[38];
    assign wire_2598 = io_tile_0_3_chanxy_out[39];
    assign io_tile_0_4_chanxy_in = {wire_5399, wire_5359, wire_5319, wire_5279, wire_2518, wire_1466, wire_1414, wire_1405, wire_1399, wire_5397, wire_5357, wire_5317, wire_5277, wire_2510, wire_1466, wire_1414, wire_1405, wire_1399, wire_5395, wire_5355, wire_5315, wire_5275, wire_2502, wire_1466, wire_1414, wire_1405, wire_1399, wire_5393, wire_5353, wire_5313, wire_5273, wire_2494, wire_1466, wire_1414, wire_1405, wire_1399, wire_5391, wire_5351, wire_5311, wire_5271, wire_2486, wire_1466, wire_1411, wire_1405, wire_1396, wire_5389, wire_5349, wire_5309, wire_5269, wire_2478, wire_1466, wire_1411, wire_1405, wire_1396, wire_5387, wire_5347, wire_5307, wire_5267, wire_2470, wire_1466, wire_1411, wire_1405, wire_1396, wire_5385, wire_5345, wire_5305, wire_5265, wire_2462, wire_1466, wire_1411, wire_1405, wire_1396, wire_5383, wire_5343, wire_5303, wire_5263, wire_2454, wire_1462, wire_1411, wire_1402, wire_1396, wire_5381, wire_5341, wire_5301, wire_5261, wire_2446, wire_1462, wire_1411, wire_1402, wire_1396, wire_5379, wire_5339, wire_5299, wire_5259, wire_2438, wire_1462, wire_1411, wire_1402, wire_1396, wire_5377, wire_5337, wire_5297, wire_5257, wire_2430, wire_1462, wire_1411, wire_1402, wire_1396, wire_5375, wire_5335, wire_5295, wire_5255, wire_2422, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5373, wire_5333, wire_5293, wire_5253, wire_2414, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5371, wire_5331, wire_5291, wire_5251, wire_2406, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5369, wire_5329, wire_5289, wire_5249, wire_2398, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5367, wire_5327, wire_5287, wire_5247, wire_2390, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5365, wire_5325, wire_5285, wire_5245, wire_2382, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5363, wire_5323, wire_5283, wire_5243, wire_2374, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5361, wire_5321, wire_5281, wire_5241, wire_2366, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5719, wire_5679, wire_5639, wire_5599, wire_2679, wire_1466, wire_1414, wire_1405, wire_1399, wire_5717, wire_5677, wire_5637, wire_5597, wire_2677, wire_1466, wire_1414, wire_1405, wire_1399, wire_5715, wire_5675, wire_5635, wire_5595, wire_2675, wire_1466, wire_1414, wire_1405, wire_1399, wire_5713, wire_5673, wire_5633, wire_5593, wire_2673, wire_1466, wire_1414, wire_1405, wire_1399, wire_5711, wire_5671, wire_5631, wire_5591, wire_2671, wire_1466, wire_1411, wire_1405, wire_1396, wire_5709, wire_5669, wire_5629, wire_5589, wire_2669, wire_1466, wire_1411, wire_1405, wire_1396, wire_5707, wire_5667, wire_5627, wire_5587, wire_2667, wire_1466, wire_1411, wire_1405, wire_1396, wire_5705, wire_5665, wire_5625, wire_5585, wire_2665, wire_1466, wire_1411, wire_1405, wire_1396, wire_5703, wire_5663, wire_5623, wire_5583, wire_2663, wire_1462, wire_1411, wire_1402, wire_1396, wire_5701, wire_5661, wire_5621, wire_5581, wire_2661, wire_1462, wire_1411, wire_1402, wire_1396, wire_5699, wire_5659, wire_5619, wire_5579, wire_2659, wire_1462, wire_1411, wire_1402, wire_1396, wire_5697, wire_5657, wire_5617, wire_5577, wire_2657, wire_1462, wire_1411, wire_1402, wire_1396, wire_5695, wire_5655, wire_5615, wire_5575, wire_2655, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5693, wire_5653, wire_5613, wire_5573, wire_2653, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5691, wire_5651, wire_5611, wire_5571, wire_2651, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5689, wire_5649, wire_5609, wire_5569, wire_2649, wire_1470, wire_1462, wire_1408, wire_1402, wire_1393, wire_5687, wire_5647, wire_5607, wire_5567, wire_2647, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5685, wire_5645, wire_5605, wire_5565, wire_2645, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5683, wire_5643, wire_5603, wire_5563, wire_2643, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393, wire_5681, wire_5641, wire_5601, wire_5561, wire_2641, wire_1470, wire_1414, wire_1408, wire_1399, wire_1393};
    // CHNAXY TOTAL: 40
    assign wire_2361 = io_tile_0_4_chanxy_out[0];
    assign wire_2369 = io_tile_0_4_chanxy_out[1];
    assign wire_2377 = io_tile_0_4_chanxy_out[2];
    assign wire_2385 = io_tile_0_4_chanxy_out[3];
    assign wire_2393 = io_tile_0_4_chanxy_out[4];
    assign wire_2401 = io_tile_0_4_chanxy_out[5];
    assign wire_2409 = io_tile_0_4_chanxy_out[6];
    assign wire_2417 = io_tile_0_4_chanxy_out[7];
    assign wire_2425 = io_tile_0_4_chanxy_out[8];
    assign wire_2433 = io_tile_0_4_chanxy_out[9];
    assign wire_2441 = io_tile_0_4_chanxy_out[10];
    assign wire_2449 = io_tile_0_4_chanxy_out[11];
    assign wire_2457 = io_tile_0_4_chanxy_out[12];
    assign wire_2465 = io_tile_0_4_chanxy_out[13];
    assign wire_2473 = io_tile_0_4_chanxy_out[14];
    assign wire_2481 = io_tile_0_4_chanxy_out[15];
    assign wire_2489 = io_tile_0_4_chanxy_out[16];
    assign wire_2497 = io_tile_0_4_chanxy_out[17];
    assign wire_2505 = io_tile_0_4_chanxy_out[18];
    assign wire_2513 = io_tile_0_4_chanxy_out[19];
    assign wire_2600 = io_tile_0_4_chanxy_out[20];
    assign wire_2602 = io_tile_0_4_chanxy_out[21];
    assign wire_2604 = io_tile_0_4_chanxy_out[22];
    assign wire_2606 = io_tile_0_4_chanxy_out[23];
    assign wire_2608 = io_tile_0_4_chanxy_out[24];
    assign wire_2610 = io_tile_0_4_chanxy_out[25];
    assign wire_2612 = io_tile_0_4_chanxy_out[26];
    assign wire_2614 = io_tile_0_4_chanxy_out[27];
    assign wire_2616 = io_tile_0_4_chanxy_out[28];
    assign wire_2618 = io_tile_0_4_chanxy_out[29];
    assign wire_2620 = io_tile_0_4_chanxy_out[30];
    assign wire_2622 = io_tile_0_4_chanxy_out[31];
    assign wire_2624 = io_tile_0_4_chanxy_out[32];
    assign wire_2626 = io_tile_0_4_chanxy_out[33];
    assign wire_2628 = io_tile_0_4_chanxy_out[34];
    assign wire_2630 = io_tile_0_4_chanxy_out[35];
    assign wire_2632 = io_tile_0_4_chanxy_out[36];
    assign wire_2634 = io_tile_0_4_chanxy_out[37];
    assign wire_2636 = io_tile_0_4_chanxy_out[38];
    assign wire_2638 = io_tile_0_4_chanxy_out[39];
    assign io_tile_0_5_chanxy_in = {wire_5889, wire_1842, wire_5719, wire_5679, wire_5639, wire_5599, wire_2512, wire_1842, wire_1790, wire_1781, wire_1775, wire_5897, wire_1842, wire_5717, wire_5677, wire_5637, wire_5597, wire_2504, wire_1842, wire_1790, wire_1781, wire_1775, wire_5905, wire_1838, wire_5715, wire_5675, wire_5635, wire_5595, wire_2496, wire_1842, wire_1790, wire_1781, wire_1775, wire_5913, wire_1838, wire_5713, wire_5673, wire_5633, wire_5593, wire_2488, wire_1842, wire_1790, wire_1781, wire_1775, wire_5921, wire_1790, wire_5711, wire_5671, wire_5631, wire_5591, wire_2480, wire_1842, wire_1787, wire_1781, wire_1772, wire_5929, wire_1790, wire_5709, wire_5669, wire_5629, wire_5589, wire_2472, wire_1842, wire_1787, wire_1781, wire_1772, wire_5937, wire_1787, wire_5707, wire_5667, wire_5627, wire_5587, wire_2464, wire_1842, wire_1787, wire_1781, wire_1772, wire_5945, wire_1787, wire_5705, wire_5665, wire_5625, wire_5585, wire_2456, wire_1842, wire_1787, wire_1781, wire_1772, wire_5953, wire_1784, wire_5703, wire_5663, wire_5623, wire_5583, wire_2448, wire_1838, wire_1787, wire_1778, wire_1772, wire_5961, wire_1784, wire_5701, wire_5661, wire_5621, wire_5581, wire_2440, wire_1838, wire_1787, wire_1778, wire_1772, wire_5969, wire_1781, wire_5699, wire_5659, wire_5619, wire_5579, wire_2432, wire_1838, wire_1787, wire_1778, wire_1772, wire_5977, wire_1781, wire_5697, wire_5657, wire_5617, wire_5577, wire_2424, wire_1838, wire_1787, wire_1778, wire_1772, wire_5985, wire_1778, wire_5695, wire_5655, wire_5615, wire_5575, wire_2416, wire_1846, wire_1838, wire_1784, wire_1778, wire_1769, wire_5993, wire_1778, wire_5693, wire_5653, wire_5613, wire_5573, wire_2408, wire_1846, wire_1838, wire_1784, wire_1778, wire_1769, wire_6001, wire_1775, wire_5691, wire_5651, wire_5611, wire_5571, wire_2400, wire_1846, wire_1838, wire_1784, wire_1778, wire_1769, wire_6009, wire_1775, wire_5689, wire_5649, wire_5609, wire_5569, wire_2392, wire_1846, wire_1838, wire_1784, wire_1778, wire_1769, wire_6017, wire_1772, wire_5687, wire_5647, wire_5607, wire_5567, wire_2384, wire_1846, wire_1790, wire_1784, wire_1775, wire_1769, wire_6025, wire_1772, wire_5685, wire_5645, wire_5605, wire_5565, wire_2376, wire_1846, wire_1790, wire_1784, wire_1775, wire_1769, wire_6033, wire_1846, wire_1769, wire_5683, wire_5643, wire_5603, wire_5563, wire_2368, wire_1846, wire_1790, wire_1784, wire_1775, wire_1769, wire_5881, wire_1846, wire_1769, wire_5681, wire_5641, wire_5601, wire_5561, wire_2360, wire_1846, wire_1790, wire_1784, wire_1775, wire_1769, wire_5883, wire_1842, wire_5891, wire_1842, wire_5899, wire_1838, wire_5907, wire_1838, wire_5915, wire_1790, wire_5923, wire_1790, wire_5931, wire_1787, wire_5939, wire_1787, wire_5947, wire_1784, wire_5955, wire_1784, wire_5963, wire_1781, wire_5971, wire_1781, wire_5979, wire_1778, wire_5987, wire_1778, wire_5995, wire_1775, wire_6003, wire_1775, wire_6011, wire_1772, wire_6019, wire_1772, wire_6027, wire_1846, wire_1769, wire_6035, wire_1846, wire_1769, wire_5885, wire_1842, wire_5893, wire_1842, wire_5901, wire_1838, wire_5909, wire_1838, wire_5917, wire_1790, wire_5925, wire_1790, wire_5933, wire_1787, wire_5941, wire_1787, wire_5949, wire_1784, wire_5957, wire_1784, wire_5965, wire_1781, wire_5973, wire_1781, wire_5981, wire_1778, wire_5989, wire_1778, wire_5997, wire_1775, wire_6005, wire_1775, wire_6013, wire_1772, wire_6021, wire_1772, wire_6029, wire_1846, wire_1769, wire_6037, wire_1846, wire_1769, wire_5887, wire_1842, wire_5895, wire_1842, wire_5903, wire_1838, wire_5911, wire_1838, wire_5919, wire_1790, wire_5927, wire_1790, wire_5935, wire_1787, wire_5943, wire_1787, wire_5951, wire_1784, wire_5959, wire_1784, wire_5967, wire_1781, wire_5975, wire_1781, wire_5983, wire_1778, wire_5991, wire_1778, wire_5999, wire_1775, wire_6007, wire_1775, wire_6015, wire_1772, wire_6023, wire_1772, wire_6031, wire_1846, wire_1769, wire_6039, wire_1846, wire_1769};
    // CHNAXY TOTAL: 100
    assign wire_2521 = io_tile_0_5_chanxy_out[0];
    assign wire_2523 = io_tile_0_5_chanxy_out[1];
    assign wire_2525 = io_tile_0_5_chanxy_out[2];
    assign wire_2527 = io_tile_0_5_chanxy_out[3];
    assign wire_2529 = io_tile_0_5_chanxy_out[4];
    assign wire_2531 = io_tile_0_5_chanxy_out[5];
    assign wire_2533 = io_tile_0_5_chanxy_out[6];
    assign wire_2535 = io_tile_0_5_chanxy_out[7];
    assign wire_2537 = io_tile_0_5_chanxy_out[8];
    assign wire_2539 = io_tile_0_5_chanxy_out[9];
    assign wire_2541 = io_tile_0_5_chanxy_out[10];
    assign wire_2543 = io_tile_0_5_chanxy_out[11];
    assign wire_2545 = io_tile_0_5_chanxy_out[12];
    assign wire_2547 = io_tile_0_5_chanxy_out[13];
    assign wire_2549 = io_tile_0_5_chanxy_out[14];
    assign wire_2551 = io_tile_0_5_chanxy_out[15];
    assign wire_2553 = io_tile_0_5_chanxy_out[16];
    assign wire_2555 = io_tile_0_5_chanxy_out[17];
    assign wire_2557 = io_tile_0_5_chanxy_out[18];
    assign wire_2559 = io_tile_0_5_chanxy_out[19];
    assign wire_2561 = io_tile_0_5_chanxy_out[20];
    assign wire_2563 = io_tile_0_5_chanxy_out[21];
    assign wire_2565 = io_tile_0_5_chanxy_out[22];
    assign wire_2567 = io_tile_0_5_chanxy_out[23];
    assign wire_2569 = io_tile_0_5_chanxy_out[24];
    assign wire_2571 = io_tile_0_5_chanxy_out[25];
    assign wire_2573 = io_tile_0_5_chanxy_out[26];
    assign wire_2575 = io_tile_0_5_chanxy_out[27];
    assign wire_2577 = io_tile_0_5_chanxy_out[28];
    assign wire_2579 = io_tile_0_5_chanxy_out[29];
    assign wire_2581 = io_tile_0_5_chanxy_out[30];
    assign wire_2583 = io_tile_0_5_chanxy_out[31];
    assign wire_2585 = io_tile_0_5_chanxy_out[32];
    assign wire_2587 = io_tile_0_5_chanxy_out[33];
    assign wire_2589 = io_tile_0_5_chanxy_out[34];
    assign wire_2591 = io_tile_0_5_chanxy_out[35];
    assign wire_2593 = io_tile_0_5_chanxy_out[36];
    assign wire_2595 = io_tile_0_5_chanxy_out[37];
    assign wire_2597 = io_tile_0_5_chanxy_out[38];
    assign wire_2599 = io_tile_0_5_chanxy_out[39];
    assign wire_2601 = io_tile_0_5_chanxy_out[40];
    assign wire_2603 = io_tile_0_5_chanxy_out[41];
    assign wire_2605 = io_tile_0_5_chanxy_out[42];
    assign wire_2607 = io_tile_0_5_chanxy_out[43];
    assign wire_2609 = io_tile_0_5_chanxy_out[44];
    assign wire_2611 = io_tile_0_5_chanxy_out[45];
    assign wire_2613 = io_tile_0_5_chanxy_out[46];
    assign wire_2615 = io_tile_0_5_chanxy_out[47];
    assign wire_2617 = io_tile_0_5_chanxy_out[48];
    assign wire_2619 = io_tile_0_5_chanxy_out[49];
    assign wire_2621 = io_tile_0_5_chanxy_out[50];
    assign wire_2623 = io_tile_0_5_chanxy_out[51];
    assign wire_2625 = io_tile_0_5_chanxy_out[52];
    assign wire_2627 = io_tile_0_5_chanxy_out[53];
    assign wire_2629 = io_tile_0_5_chanxy_out[54];
    assign wire_2631 = io_tile_0_5_chanxy_out[55];
    assign wire_2633 = io_tile_0_5_chanxy_out[56];
    assign wire_2635 = io_tile_0_5_chanxy_out[57];
    assign wire_2637 = io_tile_0_5_chanxy_out[58];
    assign wire_2639 = io_tile_0_5_chanxy_out[59];
    assign wire_2640 = io_tile_0_5_chanxy_out[60];
    assign wire_2641 = io_tile_0_5_chanxy_out[61];
    assign wire_2642 = io_tile_0_5_chanxy_out[62];
    assign wire_2643 = io_tile_0_5_chanxy_out[63];
    assign wire_2644 = io_tile_0_5_chanxy_out[64];
    assign wire_2645 = io_tile_0_5_chanxy_out[65];
    assign wire_2646 = io_tile_0_5_chanxy_out[66];
    assign wire_2647 = io_tile_0_5_chanxy_out[67];
    assign wire_2648 = io_tile_0_5_chanxy_out[68];
    assign wire_2649 = io_tile_0_5_chanxy_out[69];
    assign wire_2650 = io_tile_0_5_chanxy_out[70];
    assign wire_2651 = io_tile_0_5_chanxy_out[71];
    assign wire_2652 = io_tile_0_5_chanxy_out[72];
    assign wire_2653 = io_tile_0_5_chanxy_out[73];
    assign wire_2654 = io_tile_0_5_chanxy_out[74];
    assign wire_2655 = io_tile_0_5_chanxy_out[75];
    assign wire_2656 = io_tile_0_5_chanxy_out[76];
    assign wire_2657 = io_tile_0_5_chanxy_out[77];
    assign wire_2658 = io_tile_0_5_chanxy_out[78];
    assign wire_2659 = io_tile_0_5_chanxy_out[79];
    assign wire_2660 = io_tile_0_5_chanxy_out[80];
    assign wire_2661 = io_tile_0_5_chanxy_out[81];
    assign wire_2662 = io_tile_0_5_chanxy_out[82];
    assign wire_2663 = io_tile_0_5_chanxy_out[83];
    assign wire_2664 = io_tile_0_5_chanxy_out[84];
    assign wire_2665 = io_tile_0_5_chanxy_out[85];
    assign wire_2666 = io_tile_0_5_chanxy_out[86];
    assign wire_2667 = io_tile_0_5_chanxy_out[87];
    assign wire_2668 = io_tile_0_5_chanxy_out[88];
    assign wire_2669 = io_tile_0_5_chanxy_out[89];
    assign wire_2670 = io_tile_0_5_chanxy_out[90];
    assign wire_2671 = io_tile_0_5_chanxy_out[91];
    assign wire_2672 = io_tile_0_5_chanxy_out[92];
    assign wire_2673 = io_tile_0_5_chanxy_out[93];
    assign wire_2674 = io_tile_0_5_chanxy_out[94];
    assign wire_2675 = io_tile_0_5_chanxy_out[95];
    assign wire_2676 = io_tile_0_5_chanxy_out[96];
    assign wire_2677 = io_tile_0_5_chanxy_out[97];
    assign wire_2678 = io_tile_0_5_chanxy_out[98];
    assign wire_2679 = io_tile_0_5_chanxy_out[99];
endmodule
