



module sbcb_sp(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [839:0] io_chanxy_in,
    input [399:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[199:0] io_chanxy_out);

  wire[199:0] T0;
  wire[199:0] T1;
  wire[198:0] T2;
  wire[198:0] T3;
  wire[197:0] T4;
  wire[197:0] T5;
  wire[196:0] T6;
  wire[196:0] T7;
  wire[195:0] T8;
  wire[195:0] T9;
  wire[194:0] T10;
  wire[194:0] T11;
  wire[193:0] T12;
  wire[193:0] T13;
  wire[192:0] T14;
  wire[192:0] T15;
  wire[191:0] T16;
  wire[191:0] T17;
  wire[190:0] T18;
  wire[190:0] T19;
  wire[189:0] T20;
  wire[189:0] T21;
  wire[188:0] T22;
  wire[188:0] T23;
  wire[187:0] T24;
  wire[187:0] T25;
  wire[186:0] T26;
  wire[186:0] T27;
  wire[185:0] T28;
  wire[185:0] T29;
  wire[184:0] T30;
  wire[184:0] T31;
  wire[183:0] T32;
  wire[183:0] T33;
  wire[182:0] T34;
  wire[182:0] T35;
  wire[181:0] T36;
  wire[181:0] T37;
  wire[180:0] T38;
  wire[180:0] T39;
  wire[179:0] T40;
  wire[179:0] T41;
  wire[178:0] T42;
  wire[178:0] T43;
  wire[177:0] T44;
  wire[177:0] T45;
  wire[176:0] T46;
  wire[176:0] T47;
  wire[175:0] T48;
  wire[175:0] T49;
  wire[174:0] T50;
  wire[174:0] T51;
  wire[173:0] T52;
  wire[173:0] T53;
  wire[172:0] T54;
  wire[172:0] T55;
  wire[171:0] T56;
  wire[171:0] T57;
  wire[170:0] T58;
  wire[170:0] T59;
  wire[169:0] T60;
  wire[169:0] T61;
  wire[168:0] T62;
  wire[168:0] T63;
  wire[167:0] T64;
  wire[167:0] T65;
  wire[166:0] T66;
  wire[166:0] T67;
  wire[165:0] T68;
  wire[165:0] T69;
  wire[164:0] T70;
  wire[164:0] T71;
  wire[163:0] T72;
  wire[163:0] T73;
  wire[162:0] T74;
  wire[162:0] T75;
  wire[161:0] T76;
  wire[161:0] T77;
  wire[160:0] T78;
  wire[160:0] T79;
  wire[159:0] T80;
  wire[159:0] T81;
  wire[158:0] T82;
  wire[158:0] T83;
  wire[157:0] T84;
  wire[157:0] T85;
  wire[156:0] T86;
  wire[156:0] T87;
  wire[155:0] T88;
  wire[155:0] T89;
  wire[154:0] T90;
  wire[154:0] T91;
  wire[153:0] T92;
  wire[153:0] T93;
  wire[152:0] T94;
  wire[152:0] T95;
  wire[151:0] T96;
  wire[151:0] T97;
  wire[150:0] T98;
  wire[150:0] T99;
  wire[149:0] T100;
  wire[149:0] T101;
  wire[148:0] T102;
  wire[148:0] T103;
  wire[147:0] T104;
  wire[147:0] T105;
  wire[146:0] T106;
  wire[146:0] T107;
  wire[145:0] T108;
  wire[145:0] T109;
  wire[144:0] T110;
  wire[144:0] T111;
  wire[143:0] T112;
  wire[143:0] T113;
  wire[142:0] T114;
  wire[142:0] T115;
  wire[141:0] T116;
  wire[141:0] T117;
  wire[140:0] T118;
  wire[140:0] T119;
  wire[139:0] T120;
  wire[139:0] T121;
  wire[138:0] T122;
  wire[138:0] T123;
  wire[137:0] T124;
  wire[137:0] T125;
  wire[136:0] T126;
  wire[136:0] T127;
  wire[135:0] T128;
  wire[135:0] T129;
  wire[134:0] T130;
  wire[134:0] T131;
  wire[133:0] T132;
  wire[133:0] T133;
  wire[132:0] T134;
  wire[132:0] T135;
  wire[131:0] T136;
  wire[131:0] T137;
  wire[130:0] T138;
  wire[130:0] T139;
  wire[129:0] T140;
  wire[129:0] T141;
  wire[128:0] T142;
  wire[128:0] T143;
  wire[127:0] T144;
  wire[127:0] T145;
  wire[126:0] T146;
  wire[126:0] T147;
  wire[125:0] T148;
  wire[125:0] T149;
  wire[124:0] T150;
  wire[124:0] T151;
  wire[123:0] T152;
  wire[123:0] T153;
  wire[122:0] T154;
  wire[122:0] T155;
  wire[121:0] T156;
  wire[121:0] T157;
  wire[120:0] T158;
  wire[120:0] T159;
  wire[119:0] T160;
  wire[119:0] T161;
  wire[118:0] T162;
  wire[118:0] T163;
  wire[117:0] T164;
  wire[117:0] T165;
  wire[116:0] T166;
  wire[116:0] T167;
  wire[115:0] T168;
  wire[115:0] T169;
  wire[114:0] T170;
  wire[114:0] T171;
  wire[113:0] T172;
  wire[113:0] T173;
  wire[112:0] T174;
  wire[112:0] T175;
  wire[111:0] T176;
  wire[111:0] T177;
  wire[110:0] T178;
  wire[110:0] T179;
  wire[109:0] T180;
  wire[109:0] T181;
  wire[108:0] T182;
  wire[108:0] T183;
  wire[107:0] T184;
  wire[107:0] T185;
  wire[106:0] T186;
  wire[106:0] T187;
  wire[105:0] T188;
  wire[105:0] T189;
  wire[104:0] T190;
  wire[104:0] T191;
  wire[103:0] T192;
  wire[103:0] T193;
  wire[102:0] T194;
  wire[102:0] T195;
  wire[101:0] T196;
  wire[101:0] T197;
  wire[100:0] T198;
  wire[100:0] T199;
  wire[99:0] T200;
  wire[99:0] T201;
  wire[98:0] T202;
  wire[98:0] T203;
  wire[97:0] T204;
  wire[97:0] T205;
  wire[96:0] T206;
  wire[96:0] T207;
  wire[95:0] T208;
  wire[95:0] T209;
  wire[94:0] T210;
  wire[94:0] T211;
  wire[93:0] T212;
  wire[93:0] T213;
  wire[92:0] T214;
  wire[92:0] T215;
  wire[91:0] T216;
  wire[91:0] T217;
  wire[90:0] T218;
  wire[90:0] T219;
  wire[89:0] T220;
  wire[89:0] T221;
  wire[88:0] T222;
  wire[88:0] T223;
  wire[87:0] T224;
  wire[87:0] T225;
  wire[86:0] T226;
  wire[86:0] T227;
  wire[85:0] T228;
  wire[85:0] T229;
  wire[84:0] T230;
  wire[84:0] T231;
  wire[83:0] T232;
  wire[83:0] T233;
  wire[82:0] T234;
  wire[82:0] T235;
  wire[81:0] T236;
  wire[81:0] T237;
  wire[80:0] T238;
  wire[80:0] T239;
  wire[79:0] T240;
  wire[79:0] T241;
  wire[78:0] T242;
  wire[78:0] T243;
  wire[77:0] T244;
  wire[77:0] T245;
  wire[76:0] T246;
  wire[76:0] T247;
  wire[75:0] T248;
  wire[75:0] T249;
  wire[74:0] T250;
  wire[74:0] T251;
  wire[73:0] T252;
  wire[73:0] T253;
  wire[72:0] T254;
  wire[72:0] T255;
  wire[71:0] T256;
  wire[71:0] T257;
  wire[70:0] T258;
  wire[70:0] T259;
  wire[69:0] T260;
  wire[69:0] T261;
  wire[68:0] T262;
  wire[68:0] T263;
  wire[67:0] T264;
  wire[67:0] T265;
  wire[66:0] T266;
  wire[66:0] T267;
  wire[65:0] T268;
  wire[65:0] T269;
  wire[64:0] T270;
  wire[64:0] T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[62:0] T274;
  wire[62:0] T275;
  wire[61:0] T276;
  wire[61:0] T277;
  wire[60:0] T278;
  wire[60:0] T279;
  wire[59:0] T280;
  wire[59:0] T281;
  wire[58:0] T282;
  wire[58:0] T283;
  wire[57:0] T284;
  wire[57:0] T285;
  wire[56:0] T286;
  wire[56:0] T287;
  wire[55:0] T288;
  wire[55:0] T289;
  wire[54:0] T290;
  wire[54:0] T291;
  wire[53:0] T292;
  wire[53:0] T293;
  wire[52:0] T294;
  wire[52:0] T295;
  wire[51:0] T296;
  wire[51:0] T297;
  wire[50:0] T298;
  wire[50:0] T299;
  wire[49:0] T300;
  wire[49:0] T301;
  wire[48:0] T302;
  wire[48:0] T303;
  wire[47:0] T304;
  wire[47:0] T305;
  wire[46:0] T306;
  wire[46:0] T307;
  wire[45:0] T308;
  wire[45:0] T309;
  wire[44:0] T310;
  wire[44:0] T311;
  wire[43:0] T312;
  wire[43:0] T313;
  wire[42:0] T314;
  wire[42:0] T315;
  wire[41:0] T316;
  wire[41:0] T317;
  wire[40:0] T318;
  wire[40:0] T319;
  wire[39:0] T320;
  wire[39:0] T321;
  wire[38:0] T322;
  wire[38:0] T323;
  wire[37:0] T324;
  wire[37:0] T325;
  wire[36:0] T326;
  wire[36:0] T327;
  wire[35:0] T328;
  wire[35:0] T329;
  wire[34:0] T330;
  wire[34:0] T331;
  wire[33:0] T332;
  wire[33:0] T333;
  wire[32:0] T334;
  wire[32:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[30:0] T338;
  wire[30:0] T339;
  wire[29:0] T340;
  wire[29:0] T341;
  wire[28:0] T342;
  wire[28:0] T343;
  wire[27:0] T344;
  wire[27:0] T345;
  wire[26:0] T346;
  wire[26:0] T347;
  wire[25:0] T348;
  wire[25:0] T349;
  wire[24:0] T350;
  wire[24:0] T351;
  wire[23:0] T352;
  wire[23:0] T353;
  wire[22:0] T354;
  wire[22:0] T355;
  wire[21:0] T356;
  wire[21:0] T357;
  wire[20:0] T358;
  wire[20:0] T359;
  wire[19:0] T360;
  wire[19:0] T361;
  wire[18:0] T362;
  wire[18:0] T363;
  wire[17:0] T364;
  wire[17:0] T365;
  wire[16:0] T366;
  wire[16:0] T367;
  wire[15:0] T368;
  wire[15:0] T369;
  wire[14:0] T370;
  wire[14:0] T371;
  wire[13:0] T372;
  wire[13:0] T373;
  wire[12:0] T374;
  wire[12:0] T375;
  wire[11:0] T376;
  wire[11:0] T377;
  wire[10:0] T378;
  wire[10:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[6:0] T386;
  wire[6:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[3:0] T393;
  wire[2:0] T394;
  wire[2:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire[1:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[1:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire[2:0] T412;
  wire[2:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[1:0] T417;
  wire[1:0] T418;
  wire[1:0] T419;
  wire[2:0] T420;
  wire[2:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[10:0] T428;
  wire[10:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[2:0] T436;
  wire[2:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[1:0] T449;
  wire[1:0] T450;
  wire[1:0] T451;
  wire[2:0] T452;
  wire[2:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[1:0] T457;
  wire[1:0] T458;
  wire[1:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[10:0] T468;
  wire[10:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire[1:0] T475;
  wire[2:0] T476;
  wire[2:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[1:0] T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[2:0] T484;
  wire[2:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[1:0] T489;
  wire[1:0] T490;
  wire[1:0] T491;
  wire[2:0] T492;
  wire[2:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[2:0] T500;
  wire[2:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[10:0] T508;
  wire[10:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[1:0] T513;
  wire[1:0] T514;
  wire[1:0] T515;
  wire[2:0] T516;
  wire[2:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire[1:0] T523;
  wire[2:0] T524;
  wire[2:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[1:0] T529;
  wire[1:0] T530;
  wire[1:0] T531;
  wire[2:0] T532;
  wire[2:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[1:0] T537;
  wire[1:0] T538;
  wire[1:0] T539;
  wire[2:0] T540;
  wire[2:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[10:0] T548;
  wire[10:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[1:0] T553;
  wire[1:0] T554;
  wire[1:0] T555;
  wire[2:0] T556;
  wire[2:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[1:0] T561;
  wire[1:0] T562;
  wire[1:0] T563;
  wire[2:0] T564;
  wire[2:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[1:0] T569;
  wire[1:0] T570;
  wire[1:0] T571;
  wire[2:0] T572;
  wire[2:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[1:0] T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[2:0] T580;
  wire[2:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[10:0] T588;
  wire[10:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[1:0] T593;
  wire[1:0] T594;
  wire[1:0] T595;
  wire[2:0] T596;
  wire[2:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[3:0] T625;
  wire[3:0] T626;
  wire[3:0] T627;
  wire[10:0] T628;
  wire[10:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[3:0] T665;
  wire[3:0] T666;
  wire[3:0] T667;
  wire[10:0] T668;
  wire[10:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire[1:0] T683;
  wire[2:0] T684;
  wire[2:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[1:0] T689;
  wire[1:0] T690;
  wire[1:0] T691;
  wire[2:0] T692;
  wire[2:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[1:0] T697;
  wire[1:0] T698;
  wire[1:0] T699;
  wire[2:0] T700;
  wire[2:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[3:0] T705;
  wire[3:0] T706;
  wire[3:0] T707;
  wire[10:0] T708;
  wire[10:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[1:0] T713;
  wire[1:0] T714;
  wire[1:0] T715;
  wire[2:0] T716;
  wire[2:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[2:0] T724;
  wire[2:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[1:0] T729;
  wire[1:0] T730;
  wire[1:0] T731;
  wire[2:0] T732;
  wire[2:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[1:0] T737;
  wire[1:0] T738;
  wire[1:0] T739;
  wire[2:0] T740;
  wire[2:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[3:0] T745;
  wire[3:0] T746;
  wire[3:0] T747;
  wire[10:0] T748;
  wire[10:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[1:0] T753;
  wire[1:0] T754;
  wire[1:0] T755;
  wire[2:0] T756;
  wire[2:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[1:0] T777;
  wire[1:0] T778;
  wire[1:0] T779;
  wire[2:0] T780;
  wire[2:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[3:0] T785;
  wire[3:0] T786;
  wire[3:0] T787;
  wire[10:0] T788;
  wire[10:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[1:0] T793;
  wire[1:0] T794;
  wire[1:0] T795;
  wire[2:0] T796;
  wire[2:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[10:0] T828;
  wire[10:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[3:0] T865;
  wire[3:0] T866;
  wire[3:0] T867;
  wire[10:0] T868;
  wire[10:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[3:0] T905;
  wire[3:0] T906;
  wire[3:0] T907;
  wire[10:0] T908;
  wire[10:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire[1:0] T940;
  wire[1:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[3:0] T945;
  wire[3:0] T946;
  wire[3:0] T947;
  wire[10:0] T948;
  wire[10:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[3:0] T985;
  wire[3:0] T986;
  wire[3:0] T987;
  wire[10:0] T988;
  wire[10:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire[3:0] T1025;
  wire[3:0] T1026;
  wire[3:0] T1027;
  wire[10:0] T1028;
  wire[10:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire[3:0] T1065;
  wire[3:0] T1066;
  wire[3:0] T1067;
  wire[10:0] T1068;
  wire[10:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire[1:0] T1092;
  wire[1:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[10:0] T1108;
  wire[10:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire[1:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire[1:0] T1140;
  wire[1:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[10:0] T1148;
  wire[10:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire[1:0] T1156;
  wire[1:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire[1:0] T1172;
  wire[1:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[10:0] T1188;
  wire[10:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[1:0] T1201;
  wire[1:0] T1202;
  wire[1:0] T1203;
  wire[2:0] T1204;
  wire[2:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[1:0] T1209;
  wire[1:0] T1210;
  wire[1:0] T1211;
  wire[2:0] T1212;
  wire[2:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[2:0] T1220;
  wire[2:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[10:0] T1228;
  wire[10:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[1:0] T1233;
  wire[1:0] T1234;
  wire[1:0] T1235;
  wire[2:0] T1236;
  wire[2:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[1:0] T1241;
  wire[1:0] T1242;
  wire[1:0] T1243;
  wire[2:0] T1244;
  wire[2:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[1:0] T1249;
  wire[1:0] T1250;
  wire[1:0] T1251;
  wire[2:0] T1252;
  wire[2:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[1:0] T1257;
  wire[1:0] T1258;
  wire[1:0] T1259;
  wire[2:0] T1260;
  wire[2:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[10:0] T1268;
  wire[10:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[1:0] T1273;
  wire[1:0] T1274;
  wire[1:0] T1275;
  wire[2:0] T1276;
  wire[2:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire[1:0] T1281;
  wire[1:0] T1282;
  wire[1:0] T1283;
  wire[2:0] T1284;
  wire[2:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[1:0] T1289;
  wire[1:0] T1290;
  wire[1:0] T1291;
  wire[2:0] T1292;
  wire[2:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[1:0] T1297;
  wire[1:0] T1298;
  wire[1:0] T1299;
  wire[2:0] T1300;
  wire[2:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[10:0] T1308;
  wire[10:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[1:0] T1313;
  wire[1:0] T1314;
  wire[1:0] T1315;
  wire[2:0] T1316;
  wire[2:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[1:0] T1321;
  wire[1:0] T1322;
  wire[1:0] T1323;
  wire[2:0] T1324;
  wire[2:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[1:0] T1329;
  wire[1:0] T1330;
  wire[1:0] T1331;
  wire[2:0] T1332;
  wire[2:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[1:0] T1337;
  wire[1:0] T1338;
  wire[1:0] T1339;
  wire[2:0] T1340;
  wire[2:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[10:0] T1348;
  wire[10:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[1:0] T1353;
  wire[1:0] T1354;
  wire[1:0] T1355;
  wire[2:0] T1356;
  wire[2:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[2:0] T1364;
  wire[2:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[1:0] T1369;
  wire[1:0] T1370;
  wire[1:0] T1371;
  wire[2:0] T1372;
  wire[2:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[1:0] T1377;
  wire[1:0] T1378;
  wire[1:0] T1379;
  wire[2:0] T1380;
  wire[2:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[10:0] T1388;
  wire[10:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[1:0] T1393;
  wire[1:0] T1394;
  wire[1:0] T1395;
  wire[2:0] T1396;
  wire[2:0] T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire[1:0] T1401;
  wire[1:0] T1402;
  wire[1:0] T1403;
  wire[2:0] T1404;
  wire[2:0] T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire[1:0] T1409;
  wire[1:0] T1410;
  wire[1:0] T1411;
  wire[2:0] T1412;
  wire[2:0] T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire[1:0] T1417;
  wire[1:0] T1418;
  wire[1:0] T1419;
  wire[2:0] T1420;
  wire[2:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire[3:0] T1425;
  wire[3:0] T1426;
  wire[3:0] T1427;
  wire[10:0] T1428;
  wire[10:0] T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire[1:0] T1433;
  wire[1:0] T1434;
  wire[1:0] T1435;
  wire[2:0] T1436;
  wire[2:0] T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire[1:0] T1441;
  wire[1:0] T1442;
  wire[1:0] T1443;
  wire[2:0] T1444;
  wire[2:0] T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire[1:0] T1449;
  wire[1:0] T1450;
  wire[1:0] T1451;
  wire[2:0] T1452;
  wire[2:0] T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire[1:0] T1457;
  wire[1:0] T1458;
  wire[1:0] T1459;
  wire[2:0] T1460;
  wire[2:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[10:0] T1468;
  wire[10:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[1:0] T1473;
  wire[1:0] T1474;
  wire[1:0] T1475;
  wire[2:0] T1476;
  wire[2:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[1:0] T1481;
  wire[1:0] T1482;
  wire[1:0] T1483;
  wire[2:0] T1484;
  wire[2:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[1:0] T1489;
  wire[1:0] T1490;
  wire[1:0] T1491;
  wire[2:0] T1492;
  wire[2:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[1:0] T1497;
  wire[1:0] T1498;
  wire[1:0] T1499;
  wire[2:0] T1500;
  wire[2:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[10:0] T1508;
  wire[10:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[1:0] T1513;
  wire[1:0] T1514;
  wire[1:0] T1515;
  wire[2:0] T1516;
  wire[2:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[1:0] T1521;
  wire[1:0] T1522;
  wire[1:0] T1523;
  wire[2:0] T1524;
  wire[2:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[1:0] T1529;
  wire[1:0] T1530;
  wire[1:0] T1531;
  wire[2:0] T1532;
  wire[2:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[1:0] T1537;
  wire[1:0] T1538;
  wire[1:0] T1539;
  wire[2:0] T1540;
  wire[2:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[10:0] T1548;
  wire[10:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[1:0] T1553;
  wire[1:0] T1554;
  wire[1:0] T1555;
  wire[2:0] T1556;
  wire[2:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[1:0] T1561;
  wire[1:0] T1562;
  wire[1:0] T1563;
  wire[2:0] T1564;
  wire[2:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[1:0] T1569;
  wire[1:0] T1570;
  wire[1:0] T1571;
  wire[2:0] T1572;
  wire[2:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[1:0] T1577;
  wire[1:0] T1578;
  wire[1:0] T1579;
  wire[2:0] T1580;
  wire[2:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[10:0] T1588;
  wire[10:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[1:0] T1593;
  wire[1:0] T1594;
  wire[1:0] T1595;
  wire[2:0] T1596;
  wire[2:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire[1:0] T1604;
  wire[1:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[1:0] T1612;
  wire[1:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire[1:0] T1620;
  wire[1:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[10:0] T1628;
  wire[10:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire[1:0] T1636;
  wire[1:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire[1:0] T1644;
  wire[1:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire[1:0] T1652;
  wire[1:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire[1:0] T1660;
  wire[1:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[10:0] T1668;
  wire[10:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire[1:0] T1676;
  wire[1:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire[1:0] T1684;
  wire[1:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire T1689;
  wire T1690;
  wire T1691;
  wire[1:0] T1692;
  wire[1:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[1:0] T1700;
  wire[1:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[10:0] T1708;
  wire[10:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire[1:0] T1716;
  wire[1:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[1:0] T1724;
  wire[1:0] T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire[1:0] T1732;
  wire[1:0] T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire T1738;
  wire T1739;
  wire[1:0] T1740;
  wire[1:0] T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire[3:0] T1745;
  wire[3:0] T1746;
  wire[3:0] T1747;
  wire[10:0] T1748;
  wire[10:0] T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire T1753;
  wire T1754;
  wire T1755;
  wire[1:0] T1756;
  wire[1:0] T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire T1762;
  wire T1763;
  wire[1:0] T1764;
  wire[1:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire T1770;
  wire T1771;
  wire[1:0] T1772;
  wire[1:0] T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire T1779;
  wire[1:0] T1780;
  wire[1:0] T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire[3:0] T1785;
  wire[3:0] T1786;
  wire[3:0] T1787;
  wire[10:0] T1788;
  wire[10:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire[1:0] T1796;
  wire[1:0] T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire[1:0] T1804;
  wire[1:0] T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire[1:0] T1812;
  wire[1:0] T1813;
  wire T1814;
  wire T1815;
  wire T1816;
  wire T1817;
  wire T1818;
  wire T1819;
  wire[1:0] T1820;
  wire[1:0] T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[3:0] T1825;
  wire[3:0] T1826;
  wire[3:0] T1827;
  wire[10:0] T1828;
  wire[10:0] T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire T1834;
  wire T1835;
  wire[1:0] T1836;
  wire[1:0] T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire T1842;
  wire T1843;
  wire[1:0] T1844;
  wire[1:0] T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire T1851;
  wire[1:0] T1852;
  wire[1:0] T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire T1859;
  wire[1:0] T1860;
  wire[1:0] T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire[3:0] T1865;
  wire[3:0] T1866;
  wire[3:0] T1867;
  wire[10:0] T1868;
  wire[10:0] T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire[1:0] T1876;
  wire[1:0] T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire[1:0] T1892;
  wire[1:0] T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[1:0] T1900;
  wire[1:0] T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire[3:0] T1905;
  wire[3:0] T1906;
  wire[3:0] T1907;
  wire[10:0] T1908;
  wire[10:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire[1:0] T1916;
  wire[1:0] T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire T1921;
  wire T1922;
  wire T1923;
  wire[1:0] T1924;
  wire[1:0] T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire[1:0] T1932;
  wire[1:0] T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire T1937;
  wire T1938;
  wire T1939;
  wire[1:0] T1940;
  wire[1:0] T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire[3:0] T1945;
  wire[3:0] T1946;
  wire[3:0] T1947;
  wire[10:0] T1948;
  wire[10:0] T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire T1955;
  wire[1:0] T1956;
  wire[1:0] T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire[1:0] T1964;
  wire[1:0] T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire[1:0] T1972;
  wire[1:0] T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire[1:0] T1980;
  wire[1:0] T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire[3:0] T1985;
  wire[3:0] T1986;
  wire[3:0] T1987;
  wire[10:0] T1988;
  wire[10:0] T1989;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire[1:0] T1996;
  wire[1:0] T1997;
  wire[32:0] T1998;
  wire[32:0] T1999;
  wire[31:0] T2000;
  wire[31:0] T2001;
  wire[30:0] T2002;
  wire[30:0] T2003;
  wire[29:0] T2004;
  wire[29:0] T2005;
  wire[28:0] T2006;
  wire[28:0] T2007;
  wire[27:0] T2008;
  wire[27:0] T2009;
  wire[26:0] T2010;
  wire[26:0] T2011;
  wire[25:0] T2012;
  wire[25:0] T2013;
  wire[24:0] T2014;
  wire[24:0] T2015;
  wire[23:0] T2016;
  wire[23:0] T2017;
  wire[22:0] T2018;
  wire[22:0] T2019;
  wire[21:0] T2020;
  wire[21:0] T2021;
  wire[20:0] T2022;
  wire[20:0] T2023;
  wire[19:0] T2024;
  wire[19:0] T2025;
  wire[18:0] T2026;
  wire[18:0] T2027;
  wire[17:0] T2028;
  wire[17:0] T2029;
  wire[16:0] T2030;
  wire[16:0] T2031;
  wire[15:0] T2032;
  wire[15:0] T2033;
  wire[14:0] T2034;
  wire[14:0] T2035;
  wire[13:0] T2036;
  wire[13:0] T2037;
  wire[12:0] T2038;
  wire[12:0] T2039;
  wire[11:0] T2040;
  wire[11:0] T2041;
  wire[10:0] T2042;
  wire[10:0] T2043;
  wire[9:0] T2044;
  wire[9:0] T2045;
  wire[8:0] T2046;
  wire[8:0] T2047;
  wire[7:0] T2048;
  wire[7:0] T2049;
  wire[6:0] T2050;
  wire[6:0] T2051;
  wire[5:0] T2052;
  wire[5:0] T2053;
  wire[4:0] T2054;
  wire[4:0] T2055;
  wire[3:0] T2056;
  wire[3:0] T2057;
  wire[2:0] T2058;
  wire[2:0] T2059;
  wire[1:0] T2060;
  wire[1:0] T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire[3:0] T2065;
  wire[3:0] T2066;
  wire[3:0] T2067;
  wire[15:0] T2068;
  wire[15:0] T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire[3:0] T2073;
  wire[3:0] T2074;
  wire[3:0] T2075;
  wire[15:0] T2076;
  wire[15:0] T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[3:0] T2081;
  wire[3:0] T2082;
  wire[3:0] T2083;
  wire[15:0] T2084;
  wire[15:0] T2085;
  wire T2086;
  wire T2087;
  wire T2088;
  wire[3:0] T2089;
  wire[3:0] T2090;
  wire[3:0] T2091;
  wire[15:0] T2092;
  wire[15:0] T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire[3:0] T2097;
  wire[3:0] T2098;
  wire[3:0] T2099;
  wire[15:0] T2100;
  wire[15:0] T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire[3:0] T2105;
  wire[3:0] T2106;
  wire[3:0] T2107;
  wire[15:0] T2108;
  wire[15:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire[3:0] T2113;
  wire[3:0] T2114;
  wire[3:0] T2115;
  wire[15:0] T2116;
  wire[15:0] T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[3:0] T2121;
  wire[3:0] T2122;
  wire[3:0] T2123;
  wire[15:0] T2124;
  wire[15:0] T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire[3:0] T2129;
  wire[3:0] T2130;
  wire[3:0] T2131;
  wire[15:0] T2132;
  wire[15:0] T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire[3:0] T2137;
  wire[3:0] T2138;
  wire[3:0] T2139;
  wire[15:0] T2140;
  wire[15:0] T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire[3:0] T2145;
  wire[3:0] T2146;
  wire[3:0] T2147;
  wire[15:0] T2148;
  wire[15:0] T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire[3:0] T2153;
  wire[3:0] T2154;
  wire[3:0] T2155;
  wire[15:0] T2156;
  wire[15:0] T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire[3:0] T2161;
  wire[3:0] T2162;
  wire[3:0] T2163;
  wire[15:0] T2164;
  wire[15:0] T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire[3:0] T2169;
  wire[3:0] T2170;
  wire[3:0] T2171;
  wire[15:0] T2172;
  wire[15:0] T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  wire[3:0] T2177;
  wire[3:0] T2178;
  wire[3:0] T2179;
  wire[15:0] T2180;
  wire[15:0] T2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire[3:0] T2185;
  wire[3:0] T2186;
  wire[3:0] T2187;
  wire[15:0] T2188;
  wire[15:0] T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[3:0] T2193;
  wire[3:0] T2194;
  wire[3:0] T2195;
  wire[15:0] T2196;
  wire[15:0] T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire[3:0] T2201;
  wire[3:0] T2202;
  wire[3:0] T2203;
  wire[15:0] T2204;
  wire[15:0] T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire[3:0] T2209;
  wire[3:0] T2210;
  wire[3:0] T2211;
  wire[15:0] T2212;
  wire[15:0] T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire[3:0] T2217;
  wire[3:0] T2218;
  wire[3:0] T2219;
  wire[15:0] T2220;
  wire[15:0] T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire[3:0] T2225;
  wire[3:0] T2226;
  wire[3:0] T2227;
  wire[15:0] T2228;
  wire[15:0] T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire[3:0] T2233;
  wire[3:0] T2234;
  wire[3:0] T2235;
  wire[15:0] T2236;
  wire[15:0] T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire[3:0] T2241;
  wire[3:0] T2242;
  wire[3:0] T2243;
  wire[15:0] T2244;
  wire[15:0] T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  wire[3:0] T2249;
  wire[3:0] T2250;
  wire[3:0] T2251;
  wire[15:0] T2252;
  wire[15:0] T2253;
  wire T2254;
  wire T2255;
  wire T2256;
  wire[3:0] T2257;
  wire[3:0] T2258;
  wire[3:0] T2259;
  wire[15:0] T2260;
  wire[15:0] T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[3:0] T2265;
  wire[3:0] T2266;
  wire[3:0] T2267;
  wire[15:0] T2268;
  wire[15:0] T2269;
  wire T2270;
  wire T2271;
  wire T2272;
  wire[3:0] T2273;
  wire[3:0] T2274;
  wire[3:0] T2275;
  wire[15:0] T2276;
  wire[15:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire[3:0] T2281;
  wire[3:0] T2282;
  wire[3:0] T2283;
  wire[15:0] T2284;
  wire[15:0] T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire[3:0] T2289;
  wire[3:0] T2290;
  wire[3:0] T2291;
  wire[15:0] T2292;
  wire[15:0] T2293;
  wire T2294;
  wire T2295;
  wire T2296;
  wire[3:0] T2297;
  wire[3:0] T2298;
  wire[3:0] T2299;
  wire[15:0] T2300;
  wire[15:0] T2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire[3:0] T2305;
  wire[3:0] T2306;
  wire[3:0] T2307;
  wire[15:0] T2308;
  wire[15:0] T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire[3:0] T2313;
  wire[3:0] T2314;
  wire[3:0] T2315;
  wire[15:0] T2316;
  wire[15:0] T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  wire[3:0] T2321;
  wire[3:0] T2322;
  wire[3:0] T2323;
  wire[15:0] T2324;
  wire[15:0] T2325;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1990, T2};
  assign T2 = T3;
  assign T3 = {T1982, T4};
  assign T4 = T5;
  assign T5 = {T1974, T6};
  assign T6 = T7;
  assign T7 = {T1966, T8};
  assign T8 = T9;
  assign T9 = {T1958, T10};
  assign T10 = T11;
  assign T11 = {T1950, T12};
  assign T12 = T13;
  assign T13 = {T1942, T14};
  assign T14 = T15;
  assign T15 = {T1934, T16};
  assign T16 = T17;
  assign T17 = {T1926, T18};
  assign T18 = T19;
  assign T19 = {T1918, T20};
  assign T20 = T21;
  assign T21 = {T1910, T22};
  assign T22 = T23;
  assign T23 = {T1902, T24};
  assign T24 = T25;
  assign T25 = {T1894, T26};
  assign T26 = T27;
  assign T27 = {T1886, T28};
  assign T28 = T29;
  assign T29 = {T1878, T30};
  assign T30 = T31;
  assign T31 = {T1870, T32};
  assign T32 = T33;
  assign T33 = {T1862, T34};
  assign T34 = T35;
  assign T35 = {T1854, T36};
  assign T36 = T37;
  assign T37 = {T1846, T38};
  assign T38 = T39;
  assign T39 = {T1838, T40};
  assign T40 = T41;
  assign T41 = {T1830, T42};
  assign T42 = T43;
  assign T43 = {T1822, T44};
  assign T44 = T45;
  assign T45 = {T1814, T46};
  assign T46 = T47;
  assign T47 = {T1806, T48};
  assign T48 = T49;
  assign T49 = {T1798, T50};
  assign T50 = T51;
  assign T51 = {T1790, T52};
  assign T52 = T53;
  assign T53 = {T1782, T54};
  assign T54 = T55;
  assign T55 = {T1774, T56};
  assign T56 = T57;
  assign T57 = {T1766, T58};
  assign T58 = T59;
  assign T59 = {T1758, T60};
  assign T60 = T61;
  assign T61 = {T1750, T62};
  assign T62 = T63;
  assign T63 = {T1742, T64};
  assign T64 = T65;
  assign T65 = {T1734, T66};
  assign T66 = T67;
  assign T67 = {T1726, T68};
  assign T68 = T69;
  assign T69 = {T1718, T70};
  assign T70 = T71;
  assign T71 = {T1710, T72};
  assign T72 = T73;
  assign T73 = {T1702, T74};
  assign T74 = T75;
  assign T75 = {T1694, T76};
  assign T76 = T77;
  assign T77 = {T1686, T78};
  assign T78 = T79;
  assign T79 = {T1678, T80};
  assign T80 = T81;
  assign T81 = {T1670, T82};
  assign T82 = T83;
  assign T83 = {T1662, T84};
  assign T84 = T85;
  assign T85 = {T1654, T86};
  assign T86 = T87;
  assign T87 = {T1646, T88};
  assign T88 = T89;
  assign T89 = {T1638, T90};
  assign T90 = T91;
  assign T91 = {T1630, T92};
  assign T92 = T93;
  assign T93 = {T1622, T94};
  assign T94 = T95;
  assign T95 = {T1614, T96};
  assign T96 = T97;
  assign T97 = {T1606, T98};
  assign T98 = T99;
  assign T99 = {T1598, T100};
  assign T100 = T101;
  assign T101 = {T1590, T102};
  assign T102 = T103;
  assign T103 = {T1582, T104};
  assign T104 = T105;
  assign T105 = {T1574, T106};
  assign T106 = T107;
  assign T107 = {T1566, T108};
  assign T108 = T109;
  assign T109 = {T1558, T110};
  assign T110 = T111;
  assign T111 = {T1550, T112};
  assign T112 = T113;
  assign T113 = {T1542, T114};
  assign T114 = T115;
  assign T115 = {T1534, T116};
  assign T116 = T117;
  assign T117 = {T1526, T118};
  assign T118 = T119;
  assign T119 = {T1518, T120};
  assign T120 = T121;
  assign T121 = {T1510, T122};
  assign T122 = T123;
  assign T123 = {T1502, T124};
  assign T124 = T125;
  assign T125 = {T1494, T126};
  assign T126 = T127;
  assign T127 = {T1486, T128};
  assign T128 = T129;
  assign T129 = {T1478, T130};
  assign T130 = T131;
  assign T131 = {T1470, T132};
  assign T132 = T133;
  assign T133 = {T1462, T134};
  assign T134 = T135;
  assign T135 = {T1454, T136};
  assign T136 = T137;
  assign T137 = {T1446, T138};
  assign T138 = T139;
  assign T139 = {T1438, T140};
  assign T140 = T141;
  assign T141 = {T1430, T142};
  assign T142 = T143;
  assign T143 = {T1422, T144};
  assign T144 = T145;
  assign T145 = {T1414, T146};
  assign T146 = T147;
  assign T147 = {T1406, T148};
  assign T148 = T149;
  assign T149 = {T1398, T150};
  assign T150 = T151;
  assign T151 = {T1390, T152};
  assign T152 = T153;
  assign T153 = {T1382, T154};
  assign T154 = T155;
  assign T155 = {T1374, T156};
  assign T156 = T157;
  assign T157 = {T1366, T158};
  assign T158 = T159;
  assign T159 = {T1358, T160};
  assign T160 = T161;
  assign T161 = {T1350, T162};
  assign T162 = T163;
  assign T163 = {T1342, T164};
  assign T164 = T165;
  assign T165 = {T1334, T166};
  assign T166 = T167;
  assign T167 = {T1326, T168};
  assign T168 = T169;
  assign T169 = {T1318, T170};
  assign T170 = T171;
  assign T171 = {T1310, T172};
  assign T172 = T173;
  assign T173 = {T1302, T174};
  assign T174 = T175;
  assign T175 = {T1294, T176};
  assign T176 = T177;
  assign T177 = {T1286, T178};
  assign T178 = T179;
  assign T179 = {T1278, T180};
  assign T180 = T181;
  assign T181 = {T1270, T182};
  assign T182 = T183;
  assign T183 = {T1262, T184};
  assign T184 = T185;
  assign T185 = {T1254, T186};
  assign T186 = T187;
  assign T187 = {T1246, T188};
  assign T188 = T189;
  assign T189 = {T1238, T190};
  assign T190 = T191;
  assign T191 = {T1230, T192};
  assign T192 = T193;
  assign T193 = {T1222, T194};
  assign T194 = T195;
  assign T195 = {T1214, T196};
  assign T196 = T197;
  assign T197 = {T1206, T198};
  assign T198 = T199;
  assign T199 = {T1198, T200};
  assign T200 = T201;
  assign T201 = {T1190, T202};
  assign T202 = T203;
  assign T203 = {T1182, T204};
  assign T204 = T205;
  assign T205 = {T1174, T206};
  assign T206 = T207;
  assign T207 = {T1166, T208};
  assign T208 = T209;
  assign T209 = {T1158, T210};
  assign T210 = T211;
  assign T211 = {T1150, T212};
  assign T212 = T213;
  assign T213 = {T1142, T214};
  assign T214 = T215;
  assign T215 = {T1134, T216};
  assign T216 = T217;
  assign T217 = {T1126, T218};
  assign T218 = T219;
  assign T219 = {T1118, T220};
  assign T220 = T221;
  assign T221 = {T1110, T222};
  assign T222 = T223;
  assign T223 = {T1102, T224};
  assign T224 = T225;
  assign T225 = {T1094, T226};
  assign T226 = T227;
  assign T227 = {T1086, T228};
  assign T228 = T229;
  assign T229 = {T1078, T230};
  assign T230 = T231;
  assign T231 = {T1070, T232};
  assign T232 = T233;
  assign T233 = {T1062, T234};
  assign T234 = T235;
  assign T235 = {T1054, T236};
  assign T236 = T237;
  assign T237 = {T1046, T238};
  assign T238 = T239;
  assign T239 = {T1038, T240};
  assign T240 = T241;
  assign T241 = {T1030, T242};
  assign T242 = T243;
  assign T243 = {T1022, T244};
  assign T244 = T245;
  assign T245 = {T1014, T246};
  assign T246 = T247;
  assign T247 = {T1006, T248};
  assign T248 = T249;
  assign T249 = {T998, T250};
  assign T250 = T251;
  assign T251 = {T990, T252};
  assign T252 = T253;
  assign T253 = {T982, T254};
  assign T254 = T255;
  assign T255 = {T974, T256};
  assign T256 = T257;
  assign T257 = {T966, T258};
  assign T258 = T259;
  assign T259 = {T958, T260};
  assign T260 = T261;
  assign T261 = {T950, T262};
  assign T262 = T263;
  assign T263 = {T942, T264};
  assign T264 = T265;
  assign T265 = {T934, T266};
  assign T266 = T267;
  assign T267 = {T926, T268};
  assign T268 = T269;
  assign T269 = {T918, T270};
  assign T270 = T271;
  assign T271 = {T910, T272};
  assign T272 = T273;
  assign T273 = {T902, T274};
  assign T274 = T275;
  assign T275 = {T894, T276};
  assign T276 = T277;
  assign T277 = {T886, T278};
  assign T278 = T279;
  assign T279 = {T878, T280};
  assign T280 = T281;
  assign T281 = {T870, T282};
  assign T282 = T283;
  assign T283 = {T862, T284};
  assign T284 = T285;
  assign T285 = {T854, T286};
  assign T286 = T287;
  assign T287 = {T846, T288};
  assign T288 = T289;
  assign T289 = {T838, T290};
  assign T290 = T291;
  assign T291 = {T830, T292};
  assign T292 = T293;
  assign T293 = {T822, T294};
  assign T294 = T295;
  assign T295 = {T814, T296};
  assign T296 = T297;
  assign T297 = {T806, T298};
  assign T298 = T299;
  assign T299 = {T798, T300};
  assign T300 = T301;
  assign T301 = {T790, T302};
  assign T302 = T303;
  assign T303 = {T782, T304};
  assign T304 = T305;
  assign T305 = {T774, T306};
  assign T306 = T307;
  assign T307 = {T766, T308};
  assign T308 = T309;
  assign T309 = {T758, T310};
  assign T310 = T311;
  assign T311 = {T750, T312};
  assign T312 = T313;
  assign T313 = {T742, T314};
  assign T314 = T315;
  assign T315 = {T734, T316};
  assign T316 = T317;
  assign T317 = {T726, T318};
  assign T318 = T319;
  assign T319 = {T718, T320};
  assign T320 = T321;
  assign T321 = {T710, T322};
  assign T322 = T323;
  assign T323 = {T702, T324};
  assign T324 = T325;
  assign T325 = {T694, T326};
  assign T326 = T327;
  assign T327 = {T686, T328};
  assign T328 = T329;
  assign T329 = {T678, T330};
  assign T330 = T331;
  assign T331 = {T670, T332};
  assign T332 = T333;
  assign T333 = {T662, T334};
  assign T334 = T335;
  assign T335 = {T654, T336};
  assign T336 = T337;
  assign T337 = {T646, T338};
  assign T338 = T339;
  assign T339 = {T638, T340};
  assign T340 = T341;
  assign T341 = {T630, T342};
  assign T342 = T343;
  assign T343 = {T622, T344};
  assign T344 = T345;
  assign T345 = {T614, T346};
  assign T346 = T347;
  assign T347 = {T606, T348};
  assign T348 = T349;
  assign T349 = {T598, T350};
  assign T350 = T351;
  assign T351 = {T590, T352};
  assign T352 = T353;
  assign T353 = {T582, T354};
  assign T354 = T355;
  assign T355 = {T574, T356};
  assign T356 = T357;
  assign T357 = {T566, T358};
  assign T358 = T359;
  assign T359 = {T558, T360};
  assign T360 = T361;
  assign T361 = {T550, T362};
  assign T362 = T363;
  assign T363 = {T542, T364};
  assign T364 = T365;
  assign T365 = {T534, T366};
  assign T366 = T367;
  assign T367 = {T526, T368};
  assign T368 = T369;
  assign T369 = {T518, T370};
  assign T370 = T371;
  assign T371 = {T510, T372};
  assign T372 = T373;
  assign T373 = {T502, T374};
  assign T374 = T375;
  assign T375 = {T494, T376};
  assign T376 = T377;
  assign T377 = {T486, T378};
  assign T378 = T379;
  assign T379 = {T478, T380};
  assign T380 = T381;
  assign T381 = {T470, T382};
  assign T382 = T383;
  assign T383 = {T462, T384};
  assign T384 = T385;
  assign T385 = {T454, T386};
  assign T386 = T387;
  assign T387 = {T446, T388};
  assign T388 = T389;
  assign T389 = {T438, T390};
  assign T390 = T391;
  assign T391 = {T430, T392};
  assign T392 = T393;
  assign T393 = {T422, T394};
  assign T394 = T395;
  assign T395 = {T414, T396};
  assign T396 = T397;
  assign T397 = {T406, T398};
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[4'h9/* 9*/:3'h6/* 6*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[5'h13/* 19*/:4'h9/* 9*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[5'h1f/* 31*/:5'h1d/* 29*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[5'h15/* 21*/:5'h12/* 18*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[6'h2a/* 42*/:6'h20/* 32*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[6'h36/* 54*/:6'h34/* 52*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[6'h21/* 33*/:5'h1e/* 30*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[6'h2d/* 45*/:6'h2a/* 42*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[7'h58/* 88*/:7'h4e/* 78*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[7'h64/* 100*/:7'h62/* 98*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h39/* 57*/:6'h36/* 54*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[7'h6f/* 111*/:7'h65/* 101*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h45/* 69*/:7'h42/* 66*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'h86/* 134*/:7'h7c/* 124*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'h8c/* 140*/:8'h8a/* 138*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'h8f/* 143*/:8'h8d/* 141*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'h92/* 146*/:8'h90/* 144*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h51/* 81*/:7'h4e/* 78*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'h9d/* 157*/:8'h93/* 147*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h53/* 83*/:7'h52/* 82*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'ha0/* 160*/:8'h9e/* 158*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h55/* 85*/:7'h54/* 84*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h57/* 87*/:7'h56/* 86*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'ha6/* 166*/:8'ha4/* 164*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h59/* 89*/:7'h58/* 88*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'ha9/* 169*/:8'ha7/* 167*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hb4/* 180*/:8'haa/* 170*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hb7/* 183*/:8'hb5/* 181*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h61/* 97*/:7'h60/* 96*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hba/* 186*/:8'hb8/* 184*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h63/* 99*/:7'h62/* 98*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'hbd/* 189*/:8'hbb/* 187*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h65/* 101*/:7'h64/* 100*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'hc0/* 192*/:8'hbe/* 190*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h69/* 105*/:7'h66/* 102*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'hcb/* 203*/:8'hc1/* 193*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'hce/* 206*/:8'hcc/* 204*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'hd1/* 209*/:8'hcf/* 207*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'hd4/* 212*/:8'hd2/* 210*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h71/* 113*/:7'h70/* 112*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'hd7/* 215*/:8'hd5/* 213*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'he2/* 226*/:8'hd8/* 216*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h77/* 119*/:7'h76/* 118*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'he5/* 229*/:8'he3/* 227*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'he7/* 231*/:8'he6/* 230*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'he9/* 233*/:8'he8/* 232*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'heb/* 235*/:8'hea/* 234*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h7e/* 126*/:7'h7b/* 123*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'hf6/* 246*/:8'hec/* 236*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h86/* 134*/:8'h83/* 131*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h109/* 265*/:8'hff/* 255*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h11c/* 284*/:9'h112/* 274*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h92/* 146*/:8'h92/* 146*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h96/* 150*/:8'h93/* 147*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h12f/* 303*/:9'h125/* 293*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h135/* 309*/:9'h134/* 308*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h137/* 311*/:9'h136/* 310*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h142/* 322*/:9'h138/* 312*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'ha2/* 162*/:8'ha2/* 162*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h14a/* 330*/:9'h149/* 329*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'ha6/* 166*/:8'ha3/* 163*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h155/* 341*/:9'h14b/* 331*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h157/* 343*/:9'h156/* 342*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h159/* 345*/:9'h158/* 344*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h15b/* 347*/:9'h15a/* 346*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'haa/* 170*/:8'haa/* 170*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h15d/* 349*/:9'h15c/* 348*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hae/* 174*/:8'hab/* 171*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h168/* 360*/:9'h15e/* 350*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h16a/* 362*/:9'h169/* 361*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h16c/* 364*/:9'h16b/* 363*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h16e/* 366*/:9'h16d/* 365*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h170/* 368*/:9'h16f/* 367*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'hb6/* 182*/:8'hb3/* 179*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h17b/* 379*/:9'h171/* 369*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hb7/* 183*/:8'hb7/* 183*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h17d/* 381*/:9'h17c/* 380*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h17f/* 383*/:9'h17e/* 382*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h181/* 385*/:9'h180/* 384*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h183/* 387*/:9'h182/* 386*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'hbe/* 190*/:8'hbb/* 187*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[9'h18e/* 398*/:9'h184/* 388*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hbf/* 191*/:8'hbf/* 191*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[9'h190/* 400*/:9'h18f/* 399*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[9'h192/* 402*/:9'h191/* 401*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[9'h194/* 404*/:9'h193/* 403*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[9'h196/* 406*/:9'h195/* 405*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[9'h1a6/* 422*/:9'h1a4/* 420*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[9'h1a9/* 425*/:9'h1a7/* 423*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[9'h1ac/* 428*/:9'h1aa/* 426*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[8'hd1/* 209*/:8'hce/* 206*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[9'h1b7/* 439*/:9'h1ad/* 429*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[9'h1ba/* 442*/:9'h1b8/* 440*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[8'hd5/* 213*/:8'hd4/* 212*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[9'h1bd/* 445*/:9'h1bb/* 443*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[8'hd7/* 215*/:8'hd6/* 214*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[9'h1c0/* 448*/:9'h1be/* 446*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[9'h1c3/* 451*/:9'h1c1/* 449*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[8'hdd/* 221*/:8'hda/* 218*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[9'h1ce/* 462*/:9'h1c4/* 452*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[9'h1d1/* 465*/:9'h1cf/* 463*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[8'he1/* 225*/:8'he0/* 224*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[9'h1d4/* 468*/:9'h1d2/* 466*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[8'he3/* 227*/:8'he2/* 226*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[9'h1d7/* 471*/:9'h1d5/* 469*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[8'he5/* 229*/:8'he4/* 228*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[9'h1da/* 474*/:9'h1d8/* 472*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[8'he9/* 233*/:8'he6/* 230*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[8'heb/* 235*/:8'hea/* 234*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[9'h1e8/* 488*/:9'h1e6/* 486*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[8'hed/* 237*/:8'hec/* 236*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[9'h1eb/* 491*/:9'h1e9/* 489*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[8'hef/* 239*/:8'hee/* 238*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[9'h1ee/* 494*/:9'h1ec/* 492*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[9'h1f1/* 497*/:9'h1ef/* 495*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[8'hf5/* 245*/:8'hf2/* 242*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[9'h1fc/* 508*/:9'h1f2/* 498*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[8'hf7/* 247*/:8'hf6/* 246*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[9'h1ff/* 511*/:9'h1fd/* 509*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[8'hf9/* 249*/:8'hf8/* 248*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h202/* 514*/:10'h200/* 512*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h205/* 517*/:10'h203/* 515*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[8'hfd/* 253*/:8'hfc/* 252*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h208/* 520*/:10'h206/* 518*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h101/* 257*/:8'hfe/* 254*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h213/* 531*/:10'h209/* 521*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h103/* 259*/:9'h102/* 258*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h216/* 534*/:10'h214/* 532*/];
  assign T1398 = T1399;
  assign T1399 = T1400;
  assign T1400 = T1404[T1401];
  assign T1401 = T1402;
  assign T1402 = T1403;
  assign T1403 = io_chanxy_config[9'h105/* 261*/:9'h104/* 260*/];
  assign T1404 = T1405;
  assign T1405 = io_chanxy_in[10'h219/* 537*/:10'h217/* 535*/];
  assign T1406 = T1407;
  assign T1407 = T1408;
  assign T1408 = T1412[T1409];
  assign T1409 = T1410;
  assign T1410 = T1411;
  assign T1411 = io_chanxy_config[9'h107/* 263*/:9'h106/* 262*/];
  assign T1412 = T1413;
  assign T1413 = io_chanxy_in[10'h21c/* 540*/:10'h21a/* 538*/];
  assign T1414 = T1415;
  assign T1415 = T1416;
  assign T1416 = T1420[T1417];
  assign T1417 = T1418;
  assign T1418 = T1419;
  assign T1419 = io_chanxy_config[9'h109/* 265*/:9'h108/* 264*/];
  assign T1420 = T1421;
  assign T1421 = io_chanxy_in[10'h21f/* 543*/:10'h21d/* 541*/];
  assign T1422 = T1423;
  assign T1423 = T1424;
  assign T1424 = T1428[T1425];
  assign T1425 = T1426;
  assign T1426 = T1427;
  assign T1427 = io_chanxy_config[9'h10d/* 269*/:9'h10a/* 266*/];
  assign T1428 = T1429;
  assign T1429 = io_chanxy_in[10'h22a/* 554*/:10'h220/* 544*/];
  assign T1430 = T1431;
  assign T1431 = T1432;
  assign T1432 = T1436[T1433];
  assign T1433 = T1434;
  assign T1434 = T1435;
  assign T1435 = io_chanxy_config[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T1436 = T1437;
  assign T1437 = io_chanxy_in[10'h22d/* 557*/:10'h22b/* 555*/];
  assign T1438 = T1439;
  assign T1439 = T1440;
  assign T1440 = T1444[T1441];
  assign T1441 = T1442;
  assign T1442 = T1443;
  assign T1443 = io_chanxy_config[9'h111/* 273*/:9'h110/* 272*/];
  assign T1444 = T1445;
  assign T1445 = io_chanxy_in[10'h230/* 560*/:10'h22e/* 558*/];
  assign T1446 = T1447;
  assign T1447 = T1448;
  assign T1448 = T1452[T1449];
  assign T1449 = T1450;
  assign T1450 = T1451;
  assign T1451 = io_chanxy_config[9'h113/* 275*/:9'h112/* 274*/];
  assign T1452 = T1453;
  assign T1453 = io_chanxy_in[10'h233/* 563*/:10'h231/* 561*/];
  assign T1454 = T1455;
  assign T1455 = T1456;
  assign T1456 = T1460[T1457];
  assign T1457 = T1458;
  assign T1458 = T1459;
  assign T1459 = io_chanxy_config[9'h115/* 277*/:9'h114/* 276*/];
  assign T1460 = T1461;
  assign T1461 = io_chanxy_in[10'h236/* 566*/:10'h234/* 564*/];
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_chanxy_config[9'h119/* 281*/:9'h116/* 278*/];
  assign T1468 = T1469;
  assign T1469 = io_chanxy_in[10'h241/* 577*/:10'h237/* 567*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_chanxy_config[9'h11b/* 283*/:9'h11a/* 282*/];
  assign T1476 = T1477;
  assign T1477 = io_chanxy_in[10'h244/* 580*/:10'h242/* 578*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_chanxy_config[9'h11d/* 285*/:9'h11c/* 284*/];
  assign T1484 = T1485;
  assign T1485 = io_chanxy_in[10'h247/* 583*/:10'h245/* 581*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_chanxy_config[9'h11f/* 287*/:9'h11e/* 286*/];
  assign T1492 = T1493;
  assign T1493 = io_chanxy_in[10'h24a/* 586*/:10'h248/* 584*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_chanxy_config[9'h121/* 289*/:9'h120/* 288*/];
  assign T1500 = T1501;
  assign T1501 = io_chanxy_in[10'h24d/* 589*/:10'h24b/* 587*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_chanxy_config[9'h125/* 293*/:9'h122/* 290*/];
  assign T1508 = T1509;
  assign T1509 = io_chanxy_in[10'h258/* 600*/:10'h24e/* 590*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_chanxy_config[9'h127/* 295*/:9'h126/* 294*/];
  assign T1516 = T1517;
  assign T1517 = io_chanxy_in[10'h25b/* 603*/:10'h259/* 601*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_chanxy_config[9'h129/* 297*/:9'h128/* 296*/];
  assign T1524 = T1525;
  assign T1525 = io_chanxy_in[10'h25e/* 606*/:10'h25c/* 604*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_chanxy_config[9'h12b/* 299*/:9'h12a/* 298*/];
  assign T1532 = T1533;
  assign T1533 = io_chanxy_in[10'h261/* 609*/:10'h25f/* 607*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_chanxy_config[9'h12d/* 301*/:9'h12c/* 300*/];
  assign T1540 = T1541;
  assign T1541 = io_chanxy_in[10'h264/* 612*/:10'h262/* 610*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_chanxy_config[9'h131/* 305*/:9'h12e/* 302*/];
  assign T1548 = T1549;
  assign T1549 = io_chanxy_in[10'h26f/* 623*/:10'h265/* 613*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_chanxy_config[9'h133/* 307*/:9'h132/* 306*/];
  assign T1556 = T1557;
  assign T1557 = io_chanxy_in[10'h272/* 626*/:10'h270/* 624*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_chanxy_config[9'h135/* 309*/:9'h134/* 308*/];
  assign T1564 = T1565;
  assign T1565 = io_chanxy_in[10'h275/* 629*/:10'h273/* 627*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_chanxy_config[9'h137/* 311*/:9'h136/* 310*/];
  assign T1572 = T1573;
  assign T1573 = io_chanxy_in[10'h278/* 632*/:10'h276/* 630*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_chanxy_config[9'h139/* 313*/:9'h138/* 312*/];
  assign T1580 = T1581;
  assign T1581 = io_chanxy_in[10'h27b/* 635*/:10'h279/* 633*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_chanxy_config[9'h13d/* 317*/:9'h13a/* 314*/];
  assign T1588 = T1589;
  assign T1589 = io_chanxy_in[10'h286/* 646*/:10'h27c/* 636*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_chanxy_config[9'h13f/* 319*/:9'h13e/* 318*/];
  assign T1596 = T1597;
  assign T1597 = io_chanxy_in[10'h289/* 649*/:10'h287/* 647*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_chanxy_config[9'h140/* 320*/:9'h140/* 320*/];
  assign T1604 = T1605;
  assign T1605 = io_chanxy_in[10'h28b/* 651*/:10'h28a/* 650*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_chanxy_config[9'h141/* 321*/:9'h141/* 321*/];
  assign T1612 = T1613;
  assign T1613 = io_chanxy_in[10'h28d/* 653*/:10'h28c/* 652*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_chanxy_config[9'h142/* 322*/:9'h142/* 322*/];
  assign T1620 = T1621;
  assign T1621 = io_chanxy_in[10'h28f/* 655*/:10'h28e/* 654*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_chanxy_config[9'h146/* 326*/:9'h143/* 323*/];
  assign T1628 = T1629;
  assign T1629 = io_chanxy_in[10'h29a/* 666*/:10'h290/* 656*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_chanxy_config[9'h147/* 327*/:9'h147/* 327*/];
  assign T1636 = T1637;
  assign T1637 = io_chanxy_in[10'h29c/* 668*/:10'h29b/* 667*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_chanxy_config[9'h148/* 328*/:9'h148/* 328*/];
  assign T1644 = T1645;
  assign T1645 = io_chanxy_in[10'h29e/* 670*/:10'h29d/* 669*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1652 = T1653;
  assign T1653 = io_chanxy_in[10'h2a0/* 672*/:10'h29f/* 671*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_chanxy_config[9'h14a/* 330*/:9'h14a/* 330*/];
  assign T1660 = T1661;
  assign T1661 = io_chanxy_in[10'h2a2/* 674*/:10'h2a1/* 673*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_chanxy_config[9'h14e/* 334*/:9'h14b/* 331*/];
  assign T1668 = T1669;
  assign T1669 = io_chanxy_in[10'h2ad/* 685*/:10'h2a3/* 675*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_chanxy_config[9'h14f/* 335*/:9'h14f/* 335*/];
  assign T1676 = T1677;
  assign T1677 = io_chanxy_in[10'h2af/* 687*/:10'h2ae/* 686*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_chanxy_config[9'h150/* 336*/:9'h150/* 336*/];
  assign T1684 = T1685;
  assign T1685 = io_chanxy_in[10'h2b1/* 689*/:10'h2b0/* 688*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_chanxy_config[9'h151/* 337*/:9'h151/* 337*/];
  assign T1692 = T1693;
  assign T1693 = io_chanxy_in[10'h2b3/* 691*/:10'h2b2/* 690*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_chanxy_config[9'h152/* 338*/:9'h152/* 338*/];
  assign T1700 = T1701;
  assign T1701 = io_chanxy_in[10'h2b5/* 693*/:10'h2b4/* 692*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_chanxy_config[9'h156/* 342*/:9'h153/* 339*/];
  assign T1708 = T1709;
  assign T1709 = io_chanxy_in[10'h2c0/* 704*/:10'h2b6/* 694*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_chanxy_config[9'h157/* 343*/:9'h157/* 343*/];
  assign T1716 = T1717;
  assign T1717 = io_chanxy_in[10'h2c2/* 706*/:10'h2c1/* 705*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1724 = T1725;
  assign T1725 = io_chanxy_in[10'h2c4/* 708*/:10'h2c3/* 707*/];
  assign T1726 = T1727;
  assign T1727 = T1728;
  assign T1728 = T1732[T1729];
  assign T1729 = T1730;
  assign T1730 = T1731;
  assign T1731 = io_chanxy_config[9'h159/* 345*/:9'h159/* 345*/];
  assign T1732 = T1733;
  assign T1733 = io_chanxy_in[10'h2c6/* 710*/:10'h2c5/* 709*/];
  assign T1734 = T1735;
  assign T1735 = T1736;
  assign T1736 = T1740[T1737];
  assign T1737 = T1738;
  assign T1738 = T1739;
  assign T1739 = io_chanxy_config[9'h15a/* 346*/:9'h15a/* 346*/];
  assign T1740 = T1741;
  assign T1741 = io_chanxy_in[10'h2c8/* 712*/:10'h2c7/* 711*/];
  assign T1742 = T1743;
  assign T1743 = T1744;
  assign T1744 = T1748[T1745];
  assign T1745 = T1746;
  assign T1746 = T1747;
  assign T1747 = io_chanxy_config[9'h15e/* 350*/:9'h15b/* 347*/];
  assign T1748 = T1749;
  assign T1749 = io_chanxy_in[10'h2d3/* 723*/:10'h2c9/* 713*/];
  assign T1750 = T1751;
  assign T1751 = T1752;
  assign T1752 = T1756[T1753];
  assign T1753 = T1754;
  assign T1754 = T1755;
  assign T1755 = io_chanxy_config[9'h15f/* 351*/:9'h15f/* 351*/];
  assign T1756 = T1757;
  assign T1757 = io_chanxy_in[10'h2d5/* 725*/:10'h2d4/* 724*/];
  assign T1758 = T1759;
  assign T1759 = T1760;
  assign T1760 = T1764[T1761];
  assign T1761 = T1762;
  assign T1762 = T1763;
  assign T1763 = io_chanxy_config[9'h160/* 352*/:9'h160/* 352*/];
  assign T1764 = T1765;
  assign T1765 = io_chanxy_in[10'h2d7/* 727*/:10'h2d6/* 726*/];
  assign T1766 = T1767;
  assign T1767 = T1768;
  assign T1768 = T1772[T1769];
  assign T1769 = T1770;
  assign T1770 = T1771;
  assign T1771 = io_chanxy_config[9'h161/* 353*/:9'h161/* 353*/];
  assign T1772 = T1773;
  assign T1773 = io_chanxy_in[10'h2d9/* 729*/:10'h2d8/* 728*/];
  assign T1774 = T1775;
  assign T1775 = T1776;
  assign T1776 = T1780[T1777];
  assign T1777 = T1778;
  assign T1778 = T1779;
  assign T1779 = io_chanxy_config[9'h162/* 354*/:9'h162/* 354*/];
  assign T1780 = T1781;
  assign T1781 = io_chanxy_in[10'h2db/* 731*/:10'h2da/* 730*/];
  assign T1782 = T1783;
  assign T1783 = T1784;
  assign T1784 = T1788[T1785];
  assign T1785 = T1786;
  assign T1786 = T1787;
  assign T1787 = io_chanxy_config[9'h166/* 358*/:9'h163/* 355*/];
  assign T1788 = T1789;
  assign T1789 = io_chanxy_in[10'h2e6/* 742*/:10'h2dc/* 732*/];
  assign T1790 = T1791;
  assign T1791 = T1792;
  assign T1792 = T1796[T1793];
  assign T1793 = T1794;
  assign T1794 = T1795;
  assign T1795 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1796 = T1797;
  assign T1797 = io_chanxy_in[10'h2e8/* 744*/:10'h2e7/* 743*/];
  assign T1798 = T1799;
  assign T1799 = T1800;
  assign T1800 = T1804[T1801];
  assign T1801 = T1802;
  assign T1802 = T1803;
  assign T1803 = io_chanxy_config[9'h168/* 360*/:9'h168/* 360*/];
  assign T1804 = T1805;
  assign T1805 = io_chanxy_in[10'h2ea/* 746*/:10'h2e9/* 745*/];
  assign T1806 = T1807;
  assign T1807 = T1808;
  assign T1808 = T1812[T1809];
  assign T1809 = T1810;
  assign T1810 = T1811;
  assign T1811 = io_chanxy_config[9'h169/* 361*/:9'h169/* 361*/];
  assign T1812 = T1813;
  assign T1813 = io_chanxy_in[10'h2ec/* 748*/:10'h2eb/* 747*/];
  assign T1814 = T1815;
  assign T1815 = T1816;
  assign T1816 = T1820[T1817];
  assign T1817 = T1818;
  assign T1818 = T1819;
  assign T1819 = io_chanxy_config[9'h16a/* 362*/:9'h16a/* 362*/];
  assign T1820 = T1821;
  assign T1821 = io_chanxy_in[10'h2ee/* 750*/:10'h2ed/* 749*/];
  assign T1822 = T1823;
  assign T1823 = T1824;
  assign T1824 = T1828[T1825];
  assign T1825 = T1826;
  assign T1826 = T1827;
  assign T1827 = io_chanxy_config[9'h16e/* 366*/:9'h16b/* 363*/];
  assign T1828 = T1829;
  assign T1829 = io_chanxy_in[10'h2f9/* 761*/:10'h2ef/* 751*/];
  assign T1830 = T1831;
  assign T1831 = T1832;
  assign T1832 = T1836[T1833];
  assign T1833 = T1834;
  assign T1834 = T1835;
  assign T1835 = io_chanxy_config[9'h16f/* 367*/:9'h16f/* 367*/];
  assign T1836 = T1837;
  assign T1837 = io_chanxy_in[10'h2fb/* 763*/:10'h2fa/* 762*/];
  assign T1838 = T1839;
  assign T1839 = T1840;
  assign T1840 = T1844[T1841];
  assign T1841 = T1842;
  assign T1842 = T1843;
  assign T1843 = io_chanxy_config[9'h170/* 368*/:9'h170/* 368*/];
  assign T1844 = T1845;
  assign T1845 = io_chanxy_in[10'h2fd/* 765*/:10'h2fc/* 764*/];
  assign T1846 = T1847;
  assign T1847 = T1848;
  assign T1848 = T1852[T1849];
  assign T1849 = T1850;
  assign T1850 = T1851;
  assign T1851 = io_chanxy_config[9'h171/* 369*/:9'h171/* 369*/];
  assign T1852 = T1853;
  assign T1853 = io_chanxy_in[10'h2ff/* 767*/:10'h2fe/* 766*/];
  assign T1854 = T1855;
  assign T1855 = T1856;
  assign T1856 = T1860[T1857];
  assign T1857 = T1858;
  assign T1858 = T1859;
  assign T1859 = io_chanxy_config[9'h172/* 370*/:9'h172/* 370*/];
  assign T1860 = T1861;
  assign T1861 = io_chanxy_in[10'h301/* 769*/:10'h300/* 768*/];
  assign T1862 = T1863;
  assign T1863 = T1864;
  assign T1864 = T1868[T1865];
  assign T1865 = T1866;
  assign T1866 = T1867;
  assign T1867 = io_chanxy_config[9'h176/* 374*/:9'h173/* 371*/];
  assign T1868 = T1869;
  assign T1869 = io_chanxy_in[10'h30c/* 780*/:10'h302/* 770*/];
  assign T1870 = T1871;
  assign T1871 = T1872;
  assign T1872 = T1876[T1873];
  assign T1873 = T1874;
  assign T1874 = T1875;
  assign T1875 = io_chanxy_config[9'h177/* 375*/:9'h177/* 375*/];
  assign T1876 = T1877;
  assign T1877 = io_chanxy_in[10'h30e/* 782*/:10'h30d/* 781*/];
  assign T1878 = T1879;
  assign T1879 = T1880;
  assign T1880 = T1884[T1881];
  assign T1881 = T1882;
  assign T1882 = T1883;
  assign T1883 = io_chanxy_config[9'h178/* 376*/:9'h178/* 376*/];
  assign T1884 = T1885;
  assign T1885 = io_chanxy_in[10'h310/* 784*/:10'h30f/* 783*/];
  assign T1886 = T1887;
  assign T1887 = T1888;
  assign T1888 = T1892[T1889];
  assign T1889 = T1890;
  assign T1890 = T1891;
  assign T1891 = io_chanxy_config[9'h179/* 377*/:9'h179/* 377*/];
  assign T1892 = T1893;
  assign T1893 = io_chanxy_in[10'h312/* 786*/:10'h311/* 785*/];
  assign T1894 = T1895;
  assign T1895 = T1896;
  assign T1896 = T1900[T1897];
  assign T1897 = T1898;
  assign T1898 = T1899;
  assign T1899 = io_chanxy_config[9'h17a/* 378*/:9'h17a/* 378*/];
  assign T1900 = T1901;
  assign T1901 = io_chanxy_in[10'h314/* 788*/:10'h313/* 787*/];
  assign T1902 = T1903;
  assign T1903 = T1904;
  assign T1904 = T1908[T1905];
  assign T1905 = T1906;
  assign T1906 = T1907;
  assign T1907 = io_chanxy_config[9'h17e/* 382*/:9'h17b/* 379*/];
  assign T1908 = T1909;
  assign T1909 = io_chanxy_in[10'h31f/* 799*/:10'h315/* 789*/];
  assign T1910 = T1911;
  assign T1911 = T1912;
  assign T1912 = T1916[T1913];
  assign T1913 = T1914;
  assign T1914 = T1915;
  assign T1915 = io_chanxy_config[9'h17f/* 383*/:9'h17f/* 383*/];
  assign T1916 = T1917;
  assign T1917 = io_chanxy_in[10'h321/* 801*/:10'h320/* 800*/];
  assign T1918 = T1919;
  assign T1919 = T1920;
  assign T1920 = T1924[T1921];
  assign T1921 = T1922;
  assign T1922 = T1923;
  assign T1923 = io_chanxy_config[9'h180/* 384*/:9'h180/* 384*/];
  assign T1924 = T1925;
  assign T1925 = io_chanxy_in[10'h323/* 803*/:10'h322/* 802*/];
  assign T1926 = T1927;
  assign T1927 = T1928;
  assign T1928 = T1932[T1929];
  assign T1929 = T1930;
  assign T1930 = T1931;
  assign T1931 = io_chanxy_config[9'h181/* 385*/:9'h181/* 385*/];
  assign T1932 = T1933;
  assign T1933 = io_chanxy_in[10'h325/* 805*/:10'h324/* 804*/];
  assign T1934 = T1935;
  assign T1935 = T1936;
  assign T1936 = T1940[T1937];
  assign T1937 = T1938;
  assign T1938 = T1939;
  assign T1939 = io_chanxy_config[9'h182/* 386*/:9'h182/* 386*/];
  assign T1940 = T1941;
  assign T1941 = io_chanxy_in[10'h327/* 807*/:10'h326/* 806*/];
  assign T1942 = T1943;
  assign T1943 = T1944;
  assign T1944 = T1948[T1945];
  assign T1945 = T1946;
  assign T1946 = T1947;
  assign T1947 = io_chanxy_config[9'h186/* 390*/:9'h183/* 387*/];
  assign T1948 = T1949;
  assign T1949 = io_chanxy_in[10'h332/* 818*/:10'h328/* 808*/];
  assign T1950 = T1951;
  assign T1951 = T1952;
  assign T1952 = T1956[T1953];
  assign T1953 = T1954;
  assign T1954 = T1955;
  assign T1955 = io_chanxy_config[9'h187/* 391*/:9'h187/* 391*/];
  assign T1956 = T1957;
  assign T1957 = io_chanxy_in[10'h334/* 820*/:10'h333/* 819*/];
  assign T1958 = T1959;
  assign T1959 = T1960;
  assign T1960 = T1964[T1961];
  assign T1961 = T1962;
  assign T1962 = T1963;
  assign T1963 = io_chanxy_config[9'h188/* 392*/:9'h188/* 392*/];
  assign T1964 = T1965;
  assign T1965 = io_chanxy_in[10'h336/* 822*/:10'h335/* 821*/];
  assign T1966 = T1967;
  assign T1967 = T1968;
  assign T1968 = T1972[T1969];
  assign T1969 = T1970;
  assign T1970 = T1971;
  assign T1971 = io_chanxy_config[9'h189/* 393*/:9'h189/* 393*/];
  assign T1972 = T1973;
  assign T1973 = io_chanxy_in[10'h338/* 824*/:10'h337/* 823*/];
  assign T1974 = T1975;
  assign T1975 = T1976;
  assign T1976 = T1980[T1977];
  assign T1977 = T1978;
  assign T1978 = T1979;
  assign T1979 = io_chanxy_config[9'h18a/* 394*/:9'h18a/* 394*/];
  assign T1980 = T1981;
  assign T1981 = io_chanxy_in[10'h33a/* 826*/:10'h339/* 825*/];
  assign T1982 = T1983;
  assign T1983 = T1984;
  assign T1984 = T1988[T1985];
  assign T1985 = T1986;
  assign T1986 = T1987;
  assign T1987 = io_chanxy_config[9'h18e/* 398*/:9'h18b/* 395*/];
  assign T1988 = T1989;
  assign T1989 = io_chanxy_in[10'h345/* 837*/:10'h33b/* 827*/];
  assign T1990 = T1991;
  assign T1991 = T1992;
  assign T1992 = T1996[T1993];
  assign T1993 = T1994;
  assign T1994 = T1995;
  assign T1995 = io_chanxy_config[9'h18f/* 399*/:9'h18f/* 399*/];
  assign T1996 = T1997;
  assign T1997 = io_chanxy_in[10'h347/* 839*/:10'h346/* 838*/];
  assign io_ipin_out = T1998;
  assign T1998 = T1999;
  assign T1999 = {T2318, T2000};
  assign T2000 = T2001;
  assign T2001 = {T2310, T2002};
  assign T2002 = T2003;
  assign T2003 = {T2302, T2004};
  assign T2004 = T2005;
  assign T2005 = {T2294, T2006};
  assign T2006 = T2007;
  assign T2007 = {T2286, T2008};
  assign T2008 = T2009;
  assign T2009 = {T2278, T2010};
  assign T2010 = T2011;
  assign T2011 = {T2270, T2012};
  assign T2012 = T2013;
  assign T2013 = {T2262, T2014};
  assign T2014 = T2015;
  assign T2015 = {T2254, T2016};
  assign T2016 = T2017;
  assign T2017 = {T2246, T2018};
  assign T2018 = T2019;
  assign T2019 = {T2238, T2020};
  assign T2020 = T2021;
  assign T2021 = {T2230, T2022};
  assign T2022 = T2023;
  assign T2023 = {T2222, T2024};
  assign T2024 = T2025;
  assign T2025 = {T2214, T2026};
  assign T2026 = T2027;
  assign T2027 = {T2206, T2028};
  assign T2028 = T2029;
  assign T2029 = {T2198, T2030};
  assign T2030 = T2031;
  assign T2031 = {T2190, T2032};
  assign T2032 = T2033;
  assign T2033 = {T2182, T2034};
  assign T2034 = T2035;
  assign T2035 = {T2174, T2036};
  assign T2036 = T2037;
  assign T2037 = {T2166, T2038};
  assign T2038 = T2039;
  assign T2039 = {T2158, T2040};
  assign T2040 = T2041;
  assign T2041 = {T2150, T2042};
  assign T2042 = T2043;
  assign T2043 = {T2142, T2044};
  assign T2044 = T2045;
  assign T2045 = {T2134, T2046};
  assign T2046 = T2047;
  assign T2047 = {T2126, T2048};
  assign T2048 = T2049;
  assign T2049 = {T2118, T2050};
  assign T2050 = T2051;
  assign T2051 = {T2110, T2052};
  assign T2052 = T2053;
  assign T2053 = {T2102, T2054};
  assign T2054 = T2055;
  assign T2055 = {T2094, T2056};
  assign T2056 = T2057;
  assign T2057 = {T2086, T2058};
  assign T2058 = T2059;
  assign T2059 = {T2078, T2060};
  assign T2060 = T2061;
  assign T2061 = {T2070, T2062};
  assign T2062 = T2063;
  assign T2063 = T2064;
  assign T2064 = T2068[T2065];
  assign T2065 = T2066;
  assign T2066 = T2067;
  assign T2067 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T2068 = T2069;
  assign T2069 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T2070 = T2071;
  assign T2071 = T2072;
  assign T2072 = T2076[T2073];
  assign T2073 = T2074;
  assign T2074 = T2075;
  assign T2075 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T2076 = T2077;
  assign T2077 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T2078 = T2079;
  assign T2079 = T2080;
  assign T2080 = T2084[T2081];
  assign T2081 = T2082;
  assign T2082 = T2083;
  assign T2083 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T2084 = T2085;
  assign T2085 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T2086 = T2087;
  assign T2087 = T2088;
  assign T2088 = T2092[T2089];
  assign T2089 = T2090;
  assign T2090 = T2091;
  assign T2091 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T2092 = T2093;
  assign T2093 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T2094 = T2095;
  assign T2095 = T2096;
  assign T2096 = T2100[T2097];
  assign T2097 = T2098;
  assign T2098 = T2099;
  assign T2099 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T2100 = T2101;
  assign T2101 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T2102 = T2103;
  assign T2103 = T2104;
  assign T2104 = T2108[T2105];
  assign T2105 = T2106;
  assign T2106 = T2107;
  assign T2107 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T2108 = T2109;
  assign T2109 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T2110 = T2111;
  assign T2111 = T2112;
  assign T2112 = T2116[T2113];
  assign T2113 = T2114;
  assign T2114 = T2115;
  assign T2115 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T2116 = T2117;
  assign T2117 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T2118 = T2119;
  assign T2119 = T2120;
  assign T2120 = T2124[T2121];
  assign T2121 = T2122;
  assign T2122 = T2123;
  assign T2123 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T2124 = T2125;
  assign T2125 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T2126 = T2127;
  assign T2127 = T2128;
  assign T2128 = T2132[T2129];
  assign T2129 = T2130;
  assign T2130 = T2131;
  assign T2131 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T2132 = T2133;
  assign T2133 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T2134 = T2135;
  assign T2135 = T2136;
  assign T2136 = T2140[T2137];
  assign T2137 = T2138;
  assign T2138 = T2139;
  assign T2139 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T2140 = T2141;
  assign T2141 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T2142 = T2143;
  assign T2143 = T2144;
  assign T2144 = T2148[T2145];
  assign T2145 = T2146;
  assign T2146 = T2147;
  assign T2147 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T2148 = T2149;
  assign T2149 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T2150 = T2151;
  assign T2151 = T2152;
  assign T2152 = T2156[T2153];
  assign T2153 = T2154;
  assign T2154 = T2155;
  assign T2155 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T2156 = T2157;
  assign T2157 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T2158 = T2159;
  assign T2159 = T2160;
  assign T2160 = T2164[T2161];
  assign T2161 = T2162;
  assign T2162 = T2163;
  assign T2163 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T2164 = T2165;
  assign T2165 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T2166 = T2167;
  assign T2167 = T2168;
  assign T2168 = T2172[T2169];
  assign T2169 = T2170;
  assign T2170 = T2171;
  assign T2171 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T2172 = T2173;
  assign T2173 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T2174 = T2175;
  assign T2175 = T2176;
  assign T2176 = T2180[T2177];
  assign T2177 = T2178;
  assign T2178 = T2179;
  assign T2179 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T2180 = T2181;
  assign T2181 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T2182 = T2183;
  assign T2183 = T2184;
  assign T2184 = T2188[T2185];
  assign T2185 = T2186;
  assign T2186 = T2187;
  assign T2187 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T2188 = T2189;
  assign T2189 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T2190 = T2191;
  assign T2191 = T2192;
  assign T2192 = T2196[T2193];
  assign T2193 = T2194;
  assign T2194 = T2195;
  assign T2195 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T2196 = T2197;
  assign T2197 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T2198 = T2199;
  assign T2199 = T2200;
  assign T2200 = T2204[T2201];
  assign T2201 = T2202;
  assign T2202 = T2203;
  assign T2203 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T2204 = T2205;
  assign T2205 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T2206 = T2207;
  assign T2207 = T2208;
  assign T2208 = T2212[T2209];
  assign T2209 = T2210;
  assign T2210 = T2211;
  assign T2211 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T2212 = T2213;
  assign T2213 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T2214 = T2215;
  assign T2215 = T2216;
  assign T2216 = T2220[T2217];
  assign T2217 = T2218;
  assign T2218 = T2219;
  assign T2219 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T2220 = T2221;
  assign T2221 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T2222 = T2223;
  assign T2223 = T2224;
  assign T2224 = T2228[T2225];
  assign T2225 = T2226;
  assign T2226 = T2227;
  assign T2227 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T2228 = T2229;
  assign T2229 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T2230 = T2231;
  assign T2231 = T2232;
  assign T2232 = T2236[T2233];
  assign T2233 = T2234;
  assign T2234 = T2235;
  assign T2235 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T2236 = T2237;
  assign T2237 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T2238 = T2239;
  assign T2239 = T2240;
  assign T2240 = T2244[T2241];
  assign T2241 = T2242;
  assign T2242 = T2243;
  assign T2243 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T2244 = T2245;
  assign T2245 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T2246 = T2247;
  assign T2247 = T2248;
  assign T2248 = T2252[T2249];
  assign T2249 = T2250;
  assign T2250 = T2251;
  assign T2251 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T2252 = T2253;
  assign T2253 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T2254 = T2255;
  assign T2255 = T2256;
  assign T2256 = T2260[T2257];
  assign T2257 = T2258;
  assign T2258 = T2259;
  assign T2259 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T2260 = T2261;
  assign T2261 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T2262 = T2263;
  assign T2263 = T2264;
  assign T2264 = T2268[T2265];
  assign T2265 = T2266;
  assign T2266 = T2267;
  assign T2267 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T2268 = T2269;
  assign T2269 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T2270 = T2271;
  assign T2271 = T2272;
  assign T2272 = T2276[T2273];
  assign T2273 = T2274;
  assign T2274 = T2275;
  assign T2275 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T2276 = T2277;
  assign T2277 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T2278 = T2279;
  assign T2279 = T2280;
  assign T2280 = T2284[T2281];
  assign T2281 = T2282;
  assign T2282 = T2283;
  assign T2283 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T2284 = T2285;
  assign T2285 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T2286 = T2287;
  assign T2287 = T2288;
  assign T2288 = T2292[T2289];
  assign T2289 = T2290;
  assign T2290 = T2291;
  assign T2291 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T2292 = T2293;
  assign T2293 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T2294 = T2295;
  assign T2295 = T2296;
  assign T2296 = T2300[T2297];
  assign T2297 = T2298;
  assign T2298 = T2299;
  assign T2299 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T2300 = T2301;
  assign T2301 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T2302 = T2303;
  assign T2303 = T2304;
  assign T2304 = T2308[T2305];
  assign T2305 = T2306;
  assign T2306 = T2307;
  assign T2307 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T2308 = T2309;
  assign T2309 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T2310 = T2311;
  assign T2311 = T2312;
  assign T2312 = T2316[T2313];
  assign T2313 = T2314;
  assign T2314 = T2315;
  assign T2315 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T2316 = T2317;
  assign T2317 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T2318 = T2319;
  assign T2319 = T2320;
  assign T2320 = T2324[T2321];
  assign T2321 = T2322;
  assign T2322 = T2323;
  assign T2323 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T2324 = T2325;
  assign T2325 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_0(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [48:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [839:0] io_chanxy_in,
    output[199:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[399:0] T0;
  wire[1567:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[199:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h605/* 1541*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_49 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


module sbcb_sp_1(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[1:0] T281;
  wire[1:0] T282;
  wire[1:0] T283;
  wire[2:0] T284;
  wire[2:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[1:0] T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[1:0] T297;
  wire[1:0] T298;
  wire[1:0] T299;
  wire[2:0] T300;
  wire[2:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[1:0] T305;
  wire[1:0] T306;
  wire[1:0] T307;
  wire[2:0] T308;
  wire[2:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[10:0] T316;
  wire[10:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[1:0] T321;
  wire[1:0] T322;
  wire[1:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[1:0] T330;
  wire[1:0] T331;
  wire[2:0] T332;
  wire[2:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[1:0] T337;
  wire[1:0] T338;
  wire[1:0] T339;
  wire[2:0] T340;
  wire[2:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[1:0] T345;
  wire[1:0] T346;
  wire[1:0] T347;
  wire[2:0] T348;
  wire[2:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[10:0] T356;
  wire[10:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[1:0] T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[2:0] T364;
  wire[2:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[2:0] T372;
  wire[2:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[2:0] T380;
  wire[2:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[1:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[2:0] T388;
  wire[2:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[10:0] T396;
  wire[10:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire[1:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[1:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire[2:0] T412;
  wire[2:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[1:0] T417;
  wire[1:0] T418;
  wire[1:0] T419;
  wire[2:0] T420;
  wire[2:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T426;
  wire[1:0] T427;
  wire[2:0] T428;
  wire[2:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[3:0] T433;
  wire[3:0] T434;
  wire[3:0] T435;
  wire[10:0] T436;
  wire[10:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[1:0] T449;
  wire[1:0] T450;
  wire[1:0] T451;
  wire[2:0] T452;
  wire[2:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[1:0] T457;
  wire[1:0] T458;
  wire[1:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[1:0] T467;
  wire[2:0] T468;
  wire[2:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[3:0] T473;
  wire[3:0] T474;
  wire[3:0] T475;
  wire[10:0] T476;
  wire[10:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[1:0] T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[2:0] T484;
  wire[2:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[1:0] T489;
  wire[1:0] T490;
  wire[1:0] T491;
  wire[2:0] T492;
  wire[2:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[2:0] T500;
  wire[2:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[1:0] T505;
  wire[1:0] T506;
  wire[1:0] T507;
  wire[2:0] T508;
  wire[2:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[10:0] T516;
  wire[10:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire[1:0] T523;
  wire[2:0] T524;
  wire[2:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[1:0] T529;
  wire[1:0] T530;
  wire[1:0] T531;
  wire[2:0] T532;
  wire[2:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[1:0] T537;
  wire[1:0] T538;
  wire[1:0] T539;
  wire[2:0] T540;
  wire[2:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[1:0] T545;
  wire[1:0] T546;
  wire[1:0] T547;
  wire[2:0] T548;
  wire[2:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[3:0] T553;
  wire[3:0] T554;
  wire[3:0] T555;
  wire[10:0] T556;
  wire[10:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[1:0] T561;
  wire[1:0] T562;
  wire[1:0] T563;
  wire[2:0] T564;
  wire[2:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[1:0] T569;
  wire[1:0] T570;
  wire[1:0] T571;
  wire[2:0] T572;
  wire[2:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[1:0] T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[2:0] T580;
  wire[2:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[1:0] T585;
  wire[1:0] T586;
  wire[1:0] T587;
  wire[2:0] T588;
  wire[2:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[3:0] T593;
  wire[3:0] T594;
  wire[3:0] T595;
  wire[10:0] T596;
  wire[10:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[3:0] T633;
  wire[3:0] T634;
  wire[3:0] T635;
  wire[10:0] T636;
  wire[10:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[3:0] T673;
  wire[3:0] T674;
  wire[3:0] T675;
  wire[10:0] T676;
  wire[10:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[3:0] T713;
  wire[3:0] T714;
  wire[3:0] T715;
  wire[10:0] T716;
  wire[10:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[3:0] T753;
  wire[3:0] T754;
  wire[3:0] T755;
  wire[10:0] T756;
  wire[10:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire[1:0] T780;
  wire[1:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[3:0] T793;
  wire[3:0] T794;
  wire[3:0] T795;
  wire[10:0] T796;
  wire[10:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[3:0] T833;
  wire[3:0] T834;
  wire[3:0] T835;
  wire[10:0] T836;
  wire[10:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T875;
  wire[10:0] T876;
  wire[10:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[3:0] T913;
  wire[3:0] T914;
  wire[3:0] T915;
  wire[10:0] T916;
  wire[10:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire[1:0] T940;
  wire[1:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[3:0] T953;
  wire[3:0] T954;
  wire[3:0] T955;
  wire[10:0] T956;
  wire[10:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[3:0] T993;
  wire[3:0] T994;
  wire[3:0] T995;
  wire[10:0] T996;
  wire[10:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[3:0] T1033;
  wire[3:0] T1034;
  wire[3:0] T1035;
  wire[10:0] T1036;
  wire[10:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire[3:0] T1073;
  wire[3:0] T1074;
  wire[3:0] T1075;
  wire[10:0] T1076;
  wire[10:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire[3:0] T1081;
  wire[3:0] T1082;
  wire[3:0] T1083;
  wire[10:0] T1084;
  wire[10:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[10:0] T1092;
  wire[10:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[10:0] T1100;
  wire[10:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[10:0] T1108;
  wire[10:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[10:0] T1116;
  wire[10:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[10:0] T1124;
  wire[10:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[10:0] T1132;
  wire[10:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[10:0] T1140;
  wire[10:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[10:0] T1148;
  wire[10:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[10:0] T1156;
  wire[10:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire[3:0] T1161;
  wire[3:0] T1162;
  wire[3:0] T1163;
  wire[10:0] T1164;
  wire[10:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[10:0] T1172;
  wire[10:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[10:0] T1180;
  wire[10:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[10:0] T1188;
  wire[10:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[10:0] T1196;
  wire[10:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[3:0] T1201;
  wire[3:0] T1202;
  wire[3:0] T1203;
  wire[10:0] T1204;
  wire[10:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[10:0] T1212;
  wire[10:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[3:0] T1217;
  wire[3:0] T1218;
  wire[3:0] T1219;
  wire[10:0] T1220;
  wire[10:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[10:0] T1228;
  wire[10:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire[3:0] T1235;
  wire[10:0] T1236;
  wire[10:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[3:0] T1241;
  wire[3:0] T1242;
  wire[3:0] T1243;
  wire[10:0] T1244;
  wire[10:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[3:0] T1249;
  wire[3:0] T1250;
  wire[3:0] T1251;
  wire[10:0] T1252;
  wire[10:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[10:0] T1260;
  wire[10:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[10:0] T1268;
  wire[10:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[10:0] T1276;
  wire[10:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire[3:0] T1281;
  wire[3:0] T1282;
  wire[3:0] T1283;
  wire[10:0] T1284;
  wire[10:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[10:0] T1292;
  wire[10:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[3:0] T1297;
  wire[3:0] T1298;
  wire[3:0] T1299;
  wire[10:0] T1300;
  wire[10:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[10:0] T1308;
  wire[10:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[3:0] T1313;
  wire[3:0] T1314;
  wire[3:0] T1315;
  wire[10:0] T1316;
  wire[10:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[3:0] T1321;
  wire[3:0] T1322;
  wire[3:0] T1323;
  wire[10:0] T1324;
  wire[10:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[3:0] T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[10:0] T1332;
  wire[10:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[10:0] T1340;
  wire[10:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[10:0] T1348;
  wire[10:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[10:0] T1356;
  wire[10:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[3:0] T1361;
  wire[3:0] T1362;
  wire[3:0] T1363;
  wire[10:0] T1364;
  wire[10:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[10:0] T1372;
  wire[10:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire[3:0] T1379;
  wire[10:0] T1380;
  wire[10:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[10:0] T1388;
  wire[10:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[3:0] T1393;
  wire[3:0] T1394;
  wire[3:0] T1395;
  wire[10:0] T1396;
  wire[10:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[5'h16/* 22*/:4'hc/* 12*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[5'h1f/* 31*/:5'h1d/* 29*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[6'h22/* 34*/:6'h20/* 32*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[6'h2d/* 45*/:6'h23/* 35*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h36/* 54*/:6'h34/* 52*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[6'h39/* 57*/:6'h37/* 55*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[7'h44/* 68*/:6'h3a/* 58*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[7'h4d/* 77*/:7'h4b/* 75*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[7'h50/* 80*/:7'h4e/* 78*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[7'h5b/* 91*/:7'h51/* 81*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h35/* 53*/:6'h34/* 52*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h64/* 100*/:7'h62/* 98*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h37/* 55*/:6'h36/* 54*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h67/* 103*/:7'h65/* 101*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h72/* 114*/:7'h68/* 104*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[7'h7e/* 126*/:7'h7c/* 124*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[8'h89/* 137*/:7'h7f/* 127*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[8'h8c/* 140*/:8'h8a/* 138*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[8'h8f/* 143*/:8'h8d/* 141*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[8'h92/* 146*/:8'h90/* 144*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[8'h95/* 149*/:8'h93/* 147*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[8'ha0/* 160*/:8'h96/* 150*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[7'h55/* 85*/:7'h54/* 84*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[7'h57/* 87*/:7'h56/* 86*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[8'ha6/* 166*/:8'ha4/* 164*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[7'h59/* 89*/:7'h58/* 88*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[8'ha9/* 169*/:8'ha7/* 167*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[8'hac/* 172*/:8'haa/* 170*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[8'hb7/* 183*/:8'had/* 173*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[7'h61/* 97*/:7'h60/* 96*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[8'hba/* 186*/:8'hb8/* 184*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[7'h63/* 99*/:7'h62/* 98*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[8'hbd/* 189*/:8'hbb/* 187*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h65/* 101*/:7'h64/* 100*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[8'hc0/* 192*/:8'hbe/* 190*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h67/* 103*/:7'h66/* 102*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'hc3/* 195*/:8'hc1/* 193*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'hce/* 206*/:8'hc4/* 196*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'hd1/* 209*/:8'hcf/* 207*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'hd4/* 212*/:8'hd2/* 210*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h71/* 113*/:7'h70/* 112*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'hd7/* 215*/:8'hd5/* 213*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h73/* 115*/:7'h72/* 114*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'hda/* 218*/:8'hd8/* 216*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'he5/* 229*/:8'hdb/* 219*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'he7/* 231*/:8'he6/* 230*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'he9/* 233*/:8'he8/* 232*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'heb/* 235*/:8'hea/* 234*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h7b/* 123*/:7'h7b/* 123*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hed/* 237*/:8'hec/* 236*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hf8/* 248*/:8'hee/* 238*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'h83/* 131*/:8'h83/* 131*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[9'h10b/* 267*/:9'h101/* 257*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[9'h113/* 275*/:9'h112/* 274*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[9'h11e/* 286*/:9'h114/* 276*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'h92/* 146*/:8'h92/* 146*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'h93/* 147*/:8'h93/* 147*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h126/* 294*/:9'h125/* 293*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h131/* 305*/:9'h127/* 295*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h135/* 309*/:9'h134/* 308*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h137/* 311*/:9'h136/* 310*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h9b/* 155*/:8'h9b/* 155*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h139/* 313*/:9'h138/* 312*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h144/* 324*/:9'h13a/* 314*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'ha2/* 162*/:8'ha2/* 162*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h14a/* 330*/:9'h149/* 329*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'ha3/* 163*/:8'ha3/* 163*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h14c/* 332*/:9'h14b/* 331*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h157/* 343*/:9'h14d/* 333*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h159/* 345*/:9'h158/* 344*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h15b/* 347*/:9'h15a/* 346*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'haa/* 170*/:8'haa/* 170*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h15d/* 349*/:9'h15c/* 348*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'hab/* 171*/:8'hab/* 171*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h15f/* 351*/:9'h15e/* 350*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'haf/* 175*/:8'hac/* 172*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h16a/* 362*/:9'h160/* 352*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h16c/* 364*/:9'h16b/* 363*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h16e/* 366*/:9'h16d/* 365*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h170/* 368*/:9'h16f/* 367*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h172/* 370*/:9'h171/* 369*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h17d/* 381*/:9'h173/* 371*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h17f/* 383*/:9'h17e/* 382*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h181/* 385*/:9'h180/* 384*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h183/* 387*/:9'h182/* 386*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'hbb/* 187*/:8'hbb/* 187*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h185/* 389*/:9'h184/* 388*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h190/* 400*/:9'h186/* 390*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h192/* 402*/:9'h191/* 401*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h194/* 404*/:9'h193/* 403*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h196/* 406*/:9'h195/* 405*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hc3/* 195*/:8'hc3/* 195*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h198/* 408*/:9'h197/* 407*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'hc7/* 199*/:8'hc4/* 196*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h1a3/* 419*/:9'h199/* 409*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h1ae/* 430*/:9'h1a4/* 420*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h1b9/* 441*/:9'h1af/* 431*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h1c4/* 452*/:9'h1ba/* 442*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h1cf/* 463*/:9'h1c5/* 453*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h1da/* 474*/:9'h1d0/* 464*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h1f0/* 496*/:9'h1e6/* 486*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h1fb/* 507*/:9'h1f1/* 497*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h206/* 518*/:9'h1fc/* 508*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h211/* 529*/:10'h207/* 519*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h21c/* 540*/:10'h212/* 530*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h227/* 551*/:10'h21d/* 541*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h232/* 562*/:10'h228/* 552*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h23d/* 573*/:10'h233/* 563*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h248/* 584*/:10'h23e/* 574*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h253/* 595*/:10'h249/* 585*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h10b/* 267*/:9'h108/* 264*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h25e/* 606*/:10'h254/* 596*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h269/* 617*/:10'h25f/* 607*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h113/* 275*/:9'h110/* 272*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h274/* 628*/:10'h26a/* 618*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h117/* 279*/:9'h114/* 276*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h27f/* 639*/:10'h275/* 629*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h28a/* 650*/:10'h280/* 640*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h11f/* 287*/:9'h11c/* 284*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h295/* 661*/:10'h28b/* 651*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h123/* 291*/:9'h120/* 288*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h2a0/* 672*/:10'h296/* 662*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h2ab/* 683*/:10'h2a1/* 673*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h12b/* 299*/:9'h128/* 296*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h2b6/* 694*/:10'h2ac/* 684*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h12f/* 303*/:9'h12c/* 300*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h2c1/* 705*/:10'h2b7/* 695*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h2cc/* 716*/:10'h2c2/* 706*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h2d7/* 727*/:10'h2cd/* 717*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h13b/* 315*/:9'h138/* 312*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h2e2/* 738*/:10'h2d8/* 728*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h13f/* 319*/:9'h13c/* 316*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h2ed/* 749*/:10'h2e3/* 739*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h2f8/* 760*/:10'h2ee/* 750*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h147/* 327*/:9'h144/* 324*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h303/* 771*/:10'h2f9/* 761*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h14b/* 331*/:9'h148/* 328*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h30e/* 782*/:10'h304/* 772*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h14f/* 335*/:9'h14c/* 332*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h319/* 793*/:10'h30f/* 783*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h153/* 339*/:9'h150/* 336*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h324/* 804*/:10'h31a/* 794*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h32f/* 815*/:10'h325/* 805*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h15b/* 347*/:9'h158/* 344*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h33a/* 826*/:10'h330/* 816*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h15f/* 351*/:9'h15c/* 348*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h345/* 837*/:10'h33b/* 827*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h163/* 355*/:9'h160/* 352*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h350/* 848*/:10'h346/* 838*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h164/* 356*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h351/* 849*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_1(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_1 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_2(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[1:0] T281;
  wire[1:0] T282;
  wire[1:0] T283;
  wire[2:0] T284;
  wire[2:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[10:0] T292;
  wire[10:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[1:0] T297;
  wire[1:0] T298;
  wire[1:0] T299;
  wire[2:0] T300;
  wire[2:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[1:0] T305;
  wire[1:0] T306;
  wire[1:0] T307;
  wire[2:0] T308;
  wire[2:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[1:0] T313;
  wire[1:0] T314;
  wire[1:0] T315;
  wire[2:0] T316;
  wire[2:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[1:0] T321;
  wire[1:0] T322;
  wire[1:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[10:0] T332;
  wire[10:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[1:0] T337;
  wire[1:0] T338;
  wire[1:0] T339;
  wire[2:0] T340;
  wire[2:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[1:0] T345;
  wire[1:0] T346;
  wire[1:0] T347;
  wire[2:0] T348;
  wire[2:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[2:0] T356;
  wire[2:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[1:0] T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[2:0] T364;
  wire[2:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[10:0] T372;
  wire[10:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[1:0] T377;
  wire[1:0] T378;
  wire[1:0] T379;
  wire[2:0] T380;
  wire[2:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[1:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[2:0] T388;
  wire[2:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[1:0] T393;
  wire[1:0] T394;
  wire[1:0] T395;
  wire[2:0] T396;
  wire[2:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire[1:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[10:0] T412;
  wire[10:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[1:0] T417;
  wire[1:0] T418;
  wire[1:0] T419;
  wire[2:0] T420;
  wire[2:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T426;
  wire[1:0] T427;
  wire[2:0] T428;
  wire[2:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[2:0] T436;
  wire[2:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[3:0] T449;
  wire[3:0] T450;
  wire[3:0] T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[1:0] T457;
  wire[1:0] T458;
  wire[1:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[1:0] T467;
  wire[2:0] T468;
  wire[2:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire[1:0] T475;
  wire[2:0] T476;
  wire[2:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[1:0] T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[2:0] T484;
  wire[2:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[10:0] T492;
  wire[10:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[2:0] T500;
  wire[2:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[1:0] T505;
  wire[1:0] T506;
  wire[1:0] T507;
  wire[2:0] T508;
  wire[2:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[1:0] T513;
  wire[1:0] T514;
  wire[1:0] T515;
  wire[2:0] T516;
  wire[2:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire[1:0] T523;
  wire[2:0] T524;
  wire[2:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[10:0] T532;
  wire[10:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[1:0] T537;
  wire[1:0] T538;
  wire[1:0] T539;
  wire[2:0] T540;
  wire[2:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[1:0] T545;
  wire[1:0] T546;
  wire[1:0] T547;
  wire[2:0] T548;
  wire[2:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[1:0] T553;
  wire[1:0] T554;
  wire[1:0] T555;
  wire[2:0] T556;
  wire[2:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[1:0] T561;
  wire[1:0] T562;
  wire[1:0] T563;
  wire[2:0] T564;
  wire[2:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[3:0] T569;
  wire[3:0] T570;
  wire[3:0] T571;
  wire[10:0] T572;
  wire[10:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[1:0] T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[2:0] T580;
  wire[2:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[1:0] T585;
  wire[1:0] T586;
  wire[1:0] T587;
  wire[2:0] T588;
  wire[2:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[1:0] T593;
  wire[1:0] T594;
  wire[1:0] T595;
  wire[2:0] T596;
  wire[2:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[3:0] T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[10:0] T612;
  wire[10:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[3:0] T649;
  wire[3:0] T650;
  wire[3:0] T651;
  wire[10:0] T652;
  wire[10:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[3:0] T689;
  wire[3:0] T690;
  wire[3:0] T691;
  wire[10:0] T692;
  wire[10:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[3:0] T729;
  wire[3:0] T730;
  wire[3:0] T731;
  wire[10:0] T732;
  wire[10:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[3:0] T769;
  wire[3:0] T770;
  wire[3:0] T771;
  wire[10:0] T772;
  wire[10:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire[1:0] T780;
  wire[1:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[3:0] T809;
  wire[3:0] T810;
  wire[3:0] T811;
  wire[10:0] T812;
  wire[10:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire[3:0] T849;
  wire[3:0] T850;
  wire[3:0] T851;
  wire[10:0] T852;
  wire[10:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[3:0] T890;
  wire[3:0] T891;
  wire[10:0] T892;
  wire[10:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[3:0] T929;
  wire[3:0] T930;
  wire[3:0] T931;
  wire[10:0] T932;
  wire[10:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire[1:0] T940;
  wire[1:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[3:0] T969;
  wire[3:0] T970;
  wire[3:0] T971;
  wire[10:0] T972;
  wire[10:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire[3:0] T1009;
  wire[3:0] T1010;
  wire[3:0] T1011;
  wire[10:0] T1012;
  wire[10:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire[3:0] T1049;
  wire[3:0] T1050;
  wire[3:0] T1051;
  wire[10:0] T1052;
  wire[10:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire[3:0] T1081;
  wire[3:0] T1082;
  wire[3:0] T1083;
  wire[10:0] T1084;
  wire[10:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[10:0] T1092;
  wire[10:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[10:0] T1100;
  wire[10:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[10:0] T1108;
  wire[10:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[10:0] T1116;
  wire[10:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[10:0] T1124;
  wire[10:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[10:0] T1132;
  wire[10:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[10:0] T1140;
  wire[10:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[10:0] T1148;
  wire[10:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[10:0] T1156;
  wire[10:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire[3:0] T1161;
  wire[3:0] T1162;
  wire[3:0] T1163;
  wire[10:0] T1164;
  wire[10:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[10:0] T1172;
  wire[10:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[10:0] T1180;
  wire[10:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[10:0] T1188;
  wire[10:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[10:0] T1196;
  wire[10:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[3:0] T1201;
  wire[3:0] T1202;
  wire[3:0] T1203;
  wire[10:0] T1204;
  wire[10:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[10:0] T1212;
  wire[10:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[3:0] T1217;
  wire[3:0] T1218;
  wire[3:0] T1219;
  wire[10:0] T1220;
  wire[10:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[10:0] T1228;
  wire[10:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire[3:0] T1235;
  wire[10:0] T1236;
  wire[10:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[3:0] T1241;
  wire[3:0] T1242;
  wire[3:0] T1243;
  wire[10:0] T1244;
  wire[10:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[3:0] T1249;
  wire[3:0] T1250;
  wire[3:0] T1251;
  wire[10:0] T1252;
  wire[10:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[10:0] T1260;
  wire[10:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[10:0] T1268;
  wire[10:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[10:0] T1276;
  wire[10:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire[3:0] T1281;
  wire[3:0] T1282;
  wire[3:0] T1283;
  wire[10:0] T1284;
  wire[10:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[10:0] T1292;
  wire[10:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[3:0] T1297;
  wire[3:0] T1298;
  wire[3:0] T1299;
  wire[10:0] T1300;
  wire[10:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[10:0] T1308;
  wire[10:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[3:0] T1313;
  wire[3:0] T1314;
  wire[3:0] T1315;
  wire[10:0] T1316;
  wire[10:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[3:0] T1321;
  wire[3:0] T1322;
  wire[3:0] T1323;
  wire[10:0] T1324;
  wire[10:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[3:0] T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[10:0] T1332;
  wire[10:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[10:0] T1340;
  wire[10:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[10:0] T1348;
  wire[10:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[10:0] T1356;
  wire[10:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[3:0] T1361;
  wire[3:0] T1362;
  wire[3:0] T1363;
  wire[10:0] T1364;
  wire[10:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[10:0] T1372;
  wire[10:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire[3:0] T1379;
  wire[10:0] T1380;
  wire[10:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[10:0] T1388;
  wire[10:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[3:0] T1393;
  wire[3:0] T1394;
  wire[3:0] T1395;
  wire[10:0] T1396;
  wire[10:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[3'h5/* 5*/:2'h2/* 2*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[4'hd/* 13*/:2'h3/* 3*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[5'h10/* 16*/:4'he/* 14*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[5'h13/* 19*/:5'h11/* 17*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h11/* 17*/:4'he/* 14*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[6'h24/* 36*/:5'h1a/* 26*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[6'h27/* 39*/:6'h25/* 37*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h15/* 21*/:5'h14/* 20*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[6'h2a/* 42*/:6'h28/* 40*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h1d/* 29*/:5'h1a/* 26*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h3b/* 59*/:6'h31/* 49*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h3e/* 62*/:6'h3c/* 60*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[7'h41/* 65*/:6'h3f/* 63*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[6'h29/* 41*/:6'h26/* 38*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[7'h52/* 82*/:7'h48/* 72*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[7'h55/* 85*/:7'h53/* 83*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[7'h58/* 88*/:7'h56/* 86*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h35/* 53*/:6'h32/* 50*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h69/* 105*/:7'h5f/* 95*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h37/* 55*/:6'h36/* 54*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h6c/* 108*/:7'h6a/* 106*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h39/* 57*/:6'h38/* 56*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h41/* 65*/:6'h3e/* 62*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[8'h80/* 128*/:7'h76/* 118*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[8'h83/* 131*/:8'h81/* 129*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[8'h86/* 134*/:8'h84/* 132*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[8'h8c/* 140*/:8'h8a/* 138*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h4d/* 77*/:7'h4a/* 74*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[8'h97/* 151*/:8'h8d/* 141*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[8'h9a/* 154*/:8'h98/* 152*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[7'h51/* 81*/:7'h50/* 80*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[8'h9d/* 157*/:8'h9b/* 155*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[7'h53/* 83*/:7'h52/* 82*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[8'ha0/* 160*/:8'h9e/* 158*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[7'h55/* 85*/:7'h54/* 84*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[7'h59/* 89*/:7'h56/* 86*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[8'hae/* 174*/:8'ha4/* 164*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[8'hb1/* 177*/:8'haf/* 175*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[8'hb4/* 180*/:8'hb2/* 178*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[8'hb7/* 183*/:8'hb5/* 181*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[7'h61/* 97*/:7'h60/* 96*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[8'hba/* 186*/:8'hb8/* 184*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[7'h65/* 101*/:7'h62/* 98*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[8'hc5/* 197*/:8'hbb/* 187*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h67/* 103*/:7'h66/* 102*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[8'hc8/* 200*/:8'hc6/* 198*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h69/* 105*/:7'h68/* 104*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'hcb/* 203*/:8'hc9/* 201*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'hce/* 206*/:8'hcc/* 204*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'hd1/* 209*/:8'hcf/* 207*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h71/* 113*/:7'h6e/* 110*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'hdc/* 220*/:8'hd2/* 210*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h73/* 115*/:7'h72/* 114*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'hdf/* 223*/:8'hdd/* 221*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h75/* 117*/:7'h74/* 116*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'he2/* 226*/:8'he0/* 224*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h77/* 119*/:7'h76/* 118*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'he5/* 229*/:8'he3/* 227*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'he7/* 231*/:8'he6/* 230*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h7c/* 124*/:7'h79/* 121*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'hf2/* 242*/:8'he8/* 232*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h7d/* 125*/:7'h7d/* 125*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'hf4/* 244*/:8'hf3/* 243*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hf6/* 246*/:8'hf5/* 245*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'h84/* 132*/:8'h81/* 129*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[9'h105/* 261*/:8'hfb/* 251*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'h85/* 133*/:8'h85/* 133*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[9'h107/* 263*/:9'h106/* 262*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[9'h109/* 265*/:9'h108/* 264*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'h8c/* 140*/:8'h89/* 137*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[9'h118/* 280*/:9'h10e/* 270*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'h8d/* 141*/:8'h8d/* 141*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[9'h11a/* 282*/:9'h119/* 281*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'h94/* 148*/:8'h91/* 145*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h12b/* 299*/:9'h121/* 289*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'h95/* 149*/:8'h95/* 149*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h12d/* 301*/:9'h12c/* 300*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'h96/* 150*/:8'h96/* 150*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h9c/* 156*/:8'h99/* 153*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h13e/* 318*/:9'h134/* 308*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h9d/* 157*/:8'h9d/* 157*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h140/* 320*/:9'h13f/* 319*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'ha4/* 164*/:8'ha1/* 161*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h151/* 337*/:9'h147/* 327*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'ha5/* 165*/:8'ha5/* 165*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'ha6/* 166*/:8'ha6/* 166*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h155/* 341*/:9'h154/* 340*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h157/* 343*/:9'h156/* 342*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h159/* 345*/:9'h158/* 344*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'hac/* 172*/:8'ha9/* 169*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h164/* 356*/:9'h15a/* 346*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'had/* 173*/:8'had/* 173*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h166/* 358*/:9'h165/* 357*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h168/* 360*/:9'h167/* 359*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h16a/* 362*/:9'h169/* 361*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h16c/* 364*/:9'h16b/* 363*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'hb4/* 180*/:8'hb1/* 177*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h177/* 375*/:9'h16d/* 365*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h179/* 377*/:9'h178/* 376*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h17b/* 379*/:9'h17a/* 378*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'hb7/* 183*/:8'hb7/* 183*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h17d/* 381*/:9'h17c/* 380*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h17f/* 383*/:9'h17e/* 382*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'hbc/* 188*/:8'hb9/* 185*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h18a/* 394*/:9'h180/* 384*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h18c/* 396*/:9'h18b/* 395*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'hbe/* 190*/:8'hbe/* 190*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h18e/* 398*/:9'h18d/* 397*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'hbf/* 191*/:8'hbf/* 191*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h190/* 400*/:9'h18f/* 399*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h192/* 402*/:9'h191/* 401*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'hc4/* 196*/:8'hc1/* 193*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h19d/* 413*/:9'h193/* 403*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'hc5/* 197*/:8'hc5/* 197*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h19f/* 415*/:9'h19e/* 414*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hc6/* 198*/:8'hc6/* 198*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h1a1/* 417*/:9'h1a0/* 416*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h1ae/* 430*/:9'h1a4/* 420*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h1b9/* 441*/:9'h1af/* 431*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h1c4/* 452*/:9'h1ba/* 442*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h1cf/* 463*/:9'h1c5/* 453*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h1da/* 474*/:9'h1d0/* 464*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h1f0/* 496*/:9'h1e6/* 486*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h1fb/* 507*/:9'h1f1/* 497*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h206/* 518*/:9'h1fc/* 508*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h211/* 529*/:10'h207/* 519*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h21c/* 540*/:10'h212/* 530*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h227/* 551*/:10'h21d/* 541*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h232/* 562*/:10'h228/* 552*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h23d/* 573*/:10'h233/* 563*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h248/* 584*/:10'h23e/* 574*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h253/* 595*/:10'h249/* 585*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h10b/* 267*/:9'h108/* 264*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h25e/* 606*/:10'h254/* 596*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h269/* 617*/:10'h25f/* 607*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h113/* 275*/:9'h110/* 272*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h274/* 628*/:10'h26a/* 618*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h117/* 279*/:9'h114/* 276*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h27f/* 639*/:10'h275/* 629*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h28a/* 650*/:10'h280/* 640*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h11f/* 287*/:9'h11c/* 284*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h295/* 661*/:10'h28b/* 651*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h123/* 291*/:9'h120/* 288*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h2a0/* 672*/:10'h296/* 662*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h2ab/* 683*/:10'h2a1/* 673*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h12b/* 299*/:9'h128/* 296*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h2b6/* 694*/:10'h2ac/* 684*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h12f/* 303*/:9'h12c/* 300*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h2c1/* 705*/:10'h2b7/* 695*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h2cc/* 716*/:10'h2c2/* 706*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h2d7/* 727*/:10'h2cd/* 717*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h13b/* 315*/:9'h138/* 312*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h2e2/* 738*/:10'h2d8/* 728*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h13f/* 319*/:9'h13c/* 316*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h2ed/* 749*/:10'h2e3/* 739*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h2f8/* 760*/:10'h2ee/* 750*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h147/* 327*/:9'h144/* 324*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h303/* 771*/:10'h2f9/* 761*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h14b/* 331*/:9'h148/* 328*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h30e/* 782*/:10'h304/* 772*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h14f/* 335*/:9'h14c/* 332*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h319/* 793*/:10'h30f/* 783*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h153/* 339*/:9'h150/* 336*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h324/* 804*/:10'h31a/* 794*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h32f/* 815*/:10'h325/* 805*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h15b/* 347*/:9'h158/* 344*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h33a/* 826*/:10'h330/* 816*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h15f/* 351*/:9'h15c/* 348*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h345/* 837*/:10'h33b/* 827*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h163/* 355*/:9'h160/* 352*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h350/* 848*/:10'h346/* 838*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h164/* 356*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h351/* 849*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_2(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_2 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_3(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[1:0] T281;
  wire[1:0] T282;
  wire[1:0] T283;
  wire[2:0] T284;
  wire[2:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[1:0] T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[10:0] T300;
  wire[10:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[1:0] T305;
  wire[1:0] T306;
  wire[1:0] T307;
  wire[2:0] T308;
  wire[2:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[1:0] T313;
  wire[1:0] T314;
  wire[1:0] T315;
  wire[2:0] T316;
  wire[2:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[1:0] T321;
  wire[1:0] T322;
  wire[1:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[1:0] T330;
  wire[1:0] T331;
  wire[2:0] T332;
  wire[2:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[10:0] T340;
  wire[10:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[1:0] T345;
  wire[1:0] T346;
  wire[1:0] T347;
  wire[2:0] T348;
  wire[2:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[2:0] T356;
  wire[2:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[1:0] T361;
  wire[1:0] T362;
  wire[1:0] T363;
  wire[2:0] T364;
  wire[2:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[1:0] T369;
  wire[1:0] T370;
  wire[1:0] T371;
  wire[2:0] T372;
  wire[2:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[10:0] T380;
  wire[10:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[1:0] T385;
  wire[1:0] T386;
  wire[1:0] T387;
  wire[2:0] T388;
  wire[2:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[1:0] T393;
  wire[1:0] T394;
  wire[1:0] T395;
  wire[2:0] T396;
  wire[2:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire[1:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[1:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire[2:0] T412;
  wire[2:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[10:0] T420;
  wire[10:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T426;
  wire[1:0] T427;
  wire[2:0] T428;
  wire[2:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[2:0] T436;
  wire[2:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[1:0] T449;
  wire[1:0] T450;
  wire[1:0] T451;
  wire[2:0] T452;
  wire[2:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[10:0] T460;
  wire[10:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[1:0] T467;
  wire[2:0] T468;
  wire[2:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire[1:0] T475;
  wire[2:0] T476;
  wire[2:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[1:0] T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[2:0] T484;
  wire[2:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[1:0] T489;
  wire[1:0] T490;
  wire[1:0] T491;
  wire[2:0] T492;
  wire[2:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[10:0] T500;
  wire[10:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[1:0] T505;
  wire[1:0] T506;
  wire[1:0] T507;
  wire[2:0] T508;
  wire[2:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[1:0] T513;
  wire[1:0] T514;
  wire[1:0] T515;
  wire[2:0] T516;
  wire[2:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[1:0] T521;
  wire[1:0] T522;
  wire[1:0] T523;
  wire[2:0] T524;
  wire[2:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[1:0] T529;
  wire[1:0] T530;
  wire[1:0] T531;
  wire[2:0] T532;
  wire[2:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[10:0] T540;
  wire[10:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[1:0] T545;
  wire[1:0] T546;
  wire[1:0] T547;
  wire[2:0] T548;
  wire[2:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[1:0] T553;
  wire[1:0] T554;
  wire[1:0] T555;
  wire[2:0] T556;
  wire[2:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[1:0] T561;
  wire[1:0] T562;
  wire[1:0] T563;
  wire[2:0] T564;
  wire[2:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[1:0] T569;
  wire[1:0] T570;
  wire[1:0] T571;
  wire[2:0] T572;
  wire[2:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[10:0] T580;
  wire[10:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[1:0] T585;
  wire[1:0] T586;
  wire[1:0] T587;
  wire[2:0] T588;
  wire[2:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[1:0] T593;
  wire[1:0] T594;
  wire[1:0] T595;
  wire[2:0] T596;
  wire[2:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[3:0] T617;
  wire[3:0] T618;
  wire[3:0] T619;
  wire[10:0] T620;
  wire[10:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[3:0] T657;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[10:0] T660;
  wire[10:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[10:0] T700;
  wire[10:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[3:0] T737;
  wire[3:0] T738;
  wire[3:0] T739;
  wire[10:0] T740;
  wire[10:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[10:0] T780;
  wire[10:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[3:0] T817;
  wire[3:0] T818;
  wire[3:0] T819;
  wire[10:0] T820;
  wire[10:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[10:0] T860;
  wire[10:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[10:0] T900;
  wire[10:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[10:0] T940;
  wire[10:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[10:0] T980;
  wire[10:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire[3:0] T1017;
  wire[3:0] T1018;
  wire[3:0] T1019;
  wire[10:0] T1020;
  wire[10:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire[3:0] T1057;
  wire[3:0] T1058;
  wire[3:0] T1059;
  wire[10:0] T1060;
  wire[10:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire[3:0] T1081;
  wire[3:0] T1082;
  wire[3:0] T1083;
  wire[10:0] T1084;
  wire[10:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[10:0] T1092;
  wire[10:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[10:0] T1100;
  wire[10:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[10:0] T1108;
  wire[10:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[10:0] T1116;
  wire[10:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[10:0] T1124;
  wire[10:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[10:0] T1132;
  wire[10:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[10:0] T1140;
  wire[10:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[10:0] T1148;
  wire[10:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[10:0] T1156;
  wire[10:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire[3:0] T1161;
  wire[3:0] T1162;
  wire[3:0] T1163;
  wire[10:0] T1164;
  wire[10:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[10:0] T1172;
  wire[10:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[10:0] T1180;
  wire[10:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[10:0] T1188;
  wire[10:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[10:0] T1196;
  wire[10:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[3:0] T1201;
  wire[3:0] T1202;
  wire[3:0] T1203;
  wire[10:0] T1204;
  wire[10:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[10:0] T1212;
  wire[10:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[3:0] T1217;
  wire[3:0] T1218;
  wire[3:0] T1219;
  wire[10:0] T1220;
  wire[10:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[10:0] T1228;
  wire[10:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire[3:0] T1235;
  wire[10:0] T1236;
  wire[10:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[3:0] T1241;
  wire[3:0] T1242;
  wire[3:0] T1243;
  wire[10:0] T1244;
  wire[10:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[3:0] T1249;
  wire[3:0] T1250;
  wire[3:0] T1251;
  wire[10:0] T1252;
  wire[10:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[10:0] T1260;
  wire[10:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[10:0] T1268;
  wire[10:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[10:0] T1276;
  wire[10:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire[3:0] T1281;
  wire[3:0] T1282;
  wire[3:0] T1283;
  wire[10:0] T1284;
  wire[10:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[10:0] T1292;
  wire[10:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[3:0] T1297;
  wire[3:0] T1298;
  wire[3:0] T1299;
  wire[10:0] T1300;
  wire[10:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[10:0] T1308;
  wire[10:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[3:0] T1313;
  wire[3:0] T1314;
  wire[3:0] T1315;
  wire[10:0] T1316;
  wire[10:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[3:0] T1321;
  wire[3:0] T1322;
  wire[3:0] T1323;
  wire[10:0] T1324;
  wire[10:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[3:0] T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[10:0] T1332;
  wire[10:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[10:0] T1340;
  wire[10:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[10:0] T1348;
  wire[10:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[10:0] T1356;
  wire[10:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[3:0] T1361;
  wire[3:0] T1362;
  wire[3:0] T1363;
  wire[10:0] T1364;
  wire[10:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[10:0] T1372;
  wire[10:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire[3:0] T1379;
  wire[10:0] T1380;
  wire[10:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[10:0] T1388;
  wire[10:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[3:0] T1393;
  wire[3:0] T1394;
  wire[3:0] T1395;
  wire[10:0] T1396;
  wire[10:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[5'h10/* 16*/:3'h6/* 6*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[5'h13/* 19*/:5'h11/* 17*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[5'h16/* 22*/:5'h14/* 20*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[5'h19/* 25*/:5'h17/* 23*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[5'h1c/* 28*/:5'h1a/* 26*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[6'h27/* 39*/:5'h1d/* 29*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h15/* 21*/:5'h14/* 20*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[6'h2a/* 42*/:6'h28/* 40*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h17/* 23*/:5'h16/* 22*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[6'h2d/* 45*/:6'h2b/* 43*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h19/* 25*/:5'h18/* 24*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[6'h30/* 48*/:6'h2e/* 46*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h33/* 51*/:6'h31/* 49*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h3e/* 62*/:6'h34/* 52*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[7'h41/* 65*/:6'h3f/* 63*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[7'h44/* 68*/:7'h42/* 66*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[7'h47/* 71*/:7'h45/* 69*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[7'h4a/* 74*/:7'h48/* 72*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[7'h55/* 85*/:7'h4b/* 75*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[7'h58/* 88*/:7'h56/* 86*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[7'h5b/* 91*/:7'h59/* 89*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[7'h5e/* 94*/:7'h5c/* 92*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h33/* 51*/:6'h32/* 50*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[7'h61/* 97*/:7'h5f/* 95*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[7'h6c/* 108*/:7'h62/* 98*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h39/* 57*/:6'h38/* 56*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[8'h83/* 131*/:7'h79/* 121*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[8'h86/* 134*/:8'h84/* 132*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[8'h89/* 137*/:8'h87/* 135*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[8'h8c/* 140*/:8'h8a/* 138*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[8'h8f/* 143*/:8'h8d/* 141*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[8'h9a/* 154*/:8'h90/* 144*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[7'h51/* 81*/:7'h50/* 80*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[8'h9d/* 157*/:8'h9b/* 155*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[7'h53/* 83*/:7'h52/* 82*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[8'ha0/* 160*/:8'h9e/* 158*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[7'h55/* 85*/:7'h54/* 84*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[7'h57/* 87*/:7'h56/* 86*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[8'ha6/* 166*/:8'ha4/* 164*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[8'hb1/* 177*/:8'ha7/* 167*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[8'hb4/* 180*/:8'hb2/* 178*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[8'hb7/* 183*/:8'hb5/* 181*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[7'h61/* 97*/:7'h60/* 96*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[8'hba/* 186*/:8'hb8/* 184*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[7'h63/* 99*/:7'h62/* 98*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[8'hbd/* 189*/:8'hbb/* 187*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[8'hc8/* 200*/:8'hbe/* 190*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h69/* 105*/:7'h68/* 104*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[8'hcb/* 203*/:8'hc9/* 201*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[8'hce/* 206*/:8'hcc/* 204*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[8'hd1/* 209*/:8'hcf/* 207*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[8'hd4/* 212*/:8'hd2/* 210*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[8'hdf/* 223*/:8'hd5/* 213*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h75/* 117*/:7'h74/* 116*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[8'he2/* 226*/:8'he0/* 224*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h77/* 119*/:7'h76/* 118*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'he5/* 229*/:8'he3/* 227*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'he7/* 231*/:8'he6/* 230*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'he9/* 233*/:8'he8/* 232*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h7d/* 125*/:7'h7a/* 122*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'hf4/* 244*/:8'hea/* 234*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h7e/* 126*/:7'h7e/* 126*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'hf6/* 246*/:8'hf5/* 245*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'hf8/* 248*/:8'hf7/* 247*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'hfa/* 250*/:8'hf9/* 249*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'hfc/* 252*/:8'hfb/* 251*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[9'h107/* 263*/:8'hfd/* 253*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[9'h109/* 265*/:9'h108/* 264*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[9'h11a/* 282*/:9'h110/* 272*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'h8e/* 142*/:8'h8e/* 142*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[9'h11e/* 286*/:9'h11d/* 285*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'h95/* 149*/:8'h92/* 146*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h12d/* 301*/:9'h123/* 291*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'h96/* 150*/:8'h96/* 150*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h135/* 309*/:9'h134/* 308*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h9d/* 157*/:8'h9a/* 154*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h140/* 320*/:9'h136/* 310*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h9e/* 158*/:8'h9e/* 158*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'ha0/* 160*/:8'ha0/* 160*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'ha1/* 161*/:8'ha1/* 161*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'ha5/* 165*/:8'ha2/* 162*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h153/* 339*/:9'h149/* 329*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'ha6/* 166*/:8'ha6/* 166*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h155/* 341*/:9'h154/* 340*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h157/* 343*/:9'h156/* 342*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h159/* 345*/:9'h158/* 344*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h15b/* 347*/:9'h15a/* 346*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'had/* 173*/:8'haa/* 170*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h166/* 358*/:9'h15c/* 348*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h168/* 360*/:9'h167/* 359*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h16a/* 362*/:9'h169/* 361*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h16c/* 364*/:9'h16b/* 363*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h16e/* 366*/:9'h16d/* 365*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'hb5/* 181*/:8'hb2/* 178*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h179/* 377*/:9'h16f/* 367*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h17b/* 379*/:9'h17a/* 378*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'hb7/* 183*/:8'hb7/* 183*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h17d/* 381*/:9'h17c/* 380*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h17f/* 383*/:9'h17e/* 382*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h181/* 385*/:9'h180/* 384*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'hbd/* 189*/:8'hba/* 186*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h18c/* 396*/:9'h182/* 386*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'hbe/* 190*/:8'hbe/* 190*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h18e/* 398*/:9'h18d/* 397*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'hbf/* 191*/:8'hbf/* 191*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h190/* 400*/:9'h18f/* 399*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h192/* 402*/:9'h191/* 401*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h194/* 404*/:9'h193/* 403*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'hc5/* 197*/:8'hc2/* 194*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h19f/* 415*/:9'h195/* 405*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hc6/* 198*/:8'hc6/* 198*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h1a1/* 417*/:9'h1a0/* 416*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h1ae/* 430*/:9'h1a4/* 420*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h1b9/* 441*/:9'h1af/* 431*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h1c4/* 452*/:9'h1ba/* 442*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h1cf/* 463*/:9'h1c5/* 453*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h1da/* 474*/:9'h1d0/* 464*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h1f0/* 496*/:9'h1e6/* 486*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h1fb/* 507*/:9'h1f1/* 497*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h206/* 518*/:9'h1fc/* 508*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h211/* 529*/:10'h207/* 519*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h21c/* 540*/:10'h212/* 530*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h227/* 551*/:10'h21d/* 541*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h232/* 562*/:10'h228/* 552*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h23d/* 573*/:10'h233/* 563*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h248/* 584*/:10'h23e/* 574*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h253/* 595*/:10'h249/* 585*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h10b/* 267*/:9'h108/* 264*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h25e/* 606*/:10'h254/* 596*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h269/* 617*/:10'h25f/* 607*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h113/* 275*/:9'h110/* 272*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h274/* 628*/:10'h26a/* 618*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h117/* 279*/:9'h114/* 276*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h27f/* 639*/:10'h275/* 629*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h28a/* 650*/:10'h280/* 640*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h11f/* 287*/:9'h11c/* 284*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h295/* 661*/:10'h28b/* 651*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h123/* 291*/:9'h120/* 288*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h2a0/* 672*/:10'h296/* 662*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h2ab/* 683*/:10'h2a1/* 673*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h12b/* 299*/:9'h128/* 296*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h2b6/* 694*/:10'h2ac/* 684*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h12f/* 303*/:9'h12c/* 300*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h2c1/* 705*/:10'h2b7/* 695*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h2cc/* 716*/:10'h2c2/* 706*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h2d7/* 727*/:10'h2cd/* 717*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h13b/* 315*/:9'h138/* 312*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h2e2/* 738*/:10'h2d8/* 728*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h13f/* 319*/:9'h13c/* 316*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h2ed/* 749*/:10'h2e3/* 739*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h2f8/* 760*/:10'h2ee/* 750*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h147/* 327*/:9'h144/* 324*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h303/* 771*/:10'h2f9/* 761*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h14b/* 331*/:9'h148/* 328*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h30e/* 782*/:10'h304/* 772*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h14f/* 335*/:9'h14c/* 332*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h319/* 793*/:10'h30f/* 783*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h153/* 339*/:9'h150/* 336*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h324/* 804*/:10'h31a/* 794*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h32f/* 815*/:10'h325/* 805*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h15b/* 347*/:9'h158/* 344*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h33a/* 826*/:10'h330/* 816*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h15f/* 351*/:9'h15c/* 348*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h345/* 837*/:10'h33b/* 827*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h163/* 355*/:9'h160/* 352*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h350/* 848*/:10'h346/* 838*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h164/* 356*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h351/* 849*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_3(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_3 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_4(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [759:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[199:0] io_chanxy_out);

  wire[199:0] T0;
  wire[199:0] T1;
  wire[198:0] T2;
  wire[198:0] T3;
  wire[197:0] T4;
  wire[197:0] T5;
  wire[196:0] T6;
  wire[196:0] T7;
  wire[195:0] T8;
  wire[195:0] T9;
  wire[194:0] T10;
  wire[194:0] T11;
  wire[193:0] T12;
  wire[193:0] T13;
  wire[192:0] T14;
  wire[192:0] T15;
  wire[191:0] T16;
  wire[191:0] T17;
  wire[190:0] T18;
  wire[190:0] T19;
  wire[189:0] T20;
  wire[189:0] T21;
  wire[188:0] T22;
  wire[188:0] T23;
  wire[187:0] T24;
  wire[187:0] T25;
  wire[186:0] T26;
  wire[186:0] T27;
  wire[185:0] T28;
  wire[185:0] T29;
  wire[184:0] T30;
  wire[184:0] T31;
  wire[183:0] T32;
  wire[183:0] T33;
  wire[182:0] T34;
  wire[182:0] T35;
  wire[181:0] T36;
  wire[181:0] T37;
  wire[180:0] T38;
  wire[180:0] T39;
  wire[179:0] T40;
  wire[179:0] T41;
  wire[178:0] T42;
  wire[178:0] T43;
  wire[177:0] T44;
  wire[177:0] T45;
  wire[176:0] T46;
  wire[176:0] T47;
  wire[175:0] T48;
  wire[175:0] T49;
  wire[174:0] T50;
  wire[174:0] T51;
  wire[173:0] T52;
  wire[173:0] T53;
  wire[172:0] T54;
  wire[172:0] T55;
  wire[171:0] T56;
  wire[171:0] T57;
  wire[170:0] T58;
  wire[170:0] T59;
  wire[169:0] T60;
  wire[169:0] T61;
  wire[168:0] T62;
  wire[168:0] T63;
  wire[167:0] T64;
  wire[167:0] T65;
  wire[166:0] T66;
  wire[166:0] T67;
  wire[165:0] T68;
  wire[165:0] T69;
  wire[164:0] T70;
  wire[164:0] T71;
  wire[163:0] T72;
  wire[163:0] T73;
  wire[162:0] T74;
  wire[162:0] T75;
  wire[161:0] T76;
  wire[161:0] T77;
  wire[160:0] T78;
  wire[160:0] T79;
  wire[159:0] T80;
  wire[159:0] T81;
  wire[158:0] T82;
  wire[158:0] T83;
  wire[157:0] T84;
  wire[157:0] T85;
  wire[156:0] T86;
  wire[156:0] T87;
  wire[155:0] T88;
  wire[155:0] T89;
  wire[154:0] T90;
  wire[154:0] T91;
  wire[153:0] T92;
  wire[153:0] T93;
  wire[152:0] T94;
  wire[152:0] T95;
  wire[151:0] T96;
  wire[151:0] T97;
  wire[150:0] T98;
  wire[150:0] T99;
  wire[149:0] T100;
  wire[149:0] T101;
  wire[148:0] T102;
  wire[148:0] T103;
  wire[147:0] T104;
  wire[147:0] T105;
  wire[146:0] T106;
  wire[146:0] T107;
  wire[145:0] T108;
  wire[145:0] T109;
  wire[144:0] T110;
  wire[144:0] T111;
  wire[143:0] T112;
  wire[143:0] T113;
  wire[142:0] T114;
  wire[142:0] T115;
  wire[141:0] T116;
  wire[141:0] T117;
  wire[140:0] T118;
  wire[140:0] T119;
  wire[139:0] T120;
  wire[139:0] T121;
  wire[138:0] T122;
  wire[138:0] T123;
  wire[137:0] T124;
  wire[137:0] T125;
  wire[136:0] T126;
  wire[136:0] T127;
  wire[135:0] T128;
  wire[135:0] T129;
  wire[134:0] T130;
  wire[134:0] T131;
  wire[133:0] T132;
  wire[133:0] T133;
  wire[132:0] T134;
  wire[132:0] T135;
  wire[131:0] T136;
  wire[131:0] T137;
  wire[130:0] T138;
  wire[130:0] T139;
  wire[129:0] T140;
  wire[129:0] T141;
  wire[128:0] T142;
  wire[128:0] T143;
  wire[127:0] T144;
  wire[127:0] T145;
  wire[126:0] T146;
  wire[126:0] T147;
  wire[125:0] T148;
  wire[125:0] T149;
  wire[124:0] T150;
  wire[124:0] T151;
  wire[123:0] T152;
  wire[123:0] T153;
  wire[122:0] T154;
  wire[122:0] T155;
  wire[121:0] T156;
  wire[121:0] T157;
  wire[120:0] T158;
  wire[120:0] T159;
  wire[119:0] T160;
  wire[119:0] T161;
  wire[118:0] T162;
  wire[118:0] T163;
  wire[117:0] T164;
  wire[117:0] T165;
  wire[116:0] T166;
  wire[116:0] T167;
  wire[115:0] T168;
  wire[115:0] T169;
  wire[114:0] T170;
  wire[114:0] T171;
  wire[113:0] T172;
  wire[113:0] T173;
  wire[112:0] T174;
  wire[112:0] T175;
  wire[111:0] T176;
  wire[111:0] T177;
  wire[110:0] T178;
  wire[110:0] T179;
  wire[109:0] T180;
  wire[109:0] T181;
  wire[108:0] T182;
  wire[108:0] T183;
  wire[107:0] T184;
  wire[107:0] T185;
  wire[106:0] T186;
  wire[106:0] T187;
  wire[105:0] T188;
  wire[105:0] T189;
  wire[104:0] T190;
  wire[104:0] T191;
  wire[103:0] T192;
  wire[103:0] T193;
  wire[102:0] T194;
  wire[102:0] T195;
  wire[101:0] T196;
  wire[101:0] T197;
  wire[100:0] T198;
  wire[100:0] T199;
  wire[99:0] T200;
  wire[99:0] T201;
  wire[98:0] T202;
  wire[98:0] T203;
  wire[97:0] T204;
  wire[97:0] T205;
  wire[96:0] T206;
  wire[96:0] T207;
  wire[95:0] T208;
  wire[95:0] T209;
  wire[94:0] T210;
  wire[94:0] T211;
  wire[93:0] T212;
  wire[93:0] T213;
  wire[92:0] T214;
  wire[92:0] T215;
  wire[91:0] T216;
  wire[91:0] T217;
  wire[90:0] T218;
  wire[90:0] T219;
  wire[89:0] T220;
  wire[89:0] T221;
  wire[88:0] T222;
  wire[88:0] T223;
  wire[87:0] T224;
  wire[87:0] T225;
  wire[86:0] T226;
  wire[86:0] T227;
  wire[85:0] T228;
  wire[85:0] T229;
  wire[84:0] T230;
  wire[84:0] T231;
  wire[83:0] T232;
  wire[83:0] T233;
  wire[82:0] T234;
  wire[82:0] T235;
  wire[81:0] T236;
  wire[81:0] T237;
  wire[80:0] T238;
  wire[80:0] T239;
  wire[79:0] T240;
  wire[79:0] T241;
  wire[78:0] T242;
  wire[78:0] T243;
  wire[77:0] T244;
  wire[77:0] T245;
  wire[76:0] T246;
  wire[76:0] T247;
  wire[75:0] T248;
  wire[75:0] T249;
  wire[74:0] T250;
  wire[74:0] T251;
  wire[73:0] T252;
  wire[73:0] T253;
  wire[72:0] T254;
  wire[72:0] T255;
  wire[71:0] T256;
  wire[71:0] T257;
  wire[70:0] T258;
  wire[70:0] T259;
  wire[69:0] T260;
  wire[69:0] T261;
  wire[68:0] T262;
  wire[68:0] T263;
  wire[67:0] T264;
  wire[67:0] T265;
  wire[66:0] T266;
  wire[66:0] T267;
  wire[65:0] T268;
  wire[65:0] T269;
  wire[64:0] T270;
  wire[64:0] T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[62:0] T274;
  wire[62:0] T275;
  wire[61:0] T276;
  wire[61:0] T277;
  wire[60:0] T278;
  wire[60:0] T279;
  wire[59:0] T280;
  wire[59:0] T281;
  wire[58:0] T282;
  wire[58:0] T283;
  wire[57:0] T284;
  wire[57:0] T285;
  wire[56:0] T286;
  wire[56:0] T287;
  wire[55:0] T288;
  wire[55:0] T289;
  wire[54:0] T290;
  wire[54:0] T291;
  wire[53:0] T292;
  wire[53:0] T293;
  wire[52:0] T294;
  wire[52:0] T295;
  wire[51:0] T296;
  wire[51:0] T297;
  wire[50:0] T298;
  wire[50:0] T299;
  wire[49:0] T300;
  wire[49:0] T301;
  wire[48:0] T302;
  wire[48:0] T303;
  wire[47:0] T304;
  wire[47:0] T305;
  wire[46:0] T306;
  wire[46:0] T307;
  wire[45:0] T308;
  wire[45:0] T309;
  wire[44:0] T310;
  wire[44:0] T311;
  wire[43:0] T312;
  wire[43:0] T313;
  wire[42:0] T314;
  wire[42:0] T315;
  wire[41:0] T316;
  wire[41:0] T317;
  wire[40:0] T318;
  wire[40:0] T319;
  wire[39:0] T320;
  wire[39:0] T321;
  wire[38:0] T322;
  wire[38:0] T323;
  wire[37:0] T324;
  wire[37:0] T325;
  wire[36:0] T326;
  wire[36:0] T327;
  wire[35:0] T328;
  wire[35:0] T329;
  wire[34:0] T330;
  wire[34:0] T331;
  wire[33:0] T332;
  wire[33:0] T333;
  wire[32:0] T334;
  wire[32:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[30:0] T338;
  wire[30:0] T339;
  wire[29:0] T340;
  wire[29:0] T341;
  wire[28:0] T342;
  wire[28:0] T343;
  wire[27:0] T344;
  wire[27:0] T345;
  wire[26:0] T346;
  wire[26:0] T347;
  wire[25:0] T348;
  wire[25:0] T349;
  wire[24:0] T350;
  wire[24:0] T351;
  wire[23:0] T352;
  wire[23:0] T353;
  wire[22:0] T354;
  wire[22:0] T355;
  wire[21:0] T356;
  wire[21:0] T357;
  wire[20:0] T358;
  wire[20:0] T359;
  wire[19:0] T360;
  wire[19:0] T361;
  wire[18:0] T362;
  wire[18:0] T363;
  wire[17:0] T364;
  wire[17:0] T365;
  wire[16:0] T366;
  wire[16:0] T367;
  wire[15:0] T368;
  wire[15:0] T369;
  wire[14:0] T370;
  wire[14:0] T371;
  wire[13:0] T372;
  wire[13:0] T373;
  wire[12:0] T374;
  wire[12:0] T375;
  wire[11:0] T376;
  wire[11:0] T377;
  wire[10:0] T378;
  wire[10:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[6:0] T386;
  wire[6:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[3:0] T393;
  wire[2:0] T394;
  wire[2:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[8:0] T428;
  wire[8:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[8:0] T468;
  wire[8:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[8:0] T508;
  wire[8:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[8:0] T548;
  wire[8:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[8:0] T588;
  wire[8:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[3:0] T625;
  wire[3:0] T626;
  wire[3:0] T627;
  wire[8:0] T628;
  wire[8:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[3:0] T665;
  wire[3:0] T666;
  wire[3:0] T667;
  wire[8:0] T668;
  wire[8:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[3:0] T705;
  wire[3:0] T706;
  wire[3:0] T707;
  wire[8:0] T708;
  wire[8:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[3:0] T745;
  wire[3:0] T746;
  wire[3:0] T747;
  wire[8:0] T748;
  wire[8:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire[1:0] T780;
  wire[1:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[3:0] T785;
  wire[3:0] T786;
  wire[3:0] T787;
  wire[8:0] T788;
  wire[8:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[8:0] T828;
  wire[8:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[3:0] T865;
  wire[3:0] T866;
  wire[3:0] T867;
  wire[8:0] T868;
  wire[8:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[3:0] T905;
  wire[3:0] T906;
  wire[3:0] T907;
  wire[8:0] T908;
  wire[8:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire[1:0] T940;
  wire[1:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[3:0] T945;
  wire[3:0] T946;
  wire[3:0] T947;
  wire[8:0] T948;
  wire[8:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[3:0] T985;
  wire[3:0] T986;
  wire[3:0] T987;
  wire[8:0] T988;
  wire[8:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire[3:0] T1025;
  wire[3:0] T1026;
  wire[3:0] T1027;
  wire[8:0] T1028;
  wire[8:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire[3:0] T1065;
  wire[3:0] T1066;
  wire[3:0] T1067;
  wire[8:0] T1068;
  wire[8:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire[1:0] T1092;
  wire[1:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[8:0] T1108;
  wire[8:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire[1:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire[1:0] T1140;
  wire[1:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[8:0] T1148;
  wire[8:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire[1:0] T1156;
  wire[1:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire[1:0] T1172;
  wire[1:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[8:0] T1188;
  wire[8:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[1:0] T1201;
  wire[1:0] T1202;
  wire[1:0] T1203;
  wire[2:0] T1204;
  wire[2:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[1:0] T1209;
  wire[1:0] T1210;
  wire[1:0] T1211;
  wire[2:0] T1212;
  wire[2:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[2:0] T1220;
  wire[2:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[1:0] T1225;
  wire[1:0] T1226;
  wire[1:0] T1227;
  wire[2:0] T1228;
  wire[2:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[1:0] T1233;
  wire[1:0] T1234;
  wire[1:0] T1235;
  wire[2:0] T1236;
  wire[2:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[1:0] T1241;
  wire[1:0] T1242;
  wire[1:0] T1243;
  wire[2:0] T1244;
  wire[2:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[1:0] T1249;
  wire[1:0] T1250;
  wire[1:0] T1251;
  wire[2:0] T1252;
  wire[2:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[1:0] T1257;
  wire[1:0] T1258;
  wire[1:0] T1259;
  wire[2:0] T1260;
  wire[2:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[1:0] T1265;
  wire[1:0] T1266;
  wire[1:0] T1267;
  wire[2:0] T1268;
  wire[2:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[1:0] T1273;
  wire[1:0] T1274;
  wire[1:0] T1275;
  wire[2:0] T1276;
  wire[2:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire[1:0] T1292;
  wire[1:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire[1:0] T1308;
  wire[1:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire[1:0] T1340;
  wire[1:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire[1:0] T1356;
  wire[1:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[2:0] T1364;
  wire[2:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[1:0] T1369;
  wire[1:0] T1370;
  wire[1:0] T1371;
  wire[2:0] T1372;
  wire[2:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[1:0] T1377;
  wire[1:0] T1378;
  wire[1:0] T1379;
  wire[2:0] T1380;
  wire[2:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[1:0] T1385;
  wire[1:0] T1386;
  wire[1:0] T1387;
  wire[2:0] T1388;
  wire[2:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[1:0] T1393;
  wire[1:0] T1394;
  wire[1:0] T1395;
  wire[2:0] T1396;
  wire[2:0] T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire[1:0] T1401;
  wire[1:0] T1402;
  wire[1:0] T1403;
  wire[2:0] T1404;
  wire[2:0] T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire[1:0] T1409;
  wire[1:0] T1410;
  wire[1:0] T1411;
  wire[2:0] T1412;
  wire[2:0] T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire[1:0] T1417;
  wire[1:0] T1418;
  wire[1:0] T1419;
  wire[2:0] T1420;
  wire[2:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire[1:0] T1425;
  wire[1:0] T1426;
  wire[1:0] T1427;
  wire[2:0] T1428;
  wire[2:0] T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire[1:0] T1433;
  wire[1:0] T1434;
  wire[1:0] T1435;
  wire[2:0] T1436;
  wire[2:0] T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire[1:0] T1444;
  wire[1:0] T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire[1:0] T1452;
  wire[1:0] T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire[1:0] T1468;
  wire[1:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire T1473;
  wire T1474;
  wire T1475;
  wire[1:0] T1476;
  wire[1:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire[1:0] T1484;
  wire[1:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire[1:0] T1492;
  wire[1:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire T1497;
  wire T1498;
  wire T1499;
  wire[1:0] T1500;
  wire[1:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire[1:0] T1508;
  wire[1:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire[1:0] T1516;
  wire[1:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[1:0] T1521;
  wire[1:0] T1522;
  wire[1:0] T1523;
  wire[2:0] T1524;
  wire[2:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[1:0] T1529;
  wire[1:0] T1530;
  wire[1:0] T1531;
  wire[2:0] T1532;
  wire[2:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[1:0] T1537;
  wire[1:0] T1538;
  wire[1:0] T1539;
  wire[2:0] T1540;
  wire[2:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[1:0] T1545;
  wire[1:0] T1546;
  wire[1:0] T1547;
  wire[2:0] T1548;
  wire[2:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[1:0] T1553;
  wire[1:0] T1554;
  wire[1:0] T1555;
  wire[2:0] T1556;
  wire[2:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[1:0] T1561;
  wire[1:0] T1562;
  wire[1:0] T1563;
  wire[2:0] T1564;
  wire[2:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[1:0] T1569;
  wire[1:0] T1570;
  wire[1:0] T1571;
  wire[2:0] T1572;
  wire[2:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[1:0] T1577;
  wire[1:0] T1578;
  wire[1:0] T1579;
  wire[2:0] T1580;
  wire[2:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[1:0] T1585;
  wire[1:0] T1586;
  wire[1:0] T1587;
  wire[2:0] T1588;
  wire[2:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[1:0] T1593;
  wire[1:0] T1594;
  wire[1:0] T1595;
  wire[2:0] T1596;
  wire[2:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire[1:0] T1604;
  wire[1:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[1:0] T1612;
  wire[1:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire[1:0] T1620;
  wire[1:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire[1:0] T1628;
  wire[1:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire[1:0] T1636;
  wire[1:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire[1:0] T1644;
  wire[1:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire[1:0] T1652;
  wire[1:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire[1:0] T1660;
  wire[1:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire T1665;
  wire T1666;
  wire T1667;
  wire[1:0] T1668;
  wire[1:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire[1:0] T1676;
  wire[1:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[10:0] T1684;
  wire[10:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[1:0] T1689;
  wire[1:0] T1690;
  wire[1:0] T1691;
  wire[2:0] T1692;
  wire[2:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[10:0] T1700;
  wire[10:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[1:0] T1705;
  wire[1:0] T1706;
  wire[1:0] T1707;
  wire[2:0] T1708;
  wire[2:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[10:0] T1716;
  wire[10:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[1:0] T1721;
  wire[1:0] T1722;
  wire[1:0] T1723;
  wire[2:0] T1724;
  wire[2:0] T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire[3:0] T1729;
  wire[3:0] T1730;
  wire[3:0] T1731;
  wire[10:0] T1732;
  wire[10:0] T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire[1:0] T1737;
  wire[1:0] T1738;
  wire[1:0] T1739;
  wire[2:0] T1740;
  wire[2:0] T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire[3:0] T1745;
  wire[3:0] T1746;
  wire[3:0] T1747;
  wire[10:0] T1748;
  wire[10:0] T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire[1:0] T1753;
  wire[1:0] T1754;
  wire[1:0] T1755;
  wire[2:0] T1756;
  wire[2:0] T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire[3:0] T1761;
  wire[3:0] T1762;
  wire[3:0] T1763;
  wire[10:0] T1764;
  wire[10:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire[1:0] T1769;
  wire[1:0] T1770;
  wire[1:0] T1771;
  wire[2:0] T1772;
  wire[2:0] T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire[3:0] T1777;
  wire[3:0] T1778;
  wire[3:0] T1779;
  wire[10:0] T1780;
  wire[10:0] T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire[1:0] T1785;
  wire[1:0] T1786;
  wire[1:0] T1787;
  wire[2:0] T1788;
  wire[2:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire[3:0] T1793;
  wire[3:0] T1794;
  wire[3:0] T1795;
  wire[10:0] T1796;
  wire[10:0] T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire[1:0] T1801;
  wire[1:0] T1802;
  wire[1:0] T1803;
  wire[2:0] T1804;
  wire[2:0] T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire[3:0] T1809;
  wire[3:0] T1810;
  wire[3:0] T1811;
  wire[10:0] T1812;
  wire[10:0] T1813;
  wire T1814;
  wire T1815;
  wire T1816;
  wire[1:0] T1817;
  wire[1:0] T1818;
  wire[1:0] T1819;
  wire[2:0] T1820;
  wire[2:0] T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[3:0] T1825;
  wire[3:0] T1826;
  wire[3:0] T1827;
  wire[10:0] T1828;
  wire[10:0] T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire[1:0] T1833;
  wire[1:0] T1834;
  wire[1:0] T1835;
  wire[2:0] T1836;
  wire[2:0] T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire[3:0] T1841;
  wire[3:0] T1842;
  wire[3:0] T1843;
  wire[10:0] T1844;
  wire[10:0] T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire T1851;
  wire[1:0] T1852;
  wire[1:0] T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire[3:0] T1857;
  wire[3:0] T1858;
  wire[3:0] T1859;
  wire[10:0] T1860;
  wire[10:0] T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[1:0] T1868;
  wire[1:0] T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire[3:0] T1873;
  wire[3:0] T1874;
  wire[3:0] T1875;
  wire[10:0] T1876;
  wire[10:0] T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire[3:0] T1889;
  wire[3:0] T1890;
  wire[3:0] T1891;
  wire[10:0] T1892;
  wire[10:0] T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[1:0] T1900;
  wire[1:0] T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire[3:0] T1905;
  wire[3:0] T1906;
  wire[3:0] T1907;
  wire[10:0] T1908;
  wire[10:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire[1:0] T1916;
  wire[1:0] T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire[3:0] T1921;
  wire[3:0] T1922;
  wire[3:0] T1923;
  wire[10:0] T1924;
  wire[10:0] T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire[1:0] T1932;
  wire[1:0] T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire[3:0] T1937;
  wire[3:0] T1938;
  wire[3:0] T1939;
  wire[10:0] T1940;
  wire[10:0] T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire T1947;
  wire[1:0] T1948;
  wire[1:0] T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire[3:0] T1953;
  wire[3:0] T1954;
  wire[3:0] T1955;
  wire[10:0] T1956;
  wire[10:0] T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire[1:0] T1964;
  wire[1:0] T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire[3:0] T1969;
  wire[3:0] T1970;
  wire[3:0] T1971;
  wire[10:0] T1972;
  wire[10:0] T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire[1:0] T1980;
  wire[1:0] T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire[3:0] T1985;
  wire[3:0] T1986;
  wire[3:0] T1987;
  wire[10:0] T1988;
  wire[10:0] T1989;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire[1:0] T1996;
  wire[1:0] T1997;
  wire[32:0] T1998;
  wire[32:0] T1999;
  wire[31:0] T2000;
  wire[31:0] T2001;
  wire[30:0] T2002;
  wire[30:0] T2003;
  wire[29:0] T2004;
  wire[29:0] T2005;
  wire[28:0] T2006;
  wire[28:0] T2007;
  wire[27:0] T2008;
  wire[27:0] T2009;
  wire[26:0] T2010;
  wire[26:0] T2011;
  wire[25:0] T2012;
  wire[25:0] T2013;
  wire[24:0] T2014;
  wire[24:0] T2015;
  wire[23:0] T2016;
  wire[23:0] T2017;
  wire[22:0] T2018;
  wire[22:0] T2019;
  wire[21:0] T2020;
  wire[21:0] T2021;
  wire[20:0] T2022;
  wire[20:0] T2023;
  wire[19:0] T2024;
  wire[19:0] T2025;
  wire[18:0] T2026;
  wire[18:0] T2027;
  wire[17:0] T2028;
  wire[17:0] T2029;
  wire[16:0] T2030;
  wire[16:0] T2031;
  wire[15:0] T2032;
  wire[15:0] T2033;
  wire[14:0] T2034;
  wire[14:0] T2035;
  wire[13:0] T2036;
  wire[13:0] T2037;
  wire[12:0] T2038;
  wire[12:0] T2039;
  wire[11:0] T2040;
  wire[11:0] T2041;
  wire[10:0] T2042;
  wire[10:0] T2043;
  wire[9:0] T2044;
  wire[9:0] T2045;
  wire[8:0] T2046;
  wire[8:0] T2047;
  wire[7:0] T2048;
  wire[7:0] T2049;
  wire[6:0] T2050;
  wire[6:0] T2051;
  wire[5:0] T2052;
  wire[5:0] T2053;
  wire[4:0] T2054;
  wire[4:0] T2055;
  wire[3:0] T2056;
  wire[3:0] T2057;
  wire[2:0] T2058;
  wire[2:0] T2059;
  wire[1:0] T2060;
  wire[1:0] T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire[3:0] T2065;
  wire[3:0] T2066;
  wire[3:0] T2067;
  wire[15:0] T2068;
  wire[15:0] T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire[3:0] T2073;
  wire[3:0] T2074;
  wire[3:0] T2075;
  wire[15:0] T2076;
  wire[15:0] T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[3:0] T2081;
  wire[3:0] T2082;
  wire[3:0] T2083;
  wire[15:0] T2084;
  wire[15:0] T2085;
  wire T2086;
  wire T2087;
  wire T2088;
  wire[3:0] T2089;
  wire[3:0] T2090;
  wire[3:0] T2091;
  wire[15:0] T2092;
  wire[15:0] T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire[3:0] T2097;
  wire[3:0] T2098;
  wire[3:0] T2099;
  wire[15:0] T2100;
  wire[15:0] T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire[3:0] T2105;
  wire[3:0] T2106;
  wire[3:0] T2107;
  wire[15:0] T2108;
  wire[15:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire[3:0] T2113;
  wire[3:0] T2114;
  wire[3:0] T2115;
  wire[15:0] T2116;
  wire[15:0] T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[3:0] T2121;
  wire[3:0] T2122;
  wire[3:0] T2123;
  wire[15:0] T2124;
  wire[15:0] T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire[3:0] T2129;
  wire[3:0] T2130;
  wire[3:0] T2131;
  wire[15:0] T2132;
  wire[15:0] T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire[3:0] T2137;
  wire[3:0] T2138;
  wire[3:0] T2139;
  wire[15:0] T2140;
  wire[15:0] T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire[3:0] T2145;
  wire[3:0] T2146;
  wire[3:0] T2147;
  wire[15:0] T2148;
  wire[15:0] T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire[3:0] T2153;
  wire[3:0] T2154;
  wire[3:0] T2155;
  wire[15:0] T2156;
  wire[15:0] T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire[3:0] T2161;
  wire[3:0] T2162;
  wire[3:0] T2163;
  wire[15:0] T2164;
  wire[15:0] T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire[3:0] T2169;
  wire[3:0] T2170;
  wire[3:0] T2171;
  wire[15:0] T2172;
  wire[15:0] T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  wire[3:0] T2177;
  wire[3:0] T2178;
  wire[3:0] T2179;
  wire[15:0] T2180;
  wire[15:0] T2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire[3:0] T2185;
  wire[3:0] T2186;
  wire[3:0] T2187;
  wire[15:0] T2188;
  wire[15:0] T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[3:0] T2193;
  wire[3:0] T2194;
  wire[3:0] T2195;
  wire[15:0] T2196;
  wire[15:0] T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire[3:0] T2201;
  wire[3:0] T2202;
  wire[3:0] T2203;
  wire[15:0] T2204;
  wire[15:0] T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire[3:0] T2209;
  wire[3:0] T2210;
  wire[3:0] T2211;
  wire[15:0] T2212;
  wire[15:0] T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire[3:0] T2217;
  wire[3:0] T2218;
  wire[3:0] T2219;
  wire[15:0] T2220;
  wire[15:0] T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire[3:0] T2225;
  wire[3:0] T2226;
  wire[3:0] T2227;
  wire[15:0] T2228;
  wire[15:0] T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire[3:0] T2233;
  wire[3:0] T2234;
  wire[3:0] T2235;
  wire[15:0] T2236;
  wire[15:0] T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire[3:0] T2241;
  wire[3:0] T2242;
  wire[3:0] T2243;
  wire[15:0] T2244;
  wire[15:0] T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  wire[3:0] T2249;
  wire[3:0] T2250;
  wire[3:0] T2251;
  wire[15:0] T2252;
  wire[15:0] T2253;
  wire T2254;
  wire T2255;
  wire T2256;
  wire[3:0] T2257;
  wire[3:0] T2258;
  wire[3:0] T2259;
  wire[15:0] T2260;
  wire[15:0] T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[3:0] T2265;
  wire[3:0] T2266;
  wire[3:0] T2267;
  wire[15:0] T2268;
  wire[15:0] T2269;
  wire T2270;
  wire T2271;
  wire T2272;
  wire[3:0] T2273;
  wire[3:0] T2274;
  wire[3:0] T2275;
  wire[15:0] T2276;
  wire[15:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire[3:0] T2281;
  wire[3:0] T2282;
  wire[3:0] T2283;
  wire[15:0] T2284;
  wire[15:0] T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire[3:0] T2289;
  wire[3:0] T2290;
  wire[3:0] T2291;
  wire[15:0] T2292;
  wire[15:0] T2293;
  wire T2294;
  wire T2295;
  wire T2296;
  wire[3:0] T2297;
  wire[3:0] T2298;
  wire[3:0] T2299;
  wire[15:0] T2300;
  wire[15:0] T2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire[3:0] T2305;
  wire[3:0] T2306;
  wire[3:0] T2307;
  wire[15:0] T2308;
  wire[15:0] T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire[3:0] T2313;
  wire[3:0] T2314;
  wire[3:0] T2315;
  wire[15:0] T2316;
  wire[15:0] T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  wire[3:0] T2321;
  wire[3:0] T2322;
  wire[3:0] T2323;
  wire[15:0] T2324;
  wire[15:0] T2325;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1990, T2};
  assign T2 = T3;
  assign T3 = {T1982, T4};
  assign T4 = T5;
  assign T5 = {T1974, T6};
  assign T6 = T7;
  assign T7 = {T1966, T8};
  assign T8 = T9;
  assign T9 = {T1958, T10};
  assign T10 = T11;
  assign T11 = {T1950, T12};
  assign T12 = T13;
  assign T13 = {T1942, T14};
  assign T14 = T15;
  assign T15 = {T1934, T16};
  assign T16 = T17;
  assign T17 = {T1926, T18};
  assign T18 = T19;
  assign T19 = {T1918, T20};
  assign T20 = T21;
  assign T21 = {T1910, T22};
  assign T22 = T23;
  assign T23 = {T1902, T24};
  assign T24 = T25;
  assign T25 = {T1894, T26};
  assign T26 = T27;
  assign T27 = {T1886, T28};
  assign T28 = T29;
  assign T29 = {T1878, T30};
  assign T30 = T31;
  assign T31 = {T1870, T32};
  assign T32 = T33;
  assign T33 = {T1862, T34};
  assign T34 = T35;
  assign T35 = {T1854, T36};
  assign T36 = T37;
  assign T37 = {T1846, T38};
  assign T38 = T39;
  assign T39 = {T1838, T40};
  assign T40 = T41;
  assign T41 = {T1830, T42};
  assign T42 = T43;
  assign T43 = {T1822, T44};
  assign T44 = T45;
  assign T45 = {T1814, T46};
  assign T46 = T47;
  assign T47 = {T1806, T48};
  assign T48 = T49;
  assign T49 = {T1798, T50};
  assign T50 = T51;
  assign T51 = {T1790, T52};
  assign T52 = T53;
  assign T53 = {T1782, T54};
  assign T54 = T55;
  assign T55 = {T1774, T56};
  assign T56 = T57;
  assign T57 = {T1766, T58};
  assign T58 = T59;
  assign T59 = {T1758, T60};
  assign T60 = T61;
  assign T61 = {T1750, T62};
  assign T62 = T63;
  assign T63 = {T1742, T64};
  assign T64 = T65;
  assign T65 = {T1734, T66};
  assign T66 = T67;
  assign T67 = {T1726, T68};
  assign T68 = T69;
  assign T69 = {T1718, T70};
  assign T70 = T71;
  assign T71 = {T1710, T72};
  assign T72 = T73;
  assign T73 = {T1702, T74};
  assign T74 = T75;
  assign T75 = {T1694, T76};
  assign T76 = T77;
  assign T77 = {T1686, T78};
  assign T78 = T79;
  assign T79 = {T1678, T80};
  assign T80 = T81;
  assign T81 = {T1670, T82};
  assign T82 = T83;
  assign T83 = {T1662, T84};
  assign T84 = T85;
  assign T85 = {T1654, T86};
  assign T86 = T87;
  assign T87 = {T1646, T88};
  assign T88 = T89;
  assign T89 = {T1638, T90};
  assign T90 = T91;
  assign T91 = {T1630, T92};
  assign T92 = T93;
  assign T93 = {T1622, T94};
  assign T94 = T95;
  assign T95 = {T1614, T96};
  assign T96 = T97;
  assign T97 = {T1606, T98};
  assign T98 = T99;
  assign T99 = {T1598, T100};
  assign T100 = T101;
  assign T101 = {T1590, T102};
  assign T102 = T103;
  assign T103 = {T1582, T104};
  assign T104 = T105;
  assign T105 = {T1574, T106};
  assign T106 = T107;
  assign T107 = {T1566, T108};
  assign T108 = T109;
  assign T109 = {T1558, T110};
  assign T110 = T111;
  assign T111 = {T1550, T112};
  assign T112 = T113;
  assign T113 = {T1542, T114};
  assign T114 = T115;
  assign T115 = {T1534, T116};
  assign T116 = T117;
  assign T117 = {T1526, T118};
  assign T118 = T119;
  assign T119 = {T1518, T120};
  assign T120 = T121;
  assign T121 = {T1510, T122};
  assign T122 = T123;
  assign T123 = {T1502, T124};
  assign T124 = T125;
  assign T125 = {T1494, T126};
  assign T126 = T127;
  assign T127 = {T1486, T128};
  assign T128 = T129;
  assign T129 = {T1478, T130};
  assign T130 = T131;
  assign T131 = {T1470, T132};
  assign T132 = T133;
  assign T133 = {T1462, T134};
  assign T134 = T135;
  assign T135 = {T1454, T136};
  assign T136 = T137;
  assign T137 = {T1446, T138};
  assign T138 = T139;
  assign T139 = {T1438, T140};
  assign T140 = T141;
  assign T141 = {T1430, T142};
  assign T142 = T143;
  assign T143 = {T1422, T144};
  assign T144 = T145;
  assign T145 = {T1414, T146};
  assign T146 = T147;
  assign T147 = {T1406, T148};
  assign T148 = T149;
  assign T149 = {T1398, T150};
  assign T150 = T151;
  assign T151 = {T1390, T152};
  assign T152 = T153;
  assign T153 = {T1382, T154};
  assign T154 = T155;
  assign T155 = {T1374, T156};
  assign T156 = T157;
  assign T157 = {T1366, T158};
  assign T158 = T159;
  assign T159 = {T1358, T160};
  assign T160 = T161;
  assign T161 = {T1350, T162};
  assign T162 = T163;
  assign T163 = {T1342, T164};
  assign T164 = T165;
  assign T165 = {T1334, T166};
  assign T166 = T167;
  assign T167 = {T1326, T168};
  assign T168 = T169;
  assign T169 = {T1318, T170};
  assign T170 = T171;
  assign T171 = {T1310, T172};
  assign T172 = T173;
  assign T173 = {T1302, T174};
  assign T174 = T175;
  assign T175 = {T1294, T176};
  assign T176 = T177;
  assign T177 = {T1286, T178};
  assign T178 = T179;
  assign T179 = {T1278, T180};
  assign T180 = T181;
  assign T181 = {T1270, T182};
  assign T182 = T183;
  assign T183 = {T1262, T184};
  assign T184 = T185;
  assign T185 = {T1254, T186};
  assign T186 = T187;
  assign T187 = {T1246, T188};
  assign T188 = T189;
  assign T189 = {T1238, T190};
  assign T190 = T191;
  assign T191 = {T1230, T192};
  assign T192 = T193;
  assign T193 = {T1222, T194};
  assign T194 = T195;
  assign T195 = {T1214, T196};
  assign T196 = T197;
  assign T197 = {T1206, T198};
  assign T198 = T199;
  assign T199 = {T1198, T200};
  assign T200 = T201;
  assign T201 = {T1190, T202};
  assign T202 = T203;
  assign T203 = {T1182, T204};
  assign T204 = T205;
  assign T205 = {T1174, T206};
  assign T206 = T207;
  assign T207 = {T1166, T208};
  assign T208 = T209;
  assign T209 = {T1158, T210};
  assign T210 = T211;
  assign T211 = {T1150, T212};
  assign T212 = T213;
  assign T213 = {T1142, T214};
  assign T214 = T215;
  assign T215 = {T1134, T216};
  assign T216 = T217;
  assign T217 = {T1126, T218};
  assign T218 = T219;
  assign T219 = {T1118, T220};
  assign T220 = T221;
  assign T221 = {T1110, T222};
  assign T222 = T223;
  assign T223 = {T1102, T224};
  assign T224 = T225;
  assign T225 = {T1094, T226};
  assign T226 = T227;
  assign T227 = {T1086, T228};
  assign T228 = T229;
  assign T229 = {T1078, T230};
  assign T230 = T231;
  assign T231 = {T1070, T232};
  assign T232 = T233;
  assign T233 = {T1062, T234};
  assign T234 = T235;
  assign T235 = {T1054, T236};
  assign T236 = T237;
  assign T237 = {T1046, T238};
  assign T238 = T239;
  assign T239 = {T1038, T240};
  assign T240 = T241;
  assign T241 = {T1030, T242};
  assign T242 = T243;
  assign T243 = {T1022, T244};
  assign T244 = T245;
  assign T245 = {T1014, T246};
  assign T246 = T247;
  assign T247 = {T1006, T248};
  assign T248 = T249;
  assign T249 = {T998, T250};
  assign T250 = T251;
  assign T251 = {T990, T252};
  assign T252 = T253;
  assign T253 = {T982, T254};
  assign T254 = T255;
  assign T255 = {T974, T256};
  assign T256 = T257;
  assign T257 = {T966, T258};
  assign T258 = T259;
  assign T259 = {T958, T260};
  assign T260 = T261;
  assign T261 = {T950, T262};
  assign T262 = T263;
  assign T263 = {T942, T264};
  assign T264 = T265;
  assign T265 = {T934, T266};
  assign T266 = T267;
  assign T267 = {T926, T268};
  assign T268 = T269;
  assign T269 = {T918, T270};
  assign T270 = T271;
  assign T271 = {T910, T272};
  assign T272 = T273;
  assign T273 = {T902, T274};
  assign T274 = T275;
  assign T275 = {T894, T276};
  assign T276 = T277;
  assign T277 = {T886, T278};
  assign T278 = T279;
  assign T279 = {T878, T280};
  assign T280 = T281;
  assign T281 = {T870, T282};
  assign T282 = T283;
  assign T283 = {T862, T284};
  assign T284 = T285;
  assign T285 = {T854, T286};
  assign T286 = T287;
  assign T287 = {T846, T288};
  assign T288 = T289;
  assign T289 = {T838, T290};
  assign T290 = T291;
  assign T291 = {T830, T292};
  assign T292 = T293;
  assign T293 = {T822, T294};
  assign T294 = T295;
  assign T295 = {T814, T296};
  assign T296 = T297;
  assign T297 = {T806, T298};
  assign T298 = T299;
  assign T299 = {T798, T300};
  assign T300 = T301;
  assign T301 = {T790, T302};
  assign T302 = T303;
  assign T303 = {T782, T304};
  assign T304 = T305;
  assign T305 = {T774, T306};
  assign T306 = T307;
  assign T307 = {T766, T308};
  assign T308 = T309;
  assign T309 = {T758, T310};
  assign T310 = T311;
  assign T311 = {T750, T312};
  assign T312 = T313;
  assign T313 = {T742, T314};
  assign T314 = T315;
  assign T315 = {T734, T316};
  assign T316 = T317;
  assign T317 = {T726, T318};
  assign T318 = T319;
  assign T319 = {T718, T320};
  assign T320 = T321;
  assign T321 = {T710, T322};
  assign T322 = T323;
  assign T323 = {T702, T324};
  assign T324 = T325;
  assign T325 = {T694, T326};
  assign T326 = T327;
  assign T327 = {T686, T328};
  assign T328 = T329;
  assign T329 = {T678, T330};
  assign T330 = T331;
  assign T331 = {T670, T332};
  assign T332 = T333;
  assign T333 = {T662, T334};
  assign T334 = T335;
  assign T335 = {T654, T336};
  assign T336 = T337;
  assign T337 = {T646, T338};
  assign T338 = T339;
  assign T339 = {T638, T340};
  assign T340 = T341;
  assign T341 = {T630, T342};
  assign T342 = T343;
  assign T343 = {T622, T344};
  assign T344 = T345;
  assign T345 = {T614, T346};
  assign T346 = T347;
  assign T347 = {T606, T348};
  assign T348 = T349;
  assign T349 = {T598, T350};
  assign T350 = T351;
  assign T351 = {T590, T352};
  assign T352 = T353;
  assign T353 = {T582, T354};
  assign T354 = T355;
  assign T355 = {T574, T356};
  assign T356 = T357;
  assign T357 = {T566, T358};
  assign T358 = T359;
  assign T359 = {T558, T360};
  assign T360 = T361;
  assign T361 = {T550, T362};
  assign T362 = T363;
  assign T363 = {T542, T364};
  assign T364 = T365;
  assign T365 = {T534, T366};
  assign T366 = T367;
  assign T367 = {T526, T368};
  assign T368 = T369;
  assign T369 = {T518, T370};
  assign T370 = T371;
  assign T371 = {T510, T372};
  assign T372 = T373;
  assign T373 = {T502, T374};
  assign T374 = T375;
  assign T375 = {T494, T376};
  assign T376 = T377;
  assign T377 = {T486, T378};
  assign T378 = T379;
  assign T379 = {T478, T380};
  assign T380 = T381;
  assign T381 = {T470, T382};
  assign T382 = T383;
  assign T383 = {T462, T384};
  assign T384 = T385;
  assign T385 = {T454, T386};
  assign T386 = T387;
  assign T387 = {T446, T388};
  assign T388 = T389;
  assign T389 = {T438, T390};
  assign T390 = T391;
  assign T391 = {T430, T392};
  assign T392 = T393;
  assign T393 = {T422, T394};
  assign T394 = T395;
  assign T395 = {T414, T396};
  assign T396 = T397;
  assign T397 = {T406, T398};
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[2'h2/* 2*/:2'h2/* 2*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[3'h5/* 5*/:3'h4/* 4*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[3'h6/* 6*/:2'h3/* 3*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[4'he/* 14*/:3'h6/* 6*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[5'h10/* 16*/:4'hf/* 15*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[5'h12/* 18*/:5'h11/* 17*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[5'h14/* 20*/:5'h13/* 19*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[5'h16/* 22*/:5'h15/* 21*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[4'he/* 14*/:4'hb/* 11*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[5'h1f/* 31*/:5'h17/* 23*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[5'h16/* 22*/:5'h13/* 19*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[6'h30/* 48*/:6'h28/* 40*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[6'h32/* 50*/:6'h31/* 49*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[6'h34/* 52*/:6'h33/* 51*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[6'h36/* 54*/:6'h35/* 53*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[6'h38/* 56*/:6'h37/* 55*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[5'h1e/* 30*/:5'h1b/* 27*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[7'h41/* 65*/:6'h39/* 57*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h26/* 38*/:6'h23/* 35*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[7'h52/* 82*/:7'h4a/* 74*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h54/* 84*/:7'h53/* 83*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h56/* 86*/:7'h55/* 85*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h58/* 88*/:7'h57/* 87*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h5a/* 90*/:7'h59/* 89*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[6'h2e/* 46*/:6'h2b/* 43*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[7'h63/* 99*/:7'h5b/* 91*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[6'h2f/* 47*/:6'h2f/* 47*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[6'h36/* 54*/:6'h33/* 51*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h74/* 116*/:7'h6c/* 108*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[7'h76/* 118*/:7'h75/* 117*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[7'h78/* 120*/:7'h77/* 119*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[7'h7a/* 122*/:7'h79/* 121*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[7'h7c/* 124*/:7'h7b/* 123*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[6'h3e/* 62*/:6'h3b/* 59*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'h85/* 133*/:7'h7d/* 125*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[6'h3f/* 63*/:6'h3f/* 63*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'h87/* 135*/:8'h86/* 134*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h41/* 65*/:7'h41/* 65*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h42/* 66*/:7'h42/* 66*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h46/* 70*/:7'h43/* 67*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'h96/* 150*/:8'h8e/* 142*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h47/* 71*/:7'h47/* 71*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'h98/* 152*/:8'h97/* 151*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h48/* 72*/:7'h48/* 72*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'h9a/* 154*/:8'h99/* 153*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h49/* 73*/:7'h49/* 73*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'h9c/* 156*/:8'h9b/* 155*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'h9e/* 158*/:8'h9d/* 157*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'ha7/* 167*/:8'h9f/* 159*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'hab/* 171*/:8'haa/* 170*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'had/* 173*/:8'hac/* 172*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'haf/* 175*/:8'hae/* 174*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h56/* 86*/:7'h53/* 83*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'hb8/* 184*/:8'hb0/* 176*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'hba/* 186*/:8'hb9/* 185*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'hbc/* 188*/:8'hbb/* 187*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[8'hbe/* 190*/:8'hbd/* 189*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[7'h5a/* 90*/:7'h5a/* 90*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[8'hc0/* 192*/:8'hbf/* 191*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[7'h5e/* 94*/:7'h5b/* 91*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[8'hc9/* 201*/:8'hc1/* 193*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[7'h5f/* 95*/:7'h5f/* 95*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[8'hcb/* 203*/:8'hca/* 202*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[7'h60/* 96*/:7'h60/* 96*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[7'h61/* 97*/:7'h61/* 97*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[8'hcf/* 207*/:8'hce/* 206*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[7'h62/* 98*/:7'h62/* 98*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[7'h66/* 102*/:7'h63/* 99*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[8'hda/* 218*/:8'hd2/* 210*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[7'h67/* 103*/:7'h67/* 103*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[8'hdc/* 220*/:8'hdb/* 219*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[8'hde/* 222*/:8'hdd/* 221*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[7'h69/* 105*/:7'h69/* 105*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[8'he0/* 224*/:8'hdf/* 223*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[7'h6a/* 106*/:7'h6a/* 106*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[8'he2/* 226*/:8'he1/* 225*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[7'h6e/* 110*/:7'h6b/* 107*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[8'heb/* 235*/:8'he3/* 227*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[7'h6f/* 111*/:7'h6f/* 111*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[8'hed/* 237*/:8'hec/* 236*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[7'h70/* 112*/:7'h70/* 112*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[8'hef/* 239*/:8'hee/* 238*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[7'h71/* 113*/:7'h71/* 113*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[8'hf3/* 243*/:8'hf2/* 242*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[8'hfc/* 252*/:8'hf4/* 244*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[8'hfe/* 254*/:8'hfd/* 253*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[7'h78/* 120*/:7'h78/* 120*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h100/* 256*/:8'hff/* 255*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[7'h79/* 121*/:7'h79/* 121*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h102/* 258*/:9'h101/* 257*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[7'h7a/* 122*/:7'h7a/* 122*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h104/* 260*/:9'h103/* 259*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[7'h7e/* 126*/:7'h7b/* 123*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h10d/* 269*/:9'h105/* 261*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[7'h7f/* 127*/:7'h7f/* 127*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'h80/* 128*/:8'h80/* 128*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h113/* 275*/:9'h112/* 274*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'h82/* 130*/:8'h82/* 130*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h115/* 277*/:9'h114/* 276*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'h86/* 134*/:8'h83/* 131*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h11e/* 286*/:9'h116/* 278*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'h87/* 135*/:8'h87/* 135*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h120/* 288*/:9'h11f/* 287*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'h88/* 136*/:8'h88/* 136*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h122/* 290*/:9'h121/* 289*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'h89/* 137*/:8'h89/* 137*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h124/* 292*/:9'h123/* 291*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'h8a/* 138*/:8'h8a/* 138*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h126/* 294*/:9'h125/* 293*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'h8e/* 142*/:8'h8b/* 139*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h12f/* 303*/:9'h127/* 295*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'h8f/* 143*/:8'h8f/* 143*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h131/* 305*/:9'h130/* 304*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h133/* 307*/:9'h132/* 306*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'h91/* 145*/:8'h91/* 145*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h135/* 309*/:9'h134/* 308*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'h92/* 146*/:8'h92/* 146*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h137/* 311*/:9'h136/* 310*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'h96/* 150*/:8'h93/* 147*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[9'h140/* 320*/:9'h138/* 312*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'h97/* 151*/:8'h97/* 151*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[9'h142/* 322*/:9'h141/* 321*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'h98/* 152*/:8'h98/* 152*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[9'h144/* 324*/:9'h143/* 323*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'h99/* 153*/:8'h99/* 153*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[9'h146/* 326*/:9'h145/* 325*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[9'h151/* 337*/:9'h149/* 329*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[9'h156/* 342*/:9'h154/* 340*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[9'h159/* 345*/:9'h157/* 343*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[9'h15c/* 348*/:9'h15a/* 346*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[9'h15f/* 351*/:9'h15d/* 349*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[9'h162/* 354*/:9'h160/* 352*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[9'h165/* 357*/:9'h163/* 355*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[9'h168/* 360*/:9'h166/* 358*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[9'h16b/* 363*/:9'h169/* 361*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[9'h16e/* 366*/:9'h16c/* 364*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[9'h171/* 369*/:9'h16f/* 367*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[8'hb4/* 180*/:8'hb4/* 180*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[9'h173/* 371*/:9'h172/* 370*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[9'h175/* 373*/:9'h174/* 372*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[9'h177/* 375*/:9'h176/* 374*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[8'hb7/* 183*/:8'hb7/* 183*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[9'h179/* 377*/:9'h178/* 376*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[9'h17b/* 379*/:9'h17a/* 378*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[9'h17d/* 381*/:9'h17c/* 380*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[9'h17f/* 383*/:9'h17e/* 382*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[8'hbb/* 187*/:8'hbb/* 187*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[9'h181/* 385*/:9'h180/* 384*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[8'hbc/* 188*/:8'hbc/* 188*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[9'h183/* 387*/:9'h182/* 386*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[9'h185/* 389*/:9'h184/* 388*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[9'h188/* 392*/:9'h186/* 390*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[8'hc1/* 193*/:8'hc0/* 192*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[9'h18b/* 395*/:9'h189/* 393*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[8'hc3/* 195*/:8'hc2/* 194*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[9'h18e/* 398*/:9'h18c/* 396*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[9'h191/* 401*/:9'h18f/* 399*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[9'h194/* 404*/:9'h192/* 402*/];
  assign T1398 = T1399;
  assign T1399 = T1400;
  assign T1400 = T1404[T1401];
  assign T1401 = T1402;
  assign T1402 = T1403;
  assign T1403 = io_chanxy_config[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T1404 = T1405;
  assign T1405 = io_chanxy_in[9'h197/* 407*/:9'h195/* 405*/];
  assign T1406 = T1407;
  assign T1407 = T1408;
  assign T1408 = T1412[T1409];
  assign T1409 = T1410;
  assign T1410 = T1411;
  assign T1411 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T1412 = T1413;
  assign T1413 = io_chanxy_in[9'h19a/* 410*/:9'h198/* 408*/];
  assign T1414 = T1415;
  assign T1415 = T1416;
  assign T1416 = T1420[T1417];
  assign T1417 = T1418;
  assign T1418 = T1419;
  assign T1419 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T1420 = T1421;
  assign T1421 = io_chanxy_in[9'h19d/* 413*/:9'h19b/* 411*/];
  assign T1422 = T1423;
  assign T1423 = T1424;
  assign T1424 = T1428[T1425];
  assign T1425 = T1426;
  assign T1426 = T1427;
  assign T1427 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T1428 = T1429;
  assign T1429 = io_chanxy_in[9'h1a0/* 416*/:9'h19e/* 414*/];
  assign T1430 = T1431;
  assign T1431 = T1432;
  assign T1432 = T1436[T1433];
  assign T1433 = T1434;
  assign T1434 = T1435;
  assign T1435 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T1436 = T1437;
  assign T1437 = io_chanxy_in[9'h1a3/* 419*/:9'h1a1/* 417*/];
  assign T1438 = T1439;
  assign T1439 = T1440;
  assign T1440 = T1444[T1441];
  assign T1441 = T1442;
  assign T1442 = T1443;
  assign T1443 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T1444 = T1445;
  assign T1445 = io_chanxy_in[9'h1a5/* 421*/:9'h1a4/* 420*/];
  assign T1446 = T1447;
  assign T1447 = T1448;
  assign T1448 = T1452[T1449];
  assign T1449 = T1450;
  assign T1450 = T1451;
  assign T1451 = io_chanxy_config[8'hd3/* 211*/:8'hd3/* 211*/];
  assign T1452 = T1453;
  assign T1453 = io_chanxy_in[9'h1a7/* 423*/:9'h1a6/* 422*/];
  assign T1454 = T1455;
  assign T1455 = T1456;
  assign T1456 = T1460[T1457];
  assign T1457 = T1458;
  assign T1458 = T1459;
  assign T1459 = io_chanxy_config[8'hd4/* 212*/:8'hd4/* 212*/];
  assign T1460 = T1461;
  assign T1461 = io_chanxy_in[9'h1a9/* 425*/:9'h1a8/* 424*/];
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_chanxy_config[8'hd5/* 213*/:8'hd5/* 213*/];
  assign T1468 = T1469;
  assign T1469 = io_chanxy_in[9'h1ab/* 427*/:9'h1aa/* 426*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T1476 = T1477;
  assign T1477 = io_chanxy_in[9'h1ad/* 429*/:9'h1ac/* 428*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T1484 = T1485;
  assign T1485 = io_chanxy_in[9'h1af/* 431*/:9'h1ae/* 430*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T1492 = T1493;
  assign T1493 = io_chanxy_in[9'h1b1/* 433*/:9'h1b0/* 432*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T1500 = T1501;
  assign T1501 = io_chanxy_in[9'h1b3/* 435*/:9'h1b2/* 434*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T1508 = T1509;
  assign T1509 = io_chanxy_in[9'h1b5/* 437*/:9'h1b4/* 436*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T1516 = T1517;
  assign T1517 = io_chanxy_in[9'h1b7/* 439*/:9'h1b6/* 438*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_chanxy_config[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T1524 = T1525;
  assign T1525 = io_chanxy_in[9'h1ba/* 442*/:9'h1b8/* 440*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T1532 = T1533;
  assign T1533 = io_chanxy_in[9'h1bd/* 445*/:9'h1bb/* 443*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_chanxy_config[8'he1/* 225*/:8'he0/* 224*/];
  assign T1540 = T1541;
  assign T1541 = io_chanxy_in[9'h1c0/* 448*/:9'h1be/* 446*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_chanxy_config[8'he3/* 227*/:8'he2/* 226*/];
  assign T1548 = T1549;
  assign T1549 = io_chanxy_in[9'h1c3/* 451*/:9'h1c1/* 449*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_chanxy_config[8'he5/* 229*/:8'he4/* 228*/];
  assign T1556 = T1557;
  assign T1557 = io_chanxy_in[9'h1c6/* 454*/:9'h1c4/* 452*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_chanxy_config[8'he7/* 231*/:8'he6/* 230*/];
  assign T1564 = T1565;
  assign T1565 = io_chanxy_in[9'h1c9/* 457*/:9'h1c7/* 455*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_chanxy_config[8'he9/* 233*/:8'he8/* 232*/];
  assign T1572 = T1573;
  assign T1573 = io_chanxy_in[9'h1cc/* 460*/:9'h1ca/* 458*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_chanxy_config[8'heb/* 235*/:8'hea/* 234*/];
  assign T1580 = T1581;
  assign T1581 = io_chanxy_in[9'h1cf/* 463*/:9'h1cd/* 461*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_chanxy_config[8'hed/* 237*/:8'hec/* 236*/];
  assign T1588 = T1589;
  assign T1589 = io_chanxy_in[9'h1d2/* 466*/:9'h1d0/* 464*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_chanxy_config[8'hef/* 239*/:8'hee/* 238*/];
  assign T1596 = T1597;
  assign T1597 = io_chanxy_in[9'h1d5/* 469*/:9'h1d3/* 467*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T1604 = T1605;
  assign T1605 = io_chanxy_in[9'h1d7/* 471*/:9'h1d6/* 470*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T1612 = T1613;
  assign T1613 = io_chanxy_in[9'h1d9/* 473*/:9'h1d8/* 472*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1620 = T1621;
  assign T1621 = io_chanxy_in[9'h1db/* 475*/:9'h1da/* 474*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T1628 = T1629;
  assign T1629 = io_chanxy_in[9'h1dd/* 477*/:9'h1dc/* 476*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_chanxy_config[8'hf4/* 244*/:8'hf4/* 244*/];
  assign T1636 = T1637;
  assign T1637 = io_chanxy_in[9'h1df/* 479*/:9'h1de/* 478*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_chanxy_config[8'hf5/* 245*/:8'hf5/* 245*/];
  assign T1644 = T1645;
  assign T1645 = io_chanxy_in[9'h1e1/* 481*/:9'h1e0/* 480*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_chanxy_config[8'hf6/* 246*/:8'hf6/* 246*/];
  assign T1652 = T1653;
  assign T1653 = io_chanxy_in[9'h1e3/* 483*/:9'h1e2/* 482*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T1660 = T1661;
  assign T1661 = io_chanxy_in[9'h1e5/* 485*/:9'h1e4/* 484*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1668 = T1669;
  assign T1669 = io_chanxy_in[9'h1e7/* 487*/:9'h1e6/* 486*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T1676 = T1677;
  assign T1677 = io_chanxy_in[9'h1e9/* 489*/:9'h1e8/* 488*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_chanxy_config[8'hfd/* 253*/:8'hfa/* 250*/];
  assign T1684 = T1685;
  assign T1685 = io_chanxy_in[9'h1f4/* 500*/:9'h1ea/* 490*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_chanxy_config[8'hff/* 255*/:8'hfe/* 254*/];
  assign T1692 = T1693;
  assign T1693 = io_chanxy_in[9'h1f7/* 503*/:9'h1f5/* 501*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1700 = T1701;
  assign T1701 = io_chanxy_in[10'h202/* 514*/:9'h1f8/* 504*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_chanxy_config[9'h105/* 261*/:9'h104/* 260*/];
  assign T1708 = T1709;
  assign T1709 = io_chanxy_in[10'h205/* 517*/:10'h203/* 515*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_chanxy_config[9'h109/* 265*/:9'h106/* 262*/];
  assign T1716 = T1717;
  assign T1717 = io_chanxy_in[10'h210/* 528*/:10'h206/* 518*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_chanxy_config[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T1724 = T1725;
  assign T1725 = io_chanxy_in[10'h213/* 531*/:10'h211/* 529*/];
  assign T1726 = T1727;
  assign T1727 = T1728;
  assign T1728 = T1732[T1729];
  assign T1729 = T1730;
  assign T1730 = T1731;
  assign T1731 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1732 = T1733;
  assign T1733 = io_chanxy_in[10'h21e/* 542*/:10'h214/* 532*/];
  assign T1734 = T1735;
  assign T1735 = T1736;
  assign T1736 = T1740[T1737];
  assign T1737 = T1738;
  assign T1738 = T1739;
  assign T1739 = io_chanxy_config[9'h111/* 273*/:9'h110/* 272*/];
  assign T1740 = T1741;
  assign T1741 = io_chanxy_in[10'h221/* 545*/:10'h21f/* 543*/];
  assign T1742 = T1743;
  assign T1743 = T1744;
  assign T1744 = T1748[T1745];
  assign T1745 = T1746;
  assign T1746 = T1747;
  assign T1747 = io_chanxy_config[9'h115/* 277*/:9'h112/* 274*/];
  assign T1748 = T1749;
  assign T1749 = io_chanxy_in[10'h22c/* 556*/:10'h222/* 546*/];
  assign T1750 = T1751;
  assign T1751 = T1752;
  assign T1752 = T1756[T1753];
  assign T1753 = T1754;
  assign T1754 = T1755;
  assign T1755 = io_chanxy_config[9'h117/* 279*/:9'h116/* 278*/];
  assign T1756 = T1757;
  assign T1757 = io_chanxy_in[10'h22f/* 559*/:10'h22d/* 557*/];
  assign T1758 = T1759;
  assign T1759 = T1760;
  assign T1760 = T1764[T1761];
  assign T1761 = T1762;
  assign T1762 = T1763;
  assign T1763 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1764 = T1765;
  assign T1765 = io_chanxy_in[10'h23a/* 570*/:10'h230/* 560*/];
  assign T1766 = T1767;
  assign T1767 = T1768;
  assign T1768 = T1772[T1769];
  assign T1769 = T1770;
  assign T1770 = T1771;
  assign T1771 = io_chanxy_config[9'h11d/* 285*/:9'h11c/* 284*/];
  assign T1772 = T1773;
  assign T1773 = io_chanxy_in[10'h23d/* 573*/:10'h23b/* 571*/];
  assign T1774 = T1775;
  assign T1775 = T1776;
  assign T1776 = T1780[T1777];
  assign T1777 = T1778;
  assign T1778 = T1779;
  assign T1779 = io_chanxy_config[9'h121/* 289*/:9'h11e/* 286*/];
  assign T1780 = T1781;
  assign T1781 = io_chanxy_in[10'h248/* 584*/:10'h23e/* 574*/];
  assign T1782 = T1783;
  assign T1783 = T1784;
  assign T1784 = T1788[T1785];
  assign T1785 = T1786;
  assign T1786 = T1787;
  assign T1787 = io_chanxy_config[9'h123/* 291*/:9'h122/* 290*/];
  assign T1788 = T1789;
  assign T1789 = io_chanxy_in[10'h24b/* 587*/:10'h249/* 585*/];
  assign T1790 = T1791;
  assign T1791 = T1792;
  assign T1792 = T1796[T1793];
  assign T1793 = T1794;
  assign T1794 = T1795;
  assign T1795 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1796 = T1797;
  assign T1797 = io_chanxy_in[10'h256/* 598*/:10'h24c/* 588*/];
  assign T1798 = T1799;
  assign T1799 = T1800;
  assign T1800 = T1804[T1801];
  assign T1801 = T1802;
  assign T1802 = T1803;
  assign T1803 = io_chanxy_config[9'h129/* 297*/:9'h128/* 296*/];
  assign T1804 = T1805;
  assign T1805 = io_chanxy_in[10'h259/* 601*/:10'h257/* 599*/];
  assign T1806 = T1807;
  assign T1807 = T1808;
  assign T1808 = T1812[T1809];
  assign T1809 = T1810;
  assign T1810 = T1811;
  assign T1811 = io_chanxy_config[9'h12d/* 301*/:9'h12a/* 298*/];
  assign T1812 = T1813;
  assign T1813 = io_chanxy_in[10'h264/* 612*/:10'h25a/* 602*/];
  assign T1814 = T1815;
  assign T1815 = T1816;
  assign T1816 = T1820[T1817];
  assign T1817 = T1818;
  assign T1818 = T1819;
  assign T1819 = io_chanxy_config[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T1820 = T1821;
  assign T1821 = io_chanxy_in[10'h267/* 615*/:10'h265/* 613*/];
  assign T1822 = T1823;
  assign T1823 = T1824;
  assign T1824 = T1828[T1825];
  assign T1825 = T1826;
  assign T1826 = T1827;
  assign T1827 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1828 = T1829;
  assign T1829 = io_chanxy_in[10'h272/* 626*/:10'h268/* 616*/];
  assign T1830 = T1831;
  assign T1831 = T1832;
  assign T1832 = T1836[T1833];
  assign T1833 = T1834;
  assign T1834 = T1835;
  assign T1835 = io_chanxy_config[9'h135/* 309*/:9'h134/* 308*/];
  assign T1836 = T1837;
  assign T1837 = io_chanxy_in[10'h275/* 629*/:10'h273/* 627*/];
  assign T1838 = T1839;
  assign T1839 = T1840;
  assign T1840 = T1844[T1841];
  assign T1841 = T1842;
  assign T1842 = T1843;
  assign T1843 = io_chanxy_config[9'h139/* 313*/:9'h136/* 310*/];
  assign T1844 = T1845;
  assign T1845 = io_chanxy_in[10'h280/* 640*/:10'h276/* 630*/];
  assign T1846 = T1847;
  assign T1847 = T1848;
  assign T1848 = T1852[T1849];
  assign T1849 = T1850;
  assign T1850 = T1851;
  assign T1851 = io_chanxy_config[9'h13a/* 314*/:9'h13a/* 314*/];
  assign T1852 = T1853;
  assign T1853 = io_chanxy_in[10'h282/* 642*/:10'h281/* 641*/];
  assign T1854 = T1855;
  assign T1855 = T1856;
  assign T1856 = T1860[T1857];
  assign T1857 = T1858;
  assign T1858 = T1859;
  assign T1859 = io_chanxy_config[9'h13e/* 318*/:9'h13b/* 315*/];
  assign T1860 = T1861;
  assign T1861 = io_chanxy_in[10'h28d/* 653*/:10'h283/* 643*/];
  assign T1862 = T1863;
  assign T1863 = T1864;
  assign T1864 = T1868[T1865];
  assign T1865 = T1866;
  assign T1866 = T1867;
  assign T1867 = io_chanxy_config[9'h13f/* 319*/:9'h13f/* 319*/];
  assign T1868 = T1869;
  assign T1869 = io_chanxy_in[10'h28f/* 655*/:10'h28e/* 654*/];
  assign T1870 = T1871;
  assign T1871 = T1872;
  assign T1872 = T1876[T1873];
  assign T1873 = T1874;
  assign T1874 = T1875;
  assign T1875 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1876 = T1877;
  assign T1877 = io_chanxy_in[10'h29a/* 666*/:10'h290/* 656*/];
  assign T1878 = T1879;
  assign T1879 = T1880;
  assign T1880 = T1884[T1881];
  assign T1881 = T1882;
  assign T1882 = T1883;
  assign T1883 = io_chanxy_config[9'h144/* 324*/:9'h144/* 324*/];
  assign T1884 = T1885;
  assign T1885 = io_chanxy_in[10'h29c/* 668*/:10'h29b/* 667*/];
  assign T1886 = T1887;
  assign T1887 = T1888;
  assign T1888 = T1892[T1889];
  assign T1889 = T1890;
  assign T1890 = T1891;
  assign T1891 = io_chanxy_config[9'h148/* 328*/:9'h145/* 325*/];
  assign T1892 = T1893;
  assign T1893 = io_chanxy_in[10'h2a7/* 679*/:10'h29d/* 669*/];
  assign T1894 = T1895;
  assign T1895 = T1896;
  assign T1896 = T1900[T1897];
  assign T1897 = T1898;
  assign T1898 = T1899;
  assign T1899 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1900 = T1901;
  assign T1901 = io_chanxy_in[10'h2a9/* 681*/:10'h2a8/* 680*/];
  assign T1902 = T1903;
  assign T1903 = T1904;
  assign T1904 = T1908[T1905];
  assign T1905 = T1906;
  assign T1906 = T1907;
  assign T1907 = io_chanxy_config[9'h14d/* 333*/:9'h14a/* 330*/];
  assign T1908 = T1909;
  assign T1909 = io_chanxy_in[10'h2b4/* 692*/:10'h2aa/* 682*/];
  assign T1910 = T1911;
  assign T1911 = T1912;
  assign T1912 = T1916[T1913];
  assign T1913 = T1914;
  assign T1914 = T1915;
  assign T1915 = io_chanxy_config[9'h14e/* 334*/:9'h14e/* 334*/];
  assign T1916 = T1917;
  assign T1917 = io_chanxy_in[10'h2b6/* 694*/:10'h2b5/* 693*/];
  assign T1918 = T1919;
  assign T1919 = T1920;
  assign T1920 = T1924[T1921];
  assign T1921 = T1922;
  assign T1922 = T1923;
  assign T1923 = io_chanxy_config[9'h152/* 338*/:9'h14f/* 335*/];
  assign T1924 = T1925;
  assign T1925 = io_chanxy_in[10'h2c1/* 705*/:10'h2b7/* 695*/];
  assign T1926 = T1927;
  assign T1927 = T1928;
  assign T1928 = T1932[T1929];
  assign T1929 = T1930;
  assign T1930 = T1931;
  assign T1931 = io_chanxy_config[9'h153/* 339*/:9'h153/* 339*/];
  assign T1932 = T1933;
  assign T1933 = io_chanxy_in[10'h2c3/* 707*/:10'h2c2/* 706*/];
  assign T1934 = T1935;
  assign T1935 = T1936;
  assign T1936 = T1940[T1937];
  assign T1937 = T1938;
  assign T1938 = T1939;
  assign T1939 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1940 = T1941;
  assign T1941 = io_chanxy_in[10'h2ce/* 718*/:10'h2c4/* 708*/];
  assign T1942 = T1943;
  assign T1943 = T1944;
  assign T1944 = T1948[T1945];
  assign T1945 = T1946;
  assign T1946 = T1947;
  assign T1947 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1948 = T1949;
  assign T1949 = io_chanxy_in[10'h2d0/* 720*/:10'h2cf/* 719*/];
  assign T1950 = T1951;
  assign T1951 = T1952;
  assign T1952 = T1956[T1953];
  assign T1953 = T1954;
  assign T1954 = T1955;
  assign T1955 = io_chanxy_config[9'h15c/* 348*/:9'h159/* 345*/];
  assign T1956 = T1957;
  assign T1957 = io_chanxy_in[10'h2db/* 731*/:10'h2d1/* 721*/];
  assign T1958 = T1959;
  assign T1959 = T1960;
  assign T1960 = T1964[T1961];
  assign T1961 = T1962;
  assign T1962 = T1963;
  assign T1963 = io_chanxy_config[9'h15d/* 349*/:9'h15d/* 349*/];
  assign T1964 = T1965;
  assign T1965 = io_chanxy_in[10'h2dd/* 733*/:10'h2dc/* 732*/];
  assign T1966 = T1967;
  assign T1967 = T1968;
  assign T1968 = T1972[T1969];
  assign T1969 = T1970;
  assign T1970 = T1971;
  assign T1971 = io_chanxy_config[9'h161/* 353*/:9'h15e/* 350*/];
  assign T1972 = T1973;
  assign T1973 = io_chanxy_in[10'h2e8/* 744*/:10'h2de/* 734*/];
  assign T1974 = T1975;
  assign T1975 = T1976;
  assign T1976 = T1980[T1977];
  assign T1977 = T1978;
  assign T1978 = T1979;
  assign T1979 = io_chanxy_config[9'h162/* 354*/:9'h162/* 354*/];
  assign T1980 = T1981;
  assign T1981 = io_chanxy_in[10'h2ea/* 746*/:10'h2e9/* 745*/];
  assign T1982 = T1983;
  assign T1983 = T1984;
  assign T1984 = T1988[T1985];
  assign T1985 = T1986;
  assign T1986 = T1987;
  assign T1987 = io_chanxy_config[9'h166/* 358*/:9'h163/* 355*/];
  assign T1988 = T1989;
  assign T1989 = io_chanxy_in[10'h2f5/* 757*/:10'h2eb/* 747*/];
  assign T1990 = T1991;
  assign T1991 = T1992;
  assign T1992 = T1996[T1993];
  assign T1993 = T1994;
  assign T1994 = T1995;
  assign T1995 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1996 = T1997;
  assign T1997 = io_chanxy_in[10'h2f7/* 759*/:10'h2f6/* 758*/];
  assign io_ipin_out = T1998;
  assign T1998 = T1999;
  assign T1999 = {T2318, T2000};
  assign T2000 = T2001;
  assign T2001 = {T2310, T2002};
  assign T2002 = T2003;
  assign T2003 = {T2302, T2004};
  assign T2004 = T2005;
  assign T2005 = {T2294, T2006};
  assign T2006 = T2007;
  assign T2007 = {T2286, T2008};
  assign T2008 = T2009;
  assign T2009 = {T2278, T2010};
  assign T2010 = T2011;
  assign T2011 = {T2270, T2012};
  assign T2012 = T2013;
  assign T2013 = {T2262, T2014};
  assign T2014 = T2015;
  assign T2015 = {T2254, T2016};
  assign T2016 = T2017;
  assign T2017 = {T2246, T2018};
  assign T2018 = T2019;
  assign T2019 = {T2238, T2020};
  assign T2020 = T2021;
  assign T2021 = {T2230, T2022};
  assign T2022 = T2023;
  assign T2023 = {T2222, T2024};
  assign T2024 = T2025;
  assign T2025 = {T2214, T2026};
  assign T2026 = T2027;
  assign T2027 = {T2206, T2028};
  assign T2028 = T2029;
  assign T2029 = {T2198, T2030};
  assign T2030 = T2031;
  assign T2031 = {T2190, T2032};
  assign T2032 = T2033;
  assign T2033 = {T2182, T2034};
  assign T2034 = T2035;
  assign T2035 = {T2174, T2036};
  assign T2036 = T2037;
  assign T2037 = {T2166, T2038};
  assign T2038 = T2039;
  assign T2039 = {T2158, T2040};
  assign T2040 = T2041;
  assign T2041 = {T2150, T2042};
  assign T2042 = T2043;
  assign T2043 = {T2142, T2044};
  assign T2044 = T2045;
  assign T2045 = {T2134, T2046};
  assign T2046 = T2047;
  assign T2047 = {T2126, T2048};
  assign T2048 = T2049;
  assign T2049 = {T2118, T2050};
  assign T2050 = T2051;
  assign T2051 = {T2110, T2052};
  assign T2052 = T2053;
  assign T2053 = {T2102, T2054};
  assign T2054 = T2055;
  assign T2055 = {T2094, T2056};
  assign T2056 = T2057;
  assign T2057 = {T2086, T2058};
  assign T2058 = T2059;
  assign T2059 = {T2078, T2060};
  assign T2060 = T2061;
  assign T2061 = {T2070, T2062};
  assign T2062 = T2063;
  assign T2063 = T2064;
  assign T2064 = T2068[T2065];
  assign T2065 = T2066;
  assign T2066 = T2067;
  assign T2067 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T2068 = T2069;
  assign T2069 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T2070 = T2071;
  assign T2071 = T2072;
  assign T2072 = T2076[T2073];
  assign T2073 = T2074;
  assign T2074 = T2075;
  assign T2075 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T2076 = T2077;
  assign T2077 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T2078 = T2079;
  assign T2079 = T2080;
  assign T2080 = T2084[T2081];
  assign T2081 = T2082;
  assign T2082 = T2083;
  assign T2083 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T2084 = T2085;
  assign T2085 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T2086 = T2087;
  assign T2087 = T2088;
  assign T2088 = T2092[T2089];
  assign T2089 = T2090;
  assign T2090 = T2091;
  assign T2091 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T2092 = T2093;
  assign T2093 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T2094 = T2095;
  assign T2095 = T2096;
  assign T2096 = T2100[T2097];
  assign T2097 = T2098;
  assign T2098 = T2099;
  assign T2099 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T2100 = T2101;
  assign T2101 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T2102 = T2103;
  assign T2103 = T2104;
  assign T2104 = T2108[T2105];
  assign T2105 = T2106;
  assign T2106 = T2107;
  assign T2107 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T2108 = T2109;
  assign T2109 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T2110 = T2111;
  assign T2111 = T2112;
  assign T2112 = T2116[T2113];
  assign T2113 = T2114;
  assign T2114 = T2115;
  assign T2115 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T2116 = T2117;
  assign T2117 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T2118 = T2119;
  assign T2119 = T2120;
  assign T2120 = T2124[T2121];
  assign T2121 = T2122;
  assign T2122 = T2123;
  assign T2123 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T2124 = T2125;
  assign T2125 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T2126 = T2127;
  assign T2127 = T2128;
  assign T2128 = T2132[T2129];
  assign T2129 = T2130;
  assign T2130 = T2131;
  assign T2131 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T2132 = T2133;
  assign T2133 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T2134 = T2135;
  assign T2135 = T2136;
  assign T2136 = T2140[T2137];
  assign T2137 = T2138;
  assign T2138 = T2139;
  assign T2139 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T2140 = T2141;
  assign T2141 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T2142 = T2143;
  assign T2143 = T2144;
  assign T2144 = T2148[T2145];
  assign T2145 = T2146;
  assign T2146 = T2147;
  assign T2147 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T2148 = T2149;
  assign T2149 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T2150 = T2151;
  assign T2151 = T2152;
  assign T2152 = T2156[T2153];
  assign T2153 = T2154;
  assign T2154 = T2155;
  assign T2155 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T2156 = T2157;
  assign T2157 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T2158 = T2159;
  assign T2159 = T2160;
  assign T2160 = T2164[T2161];
  assign T2161 = T2162;
  assign T2162 = T2163;
  assign T2163 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T2164 = T2165;
  assign T2165 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T2166 = T2167;
  assign T2167 = T2168;
  assign T2168 = T2172[T2169];
  assign T2169 = T2170;
  assign T2170 = T2171;
  assign T2171 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T2172 = T2173;
  assign T2173 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T2174 = T2175;
  assign T2175 = T2176;
  assign T2176 = T2180[T2177];
  assign T2177 = T2178;
  assign T2178 = T2179;
  assign T2179 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T2180 = T2181;
  assign T2181 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T2182 = T2183;
  assign T2183 = T2184;
  assign T2184 = T2188[T2185];
  assign T2185 = T2186;
  assign T2186 = T2187;
  assign T2187 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T2188 = T2189;
  assign T2189 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T2190 = T2191;
  assign T2191 = T2192;
  assign T2192 = T2196[T2193];
  assign T2193 = T2194;
  assign T2194 = T2195;
  assign T2195 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T2196 = T2197;
  assign T2197 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T2198 = T2199;
  assign T2199 = T2200;
  assign T2200 = T2204[T2201];
  assign T2201 = T2202;
  assign T2202 = T2203;
  assign T2203 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T2204 = T2205;
  assign T2205 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T2206 = T2207;
  assign T2207 = T2208;
  assign T2208 = T2212[T2209];
  assign T2209 = T2210;
  assign T2210 = T2211;
  assign T2211 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T2212 = T2213;
  assign T2213 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T2214 = T2215;
  assign T2215 = T2216;
  assign T2216 = T2220[T2217];
  assign T2217 = T2218;
  assign T2218 = T2219;
  assign T2219 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T2220 = T2221;
  assign T2221 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T2222 = T2223;
  assign T2223 = T2224;
  assign T2224 = T2228[T2225];
  assign T2225 = T2226;
  assign T2226 = T2227;
  assign T2227 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T2228 = T2229;
  assign T2229 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T2230 = T2231;
  assign T2231 = T2232;
  assign T2232 = T2236[T2233];
  assign T2233 = T2234;
  assign T2234 = T2235;
  assign T2235 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T2236 = T2237;
  assign T2237 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T2238 = T2239;
  assign T2239 = T2240;
  assign T2240 = T2244[T2241];
  assign T2241 = T2242;
  assign T2242 = T2243;
  assign T2243 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T2244 = T2245;
  assign T2245 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T2246 = T2247;
  assign T2247 = T2248;
  assign T2248 = T2252[T2249];
  assign T2249 = T2250;
  assign T2250 = T2251;
  assign T2251 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T2252 = T2253;
  assign T2253 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T2254 = T2255;
  assign T2255 = T2256;
  assign T2256 = T2260[T2257];
  assign T2257 = T2258;
  assign T2258 = T2259;
  assign T2259 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T2260 = T2261;
  assign T2261 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T2262 = T2263;
  assign T2263 = T2264;
  assign T2264 = T2268[T2265];
  assign T2265 = T2266;
  assign T2266 = T2267;
  assign T2267 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T2268 = T2269;
  assign T2269 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T2270 = T2271;
  assign T2271 = T2272;
  assign T2272 = T2276[T2273];
  assign T2273 = T2274;
  assign T2274 = T2275;
  assign T2275 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T2276 = T2277;
  assign T2277 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T2278 = T2279;
  assign T2279 = T2280;
  assign T2280 = T2284[T2281];
  assign T2281 = T2282;
  assign T2282 = T2283;
  assign T2283 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T2284 = T2285;
  assign T2285 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T2286 = T2287;
  assign T2287 = T2288;
  assign T2288 = T2292[T2289];
  assign T2289 = T2290;
  assign T2290 = T2291;
  assign T2291 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T2292 = T2293;
  assign T2293 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T2294 = T2295;
  assign T2295 = T2296;
  assign T2296 = T2300[T2297];
  assign T2297 = T2298;
  assign T2298 = T2299;
  assign T2299 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T2300 = T2301;
  assign T2301 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T2302 = T2303;
  assign T2303 = T2304;
  assign T2304 = T2308[T2305];
  assign T2305 = T2306;
  assign T2306 = T2307;
  assign T2307 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T2308 = T2309;
  assign T2309 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T2310 = T2311;
  assign T2311 = T2312;
  assign T2312 = T2316[T2313];
  assign T2313 = T2314;
  assign T2314 = T2315;
  assign T2315 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T2316 = T2317;
  assign T2317 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T2318 = T2319;
  assign T2319 = T2320;
  assign T2320 = T2324[T2321];
  assign T2321 = T2322;
  assign T2322 = T2323;
  assign T2323 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T2324 = T2325;
  assign T2325 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_4(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [759:0] io_chanxy_in,
    output[199:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[199:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_4 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


module sbcb_sp_5(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [775:0] io_chanxy_in,
    input [367:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[199:0] io_chanxy_out);

  wire[199:0] T0;
  wire[199:0] T1;
  wire[198:0] T2;
  wire[198:0] T3;
  wire[197:0] T4;
  wire[197:0] T5;
  wire[196:0] T6;
  wire[196:0] T7;
  wire[195:0] T8;
  wire[195:0] T9;
  wire[194:0] T10;
  wire[194:0] T11;
  wire[193:0] T12;
  wire[193:0] T13;
  wire[192:0] T14;
  wire[192:0] T15;
  wire[191:0] T16;
  wire[191:0] T17;
  wire[190:0] T18;
  wire[190:0] T19;
  wire[189:0] T20;
  wire[189:0] T21;
  wire[188:0] T22;
  wire[188:0] T23;
  wire[187:0] T24;
  wire[187:0] T25;
  wire[186:0] T26;
  wire[186:0] T27;
  wire[185:0] T28;
  wire[185:0] T29;
  wire[184:0] T30;
  wire[184:0] T31;
  wire[183:0] T32;
  wire[183:0] T33;
  wire[182:0] T34;
  wire[182:0] T35;
  wire[181:0] T36;
  wire[181:0] T37;
  wire[180:0] T38;
  wire[180:0] T39;
  wire[179:0] T40;
  wire[179:0] T41;
  wire[178:0] T42;
  wire[178:0] T43;
  wire[177:0] T44;
  wire[177:0] T45;
  wire[176:0] T46;
  wire[176:0] T47;
  wire[175:0] T48;
  wire[175:0] T49;
  wire[174:0] T50;
  wire[174:0] T51;
  wire[173:0] T52;
  wire[173:0] T53;
  wire[172:0] T54;
  wire[172:0] T55;
  wire[171:0] T56;
  wire[171:0] T57;
  wire[170:0] T58;
  wire[170:0] T59;
  wire[169:0] T60;
  wire[169:0] T61;
  wire[168:0] T62;
  wire[168:0] T63;
  wire[167:0] T64;
  wire[167:0] T65;
  wire[166:0] T66;
  wire[166:0] T67;
  wire[165:0] T68;
  wire[165:0] T69;
  wire[164:0] T70;
  wire[164:0] T71;
  wire[163:0] T72;
  wire[163:0] T73;
  wire[162:0] T74;
  wire[162:0] T75;
  wire[161:0] T76;
  wire[161:0] T77;
  wire[160:0] T78;
  wire[160:0] T79;
  wire[159:0] T80;
  wire[159:0] T81;
  wire[158:0] T82;
  wire[158:0] T83;
  wire[157:0] T84;
  wire[157:0] T85;
  wire[156:0] T86;
  wire[156:0] T87;
  wire[155:0] T88;
  wire[155:0] T89;
  wire[154:0] T90;
  wire[154:0] T91;
  wire[153:0] T92;
  wire[153:0] T93;
  wire[152:0] T94;
  wire[152:0] T95;
  wire[151:0] T96;
  wire[151:0] T97;
  wire[150:0] T98;
  wire[150:0] T99;
  wire[149:0] T100;
  wire[149:0] T101;
  wire[148:0] T102;
  wire[148:0] T103;
  wire[147:0] T104;
  wire[147:0] T105;
  wire[146:0] T106;
  wire[146:0] T107;
  wire[145:0] T108;
  wire[145:0] T109;
  wire[144:0] T110;
  wire[144:0] T111;
  wire[143:0] T112;
  wire[143:0] T113;
  wire[142:0] T114;
  wire[142:0] T115;
  wire[141:0] T116;
  wire[141:0] T117;
  wire[140:0] T118;
  wire[140:0] T119;
  wire[139:0] T120;
  wire[139:0] T121;
  wire[138:0] T122;
  wire[138:0] T123;
  wire[137:0] T124;
  wire[137:0] T125;
  wire[136:0] T126;
  wire[136:0] T127;
  wire[135:0] T128;
  wire[135:0] T129;
  wire[134:0] T130;
  wire[134:0] T131;
  wire[133:0] T132;
  wire[133:0] T133;
  wire[132:0] T134;
  wire[132:0] T135;
  wire[131:0] T136;
  wire[131:0] T137;
  wire[130:0] T138;
  wire[130:0] T139;
  wire[129:0] T140;
  wire[129:0] T141;
  wire[128:0] T142;
  wire[128:0] T143;
  wire[127:0] T144;
  wire[127:0] T145;
  wire[126:0] T146;
  wire[126:0] T147;
  wire[125:0] T148;
  wire[125:0] T149;
  wire[124:0] T150;
  wire[124:0] T151;
  wire[123:0] T152;
  wire[123:0] T153;
  wire[122:0] T154;
  wire[122:0] T155;
  wire[121:0] T156;
  wire[121:0] T157;
  wire[120:0] T158;
  wire[120:0] T159;
  wire[119:0] T160;
  wire[119:0] T161;
  wire[118:0] T162;
  wire[118:0] T163;
  wire[117:0] T164;
  wire[117:0] T165;
  wire[116:0] T166;
  wire[116:0] T167;
  wire[115:0] T168;
  wire[115:0] T169;
  wire[114:0] T170;
  wire[114:0] T171;
  wire[113:0] T172;
  wire[113:0] T173;
  wire[112:0] T174;
  wire[112:0] T175;
  wire[111:0] T176;
  wire[111:0] T177;
  wire[110:0] T178;
  wire[110:0] T179;
  wire[109:0] T180;
  wire[109:0] T181;
  wire[108:0] T182;
  wire[108:0] T183;
  wire[107:0] T184;
  wire[107:0] T185;
  wire[106:0] T186;
  wire[106:0] T187;
  wire[105:0] T188;
  wire[105:0] T189;
  wire[104:0] T190;
  wire[104:0] T191;
  wire[103:0] T192;
  wire[103:0] T193;
  wire[102:0] T194;
  wire[102:0] T195;
  wire[101:0] T196;
  wire[101:0] T197;
  wire[100:0] T198;
  wire[100:0] T199;
  wire[99:0] T200;
  wire[99:0] T201;
  wire[98:0] T202;
  wire[98:0] T203;
  wire[97:0] T204;
  wire[97:0] T205;
  wire[96:0] T206;
  wire[96:0] T207;
  wire[95:0] T208;
  wire[95:0] T209;
  wire[94:0] T210;
  wire[94:0] T211;
  wire[93:0] T212;
  wire[93:0] T213;
  wire[92:0] T214;
  wire[92:0] T215;
  wire[91:0] T216;
  wire[91:0] T217;
  wire[90:0] T218;
  wire[90:0] T219;
  wire[89:0] T220;
  wire[89:0] T221;
  wire[88:0] T222;
  wire[88:0] T223;
  wire[87:0] T224;
  wire[87:0] T225;
  wire[86:0] T226;
  wire[86:0] T227;
  wire[85:0] T228;
  wire[85:0] T229;
  wire[84:0] T230;
  wire[84:0] T231;
  wire[83:0] T232;
  wire[83:0] T233;
  wire[82:0] T234;
  wire[82:0] T235;
  wire[81:0] T236;
  wire[81:0] T237;
  wire[80:0] T238;
  wire[80:0] T239;
  wire[79:0] T240;
  wire[79:0] T241;
  wire[78:0] T242;
  wire[78:0] T243;
  wire[77:0] T244;
  wire[77:0] T245;
  wire[76:0] T246;
  wire[76:0] T247;
  wire[75:0] T248;
  wire[75:0] T249;
  wire[74:0] T250;
  wire[74:0] T251;
  wire[73:0] T252;
  wire[73:0] T253;
  wire[72:0] T254;
  wire[72:0] T255;
  wire[71:0] T256;
  wire[71:0] T257;
  wire[70:0] T258;
  wire[70:0] T259;
  wire[69:0] T260;
  wire[69:0] T261;
  wire[68:0] T262;
  wire[68:0] T263;
  wire[67:0] T264;
  wire[67:0] T265;
  wire[66:0] T266;
  wire[66:0] T267;
  wire[65:0] T268;
  wire[65:0] T269;
  wire[64:0] T270;
  wire[64:0] T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[62:0] T274;
  wire[62:0] T275;
  wire[61:0] T276;
  wire[61:0] T277;
  wire[60:0] T278;
  wire[60:0] T279;
  wire[59:0] T280;
  wire[59:0] T281;
  wire[58:0] T282;
  wire[58:0] T283;
  wire[57:0] T284;
  wire[57:0] T285;
  wire[56:0] T286;
  wire[56:0] T287;
  wire[55:0] T288;
  wire[55:0] T289;
  wire[54:0] T290;
  wire[54:0] T291;
  wire[53:0] T292;
  wire[53:0] T293;
  wire[52:0] T294;
  wire[52:0] T295;
  wire[51:0] T296;
  wire[51:0] T297;
  wire[50:0] T298;
  wire[50:0] T299;
  wire[49:0] T300;
  wire[49:0] T301;
  wire[48:0] T302;
  wire[48:0] T303;
  wire[47:0] T304;
  wire[47:0] T305;
  wire[46:0] T306;
  wire[46:0] T307;
  wire[45:0] T308;
  wire[45:0] T309;
  wire[44:0] T310;
  wire[44:0] T311;
  wire[43:0] T312;
  wire[43:0] T313;
  wire[42:0] T314;
  wire[42:0] T315;
  wire[41:0] T316;
  wire[41:0] T317;
  wire[40:0] T318;
  wire[40:0] T319;
  wire[39:0] T320;
  wire[39:0] T321;
  wire[38:0] T322;
  wire[38:0] T323;
  wire[37:0] T324;
  wire[37:0] T325;
  wire[36:0] T326;
  wire[36:0] T327;
  wire[35:0] T328;
  wire[35:0] T329;
  wire[34:0] T330;
  wire[34:0] T331;
  wire[33:0] T332;
  wire[33:0] T333;
  wire[32:0] T334;
  wire[32:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[30:0] T338;
  wire[30:0] T339;
  wire[29:0] T340;
  wire[29:0] T341;
  wire[28:0] T342;
  wire[28:0] T343;
  wire[27:0] T344;
  wire[27:0] T345;
  wire[26:0] T346;
  wire[26:0] T347;
  wire[25:0] T348;
  wire[25:0] T349;
  wire[24:0] T350;
  wire[24:0] T351;
  wire[23:0] T352;
  wire[23:0] T353;
  wire[22:0] T354;
  wire[22:0] T355;
  wire[21:0] T356;
  wire[21:0] T357;
  wire[20:0] T358;
  wire[20:0] T359;
  wire[19:0] T360;
  wire[19:0] T361;
  wire[18:0] T362;
  wire[18:0] T363;
  wire[17:0] T364;
  wire[17:0] T365;
  wire[16:0] T366;
  wire[16:0] T367;
  wire[15:0] T368;
  wire[15:0] T369;
  wire[14:0] T370;
  wire[14:0] T371;
  wire[13:0] T372;
  wire[13:0] T373;
  wire[12:0] T374;
  wire[12:0] T375;
  wire[11:0] T376;
  wire[11:0] T377;
  wire[10:0] T378;
  wire[10:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[6:0] T386;
  wire[6:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[3:0] T393;
  wire[2:0] T394;
  wire[2:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[1:0] T401;
  wire[1:0] T402;
  wire[1:0] T403;
  wire[2:0] T404;
  wire[2:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[1:0] T409;
  wire[1:0] T410;
  wire[1:0] T411;
  wire[2:0] T412;
  wire[2:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[1:0] T417;
  wire[1:0] T418;
  wire[1:0] T419;
  wire[2:0] T420;
  wire[2:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[1:0] T425;
  wire[1:0] T426;
  wire[1:0] T427;
  wire[2:0] T428;
  wire[2:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[1:0] T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[2:0] T436;
  wire[2:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[1:0] T449;
  wire[1:0] T450;
  wire[1:0] T451;
  wire[2:0] T452;
  wire[2:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[1:0] T457;
  wire[1:0] T458;
  wire[1:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[1:0] T467;
  wire[2:0] T468;
  wire[2:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire[1:0] T475;
  wire[2:0] T476;
  wire[2:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[1:0] T561;
  wire[1:0] T562;
  wire[1:0] T563;
  wire[2:0] T564;
  wire[2:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[1:0] T569;
  wire[1:0] T570;
  wire[1:0] T571;
  wire[2:0] T572;
  wire[2:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[1:0] T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[2:0] T580;
  wire[2:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[1:0] T585;
  wire[1:0] T586;
  wire[1:0] T587;
  wire[2:0] T588;
  wire[2:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[1:0] T593;
  wire[1:0] T594;
  wire[1:0] T595;
  wire[2:0] T596;
  wire[2:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[2:0] T724;
  wire[2:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[1:0] T729;
  wire[1:0] T730;
  wire[1:0] T731;
  wire[2:0] T732;
  wire[2:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[1:0] T737;
  wire[1:0] T738;
  wire[1:0] T739;
  wire[2:0] T740;
  wire[2:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[1:0] T745;
  wire[1:0] T746;
  wire[1:0] T747;
  wire[2:0] T748;
  wire[2:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[1:0] T753;
  wire[1:0] T754;
  wire[1:0] T755;
  wire[2:0] T756;
  wire[2:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[1:0] T777;
  wire[1:0] T778;
  wire[1:0] T779;
  wire[2:0] T780;
  wire[2:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[1:0] T793;
  wire[1:0] T794;
  wire[1:0] T795;
  wire[2:0] T796;
  wire[2:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[3:0] T881;
  wire[3:0] T882;
  wire[3:0] T883;
  wire[10:0] T884;
  wire[10:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[1:0] T889;
  wire[1:0] T890;
  wire[1:0] T891;
  wire[2:0] T892;
  wire[2:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[10:0] T900;
  wire[10:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[1:0] T905;
  wire[1:0] T906;
  wire[1:0] T907;
  wire[2:0] T908;
  wire[2:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[3:0] T913;
  wire[3:0] T914;
  wire[3:0] T915;
  wire[10:0] T916;
  wire[10:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire[1:0] T922;
  wire[1:0] T923;
  wire[2:0] T924;
  wire[2:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[3:0] T929;
  wire[3:0] T930;
  wire[3:0] T931;
  wire[10:0] T932;
  wire[10:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[1:0] T937;
  wire[1:0] T938;
  wire[1:0] T939;
  wire[2:0] T940;
  wire[2:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[3:0] T945;
  wire[3:0] T946;
  wire[3:0] T947;
  wire[10:0] T948;
  wire[10:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[1:0] T953;
  wire[1:0] T954;
  wire[1:0] T955;
  wire[2:0] T956;
  wire[2:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[3:0] T961;
  wire[3:0] T962;
  wire[3:0] T963;
  wire[10:0] T964;
  wire[10:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[1:0] T969;
  wire[1:0] T970;
  wire[1:0] T971;
  wire[2:0] T972;
  wire[2:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[10:0] T980;
  wire[10:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[1:0] T985;
  wire[1:0] T986;
  wire[1:0] T987;
  wire[2:0] T988;
  wire[2:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[3:0] T993;
  wire[3:0] T994;
  wire[3:0] T995;
  wire[10:0] T996;
  wire[10:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire[1:0] T1001;
  wire[1:0] T1002;
  wire[1:0] T1003;
  wire[2:0] T1004;
  wire[2:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire[3:0] T1009;
  wire[3:0] T1010;
  wire[3:0] T1011;
  wire[10:0] T1012;
  wire[10:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire[1:0] T1017;
  wire[1:0] T1018;
  wire[1:0] T1019;
  wire[2:0] T1020;
  wire[2:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire[3:0] T1025;
  wire[3:0] T1026;
  wire[3:0] T1027;
  wire[10:0] T1028;
  wire[10:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[1:0] T1033;
  wire[1:0] T1034;
  wire[1:0] T1035;
  wire[2:0] T1036;
  wire[2:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire[3:0] T1041;
  wire[3:0] T1042;
  wire[3:0] T1043;
  wire[10:0] T1044;
  wire[10:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire[3:0] T1057;
  wire[3:0] T1058;
  wire[3:0] T1059;
  wire[10:0] T1060;
  wire[10:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire[3:0] T1073;
  wire[3:0] T1074;
  wire[3:0] T1075;
  wire[10:0] T1076;
  wire[10:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[10:0] T1092;
  wire[10:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[10:0] T1108;
  wire[10:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[10:0] T1124;
  wire[10:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[10:0] T1140;
  wire[10:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire[1:0] T1148;
  wire[1:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[10:0] T1156;
  wire[10:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[10:0] T1172;
  wire[10:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[10:0] T1188;
  wire[10:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[1:0] T1201;
  wire[1:0] T1202;
  wire[1:0] T1203;
  wire[2:0] T1204;
  wire[2:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[1:0] T1209;
  wire[1:0] T1210;
  wire[1:0] T1211;
  wire[2:0] T1212;
  wire[2:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[2:0] T1220;
  wire[2:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[9:0] T1228;
  wire[9:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[1:0] T1233;
  wire[1:0] T1234;
  wire[1:0] T1235;
  wire[2:0] T1236;
  wire[2:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[1:0] T1241;
  wire[1:0] T1242;
  wire[1:0] T1243;
  wire[2:0] T1244;
  wire[2:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[1:0] T1249;
  wire[1:0] T1250;
  wire[1:0] T1251;
  wire[2:0] T1252;
  wire[2:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[1:0] T1257;
  wire[1:0] T1258;
  wire[1:0] T1259;
  wire[2:0] T1260;
  wire[2:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[9:0] T1268;
  wire[9:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[1:0] T1273;
  wire[1:0] T1274;
  wire[1:0] T1275;
  wire[2:0] T1276;
  wire[2:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire[1:0] T1292;
  wire[1:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[9:0] T1308;
  wire[9:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire[1:0] T1340;
  wire[1:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[9:0] T1348;
  wire[9:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire[1:0] T1356;
  wire[1:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire[1:0] T1364;
  wire[1:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire[1:0] T1372;
  wire[1:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire[1:0] T1380;
  wire[1:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[9:0] T1388;
  wire[9:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[1:0] T1396;
  wire[1:0] T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire T1401;
  wire T1402;
  wire T1403;
  wire[1:0] T1404;
  wire[1:0] T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire[1:0] T1412;
  wire[1:0] T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire[1:0] T1420;
  wire[1:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire[3:0] T1425;
  wire[3:0] T1426;
  wire[3:0] T1427;
  wire[9:0] T1428;
  wire[9:0] T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire T1435;
  wire[1:0] T1436;
  wire[1:0] T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire[1:0] T1444;
  wire[1:0] T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire[1:0] T1452;
  wire[1:0] T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[9:0] T1468;
  wire[9:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire T1473;
  wire T1474;
  wire T1475;
  wire[1:0] T1476;
  wire[1:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire[1:0] T1484;
  wire[1:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire[1:0] T1492;
  wire[1:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire T1497;
  wire T1498;
  wire T1499;
  wire[1:0] T1500;
  wire[1:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[9:0] T1508;
  wire[9:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire[1:0] T1516;
  wire[1:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire[1:0] T1524;
  wire[1:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire[1:0] T1532;
  wire[1:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[8:0] T1548;
  wire[8:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire[1:0] T1556;
  wire[1:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire[1:0] T1564;
  wire[1:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire[1:0] T1572;
  wire[1:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire T1577;
  wire T1578;
  wire T1579;
  wire[1:0] T1580;
  wire[1:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[8:0] T1588;
  wire[8:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire[1:0] T1596;
  wire[1:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire[1:0] T1604;
  wire[1:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[1:0] T1612;
  wire[1:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire[1:0] T1620;
  wire[1:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[8:0] T1628;
  wire[8:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire[1:0] T1636;
  wire[1:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire[1:0] T1644;
  wire[1:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire[1:0] T1652;
  wire[1:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire[1:0] T1660;
  wire[1:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[8:0] T1668;
  wire[8:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire[1:0] T1676;
  wire[1:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire[1:0] T1684;
  wire[1:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire T1689;
  wire T1690;
  wire T1691;
  wire[1:0] T1692;
  wire[1:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[1:0] T1700;
  wire[1:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[8:0] T1708;
  wire[8:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire[1:0] T1716;
  wire[1:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[1:0] T1724;
  wire[1:0] T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire[1:0] T1732;
  wire[1:0] T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire T1738;
  wire T1739;
  wire[1:0] T1740;
  wire[1:0] T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire[3:0] T1745;
  wire[3:0] T1746;
  wire[3:0] T1747;
  wire[8:0] T1748;
  wire[8:0] T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire T1753;
  wire T1754;
  wire T1755;
  wire[1:0] T1756;
  wire[1:0] T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire T1762;
  wire T1763;
  wire[1:0] T1764;
  wire[1:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire T1770;
  wire T1771;
  wire[1:0] T1772;
  wire[1:0] T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire T1779;
  wire[1:0] T1780;
  wire[1:0] T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire[3:0] T1785;
  wire[3:0] T1786;
  wire[3:0] T1787;
  wire[8:0] T1788;
  wire[8:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire[1:0] T1796;
  wire[1:0] T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire[1:0] T1804;
  wire[1:0] T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire[1:0] T1812;
  wire[1:0] T1813;
  wire T1814;
  wire T1815;
  wire T1816;
  wire T1817;
  wire T1818;
  wire T1819;
  wire[1:0] T1820;
  wire[1:0] T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[3:0] T1825;
  wire[3:0] T1826;
  wire[3:0] T1827;
  wire[8:0] T1828;
  wire[8:0] T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire T1834;
  wire T1835;
  wire[1:0] T1836;
  wire[1:0] T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire T1842;
  wire T1843;
  wire[1:0] T1844;
  wire[1:0] T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire T1851;
  wire[1:0] T1852;
  wire[1:0] T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire T1859;
  wire[1:0] T1860;
  wire[1:0] T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire[3:0] T1865;
  wire[3:0] T1866;
  wire[3:0] T1867;
  wire[8:0] T1868;
  wire[8:0] T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire[1:0] T1876;
  wire[1:0] T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire[1:0] T1892;
  wire[1:0] T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[1:0] T1900;
  wire[1:0] T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire[3:0] T1905;
  wire[3:0] T1906;
  wire[3:0] T1907;
  wire[8:0] T1908;
  wire[8:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire[1:0] T1916;
  wire[1:0] T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire T1921;
  wire T1922;
  wire T1923;
  wire[1:0] T1924;
  wire[1:0] T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire[1:0] T1932;
  wire[1:0] T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire T1937;
  wire T1938;
  wire T1939;
  wire[1:0] T1940;
  wire[1:0] T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire[3:0] T1945;
  wire[3:0] T1946;
  wire[3:0] T1947;
  wire[8:0] T1948;
  wire[8:0] T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire T1955;
  wire[1:0] T1956;
  wire[1:0] T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire[1:0] T1964;
  wire[1:0] T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire T1969;
  wire T1970;
  wire T1971;
  wire[1:0] T1972;
  wire[1:0] T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire[1:0] T1980;
  wire[1:0] T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire[3:0] T1985;
  wire[3:0] T1986;
  wire[3:0] T1987;
  wire[8:0] T1988;
  wire[8:0] T1989;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire[1:0] T1996;
  wire[1:0] T1997;
  wire[32:0] T1998;
  wire[32:0] T1999;
  wire[31:0] T2000;
  wire[31:0] T2001;
  wire[30:0] T2002;
  wire[30:0] T2003;
  wire[29:0] T2004;
  wire[29:0] T2005;
  wire[28:0] T2006;
  wire[28:0] T2007;
  wire[27:0] T2008;
  wire[27:0] T2009;
  wire[26:0] T2010;
  wire[26:0] T2011;
  wire[25:0] T2012;
  wire[25:0] T2013;
  wire[24:0] T2014;
  wire[24:0] T2015;
  wire[23:0] T2016;
  wire[23:0] T2017;
  wire[22:0] T2018;
  wire[22:0] T2019;
  wire[21:0] T2020;
  wire[21:0] T2021;
  wire[20:0] T2022;
  wire[20:0] T2023;
  wire[19:0] T2024;
  wire[19:0] T2025;
  wire[18:0] T2026;
  wire[18:0] T2027;
  wire[17:0] T2028;
  wire[17:0] T2029;
  wire[16:0] T2030;
  wire[16:0] T2031;
  wire[15:0] T2032;
  wire[15:0] T2033;
  wire[14:0] T2034;
  wire[14:0] T2035;
  wire[13:0] T2036;
  wire[13:0] T2037;
  wire[12:0] T2038;
  wire[12:0] T2039;
  wire[11:0] T2040;
  wire[11:0] T2041;
  wire[10:0] T2042;
  wire[10:0] T2043;
  wire[9:0] T2044;
  wire[9:0] T2045;
  wire[8:0] T2046;
  wire[8:0] T2047;
  wire[7:0] T2048;
  wire[7:0] T2049;
  wire[6:0] T2050;
  wire[6:0] T2051;
  wire[5:0] T2052;
  wire[5:0] T2053;
  wire[4:0] T2054;
  wire[4:0] T2055;
  wire[3:0] T2056;
  wire[3:0] T2057;
  wire[2:0] T2058;
  wire[2:0] T2059;
  wire[1:0] T2060;
  wire[1:0] T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire[3:0] T2065;
  wire[3:0] T2066;
  wire[3:0] T2067;
  wire[15:0] T2068;
  wire[15:0] T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire[3:0] T2073;
  wire[3:0] T2074;
  wire[3:0] T2075;
  wire[15:0] T2076;
  wire[15:0] T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[3:0] T2081;
  wire[3:0] T2082;
  wire[3:0] T2083;
  wire[15:0] T2084;
  wire[15:0] T2085;
  wire T2086;
  wire T2087;
  wire T2088;
  wire[3:0] T2089;
  wire[3:0] T2090;
  wire[3:0] T2091;
  wire[15:0] T2092;
  wire[15:0] T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire[3:0] T2097;
  wire[3:0] T2098;
  wire[3:0] T2099;
  wire[15:0] T2100;
  wire[15:0] T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire[3:0] T2105;
  wire[3:0] T2106;
  wire[3:0] T2107;
  wire[15:0] T2108;
  wire[15:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire[3:0] T2113;
  wire[3:0] T2114;
  wire[3:0] T2115;
  wire[15:0] T2116;
  wire[15:0] T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[3:0] T2121;
  wire[3:0] T2122;
  wire[3:0] T2123;
  wire[15:0] T2124;
  wire[15:0] T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire[3:0] T2129;
  wire[3:0] T2130;
  wire[3:0] T2131;
  wire[15:0] T2132;
  wire[15:0] T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire[3:0] T2137;
  wire[3:0] T2138;
  wire[3:0] T2139;
  wire[15:0] T2140;
  wire[15:0] T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire[3:0] T2145;
  wire[3:0] T2146;
  wire[3:0] T2147;
  wire[15:0] T2148;
  wire[15:0] T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire[3:0] T2153;
  wire[3:0] T2154;
  wire[3:0] T2155;
  wire[15:0] T2156;
  wire[15:0] T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire[3:0] T2161;
  wire[3:0] T2162;
  wire[3:0] T2163;
  wire[15:0] T2164;
  wire[15:0] T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire[3:0] T2169;
  wire[3:0] T2170;
  wire[3:0] T2171;
  wire[15:0] T2172;
  wire[15:0] T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  wire[3:0] T2177;
  wire[3:0] T2178;
  wire[3:0] T2179;
  wire[15:0] T2180;
  wire[15:0] T2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire[3:0] T2185;
  wire[3:0] T2186;
  wire[3:0] T2187;
  wire[15:0] T2188;
  wire[15:0] T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[3:0] T2193;
  wire[3:0] T2194;
  wire[3:0] T2195;
  wire[15:0] T2196;
  wire[15:0] T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire[3:0] T2201;
  wire[3:0] T2202;
  wire[3:0] T2203;
  wire[15:0] T2204;
  wire[15:0] T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire[3:0] T2209;
  wire[3:0] T2210;
  wire[3:0] T2211;
  wire[15:0] T2212;
  wire[15:0] T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire[3:0] T2217;
  wire[3:0] T2218;
  wire[3:0] T2219;
  wire[15:0] T2220;
  wire[15:0] T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire[3:0] T2225;
  wire[3:0] T2226;
  wire[3:0] T2227;
  wire[15:0] T2228;
  wire[15:0] T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire[3:0] T2233;
  wire[3:0] T2234;
  wire[3:0] T2235;
  wire[15:0] T2236;
  wire[15:0] T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire[3:0] T2241;
  wire[3:0] T2242;
  wire[3:0] T2243;
  wire[15:0] T2244;
  wire[15:0] T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  wire[3:0] T2249;
  wire[3:0] T2250;
  wire[3:0] T2251;
  wire[15:0] T2252;
  wire[15:0] T2253;
  wire T2254;
  wire T2255;
  wire T2256;
  wire[3:0] T2257;
  wire[3:0] T2258;
  wire[3:0] T2259;
  wire[15:0] T2260;
  wire[15:0] T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[3:0] T2265;
  wire[3:0] T2266;
  wire[3:0] T2267;
  wire[15:0] T2268;
  wire[15:0] T2269;
  wire T2270;
  wire T2271;
  wire T2272;
  wire[3:0] T2273;
  wire[3:0] T2274;
  wire[3:0] T2275;
  wire[15:0] T2276;
  wire[15:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire[3:0] T2281;
  wire[3:0] T2282;
  wire[3:0] T2283;
  wire[15:0] T2284;
  wire[15:0] T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire[3:0] T2289;
  wire[3:0] T2290;
  wire[3:0] T2291;
  wire[15:0] T2292;
  wire[15:0] T2293;
  wire T2294;
  wire T2295;
  wire T2296;
  wire[3:0] T2297;
  wire[3:0] T2298;
  wire[3:0] T2299;
  wire[15:0] T2300;
  wire[15:0] T2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire[3:0] T2305;
  wire[3:0] T2306;
  wire[3:0] T2307;
  wire[15:0] T2308;
  wire[15:0] T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire[3:0] T2313;
  wire[3:0] T2314;
  wire[3:0] T2315;
  wire[15:0] T2316;
  wire[15:0] T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  wire[3:0] T2321;
  wire[3:0] T2322;
  wire[3:0] T2323;
  wire[15:0] T2324;
  wire[15:0] T2325;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1990, T2};
  assign T2 = T3;
  assign T3 = {T1982, T4};
  assign T4 = T5;
  assign T5 = {T1974, T6};
  assign T6 = T7;
  assign T7 = {T1966, T8};
  assign T8 = T9;
  assign T9 = {T1958, T10};
  assign T10 = T11;
  assign T11 = {T1950, T12};
  assign T12 = T13;
  assign T13 = {T1942, T14};
  assign T14 = T15;
  assign T15 = {T1934, T16};
  assign T16 = T17;
  assign T17 = {T1926, T18};
  assign T18 = T19;
  assign T19 = {T1918, T20};
  assign T20 = T21;
  assign T21 = {T1910, T22};
  assign T22 = T23;
  assign T23 = {T1902, T24};
  assign T24 = T25;
  assign T25 = {T1894, T26};
  assign T26 = T27;
  assign T27 = {T1886, T28};
  assign T28 = T29;
  assign T29 = {T1878, T30};
  assign T30 = T31;
  assign T31 = {T1870, T32};
  assign T32 = T33;
  assign T33 = {T1862, T34};
  assign T34 = T35;
  assign T35 = {T1854, T36};
  assign T36 = T37;
  assign T37 = {T1846, T38};
  assign T38 = T39;
  assign T39 = {T1838, T40};
  assign T40 = T41;
  assign T41 = {T1830, T42};
  assign T42 = T43;
  assign T43 = {T1822, T44};
  assign T44 = T45;
  assign T45 = {T1814, T46};
  assign T46 = T47;
  assign T47 = {T1806, T48};
  assign T48 = T49;
  assign T49 = {T1798, T50};
  assign T50 = T51;
  assign T51 = {T1790, T52};
  assign T52 = T53;
  assign T53 = {T1782, T54};
  assign T54 = T55;
  assign T55 = {T1774, T56};
  assign T56 = T57;
  assign T57 = {T1766, T58};
  assign T58 = T59;
  assign T59 = {T1758, T60};
  assign T60 = T61;
  assign T61 = {T1750, T62};
  assign T62 = T63;
  assign T63 = {T1742, T64};
  assign T64 = T65;
  assign T65 = {T1734, T66};
  assign T66 = T67;
  assign T67 = {T1726, T68};
  assign T68 = T69;
  assign T69 = {T1718, T70};
  assign T70 = T71;
  assign T71 = {T1710, T72};
  assign T72 = T73;
  assign T73 = {T1702, T74};
  assign T74 = T75;
  assign T75 = {T1694, T76};
  assign T76 = T77;
  assign T77 = {T1686, T78};
  assign T78 = T79;
  assign T79 = {T1678, T80};
  assign T80 = T81;
  assign T81 = {T1670, T82};
  assign T82 = T83;
  assign T83 = {T1662, T84};
  assign T84 = T85;
  assign T85 = {T1654, T86};
  assign T86 = T87;
  assign T87 = {T1646, T88};
  assign T88 = T89;
  assign T89 = {T1638, T90};
  assign T90 = T91;
  assign T91 = {T1630, T92};
  assign T92 = T93;
  assign T93 = {T1622, T94};
  assign T94 = T95;
  assign T95 = {T1614, T96};
  assign T96 = T97;
  assign T97 = {T1606, T98};
  assign T98 = T99;
  assign T99 = {T1598, T100};
  assign T100 = T101;
  assign T101 = {T1590, T102};
  assign T102 = T103;
  assign T103 = {T1582, T104};
  assign T104 = T105;
  assign T105 = {T1574, T106};
  assign T106 = T107;
  assign T107 = {T1566, T108};
  assign T108 = T109;
  assign T109 = {T1558, T110};
  assign T110 = T111;
  assign T111 = {T1550, T112};
  assign T112 = T113;
  assign T113 = {T1542, T114};
  assign T114 = T115;
  assign T115 = {T1534, T116};
  assign T116 = T117;
  assign T117 = {T1526, T118};
  assign T118 = T119;
  assign T119 = {T1518, T120};
  assign T120 = T121;
  assign T121 = {T1510, T122};
  assign T122 = T123;
  assign T123 = {T1502, T124};
  assign T124 = T125;
  assign T125 = {T1494, T126};
  assign T126 = T127;
  assign T127 = {T1486, T128};
  assign T128 = T129;
  assign T129 = {T1478, T130};
  assign T130 = T131;
  assign T131 = {T1470, T132};
  assign T132 = T133;
  assign T133 = {T1462, T134};
  assign T134 = T135;
  assign T135 = {T1454, T136};
  assign T136 = T137;
  assign T137 = {T1446, T138};
  assign T138 = T139;
  assign T139 = {T1438, T140};
  assign T140 = T141;
  assign T141 = {T1430, T142};
  assign T142 = T143;
  assign T143 = {T1422, T144};
  assign T144 = T145;
  assign T145 = {T1414, T146};
  assign T146 = T147;
  assign T147 = {T1406, T148};
  assign T148 = T149;
  assign T149 = {T1398, T150};
  assign T150 = T151;
  assign T151 = {T1390, T152};
  assign T152 = T153;
  assign T153 = {T1382, T154};
  assign T154 = T155;
  assign T155 = {T1374, T156};
  assign T156 = T157;
  assign T157 = {T1366, T158};
  assign T158 = T159;
  assign T159 = {T1358, T160};
  assign T160 = T161;
  assign T161 = {T1350, T162};
  assign T162 = T163;
  assign T163 = {T1342, T164};
  assign T164 = T165;
  assign T165 = {T1334, T166};
  assign T166 = T167;
  assign T167 = {T1326, T168};
  assign T168 = T169;
  assign T169 = {T1318, T170};
  assign T170 = T171;
  assign T171 = {T1310, T172};
  assign T172 = T173;
  assign T173 = {T1302, T174};
  assign T174 = T175;
  assign T175 = {T1294, T176};
  assign T176 = T177;
  assign T177 = {T1286, T178};
  assign T178 = T179;
  assign T179 = {T1278, T180};
  assign T180 = T181;
  assign T181 = {T1270, T182};
  assign T182 = T183;
  assign T183 = {T1262, T184};
  assign T184 = T185;
  assign T185 = {T1254, T186};
  assign T186 = T187;
  assign T187 = {T1246, T188};
  assign T188 = T189;
  assign T189 = {T1238, T190};
  assign T190 = T191;
  assign T191 = {T1230, T192};
  assign T192 = T193;
  assign T193 = {T1222, T194};
  assign T194 = T195;
  assign T195 = {T1214, T196};
  assign T196 = T197;
  assign T197 = {T1206, T198};
  assign T198 = T199;
  assign T199 = {T1198, T200};
  assign T200 = T201;
  assign T201 = {T1190, T202};
  assign T202 = T203;
  assign T203 = {T1182, T204};
  assign T204 = T205;
  assign T205 = {T1174, T206};
  assign T206 = T207;
  assign T207 = {T1166, T208};
  assign T208 = T209;
  assign T209 = {T1158, T210};
  assign T210 = T211;
  assign T211 = {T1150, T212};
  assign T212 = T213;
  assign T213 = {T1142, T214};
  assign T214 = T215;
  assign T215 = {T1134, T216};
  assign T216 = T217;
  assign T217 = {T1126, T218};
  assign T218 = T219;
  assign T219 = {T1118, T220};
  assign T220 = T221;
  assign T221 = {T1110, T222};
  assign T222 = T223;
  assign T223 = {T1102, T224};
  assign T224 = T225;
  assign T225 = {T1094, T226};
  assign T226 = T227;
  assign T227 = {T1086, T228};
  assign T228 = T229;
  assign T229 = {T1078, T230};
  assign T230 = T231;
  assign T231 = {T1070, T232};
  assign T232 = T233;
  assign T233 = {T1062, T234};
  assign T234 = T235;
  assign T235 = {T1054, T236};
  assign T236 = T237;
  assign T237 = {T1046, T238};
  assign T238 = T239;
  assign T239 = {T1038, T240};
  assign T240 = T241;
  assign T241 = {T1030, T242};
  assign T242 = T243;
  assign T243 = {T1022, T244};
  assign T244 = T245;
  assign T245 = {T1014, T246};
  assign T246 = T247;
  assign T247 = {T1006, T248};
  assign T248 = T249;
  assign T249 = {T998, T250};
  assign T250 = T251;
  assign T251 = {T990, T252};
  assign T252 = T253;
  assign T253 = {T982, T254};
  assign T254 = T255;
  assign T255 = {T974, T256};
  assign T256 = T257;
  assign T257 = {T966, T258};
  assign T258 = T259;
  assign T259 = {T958, T260};
  assign T260 = T261;
  assign T261 = {T950, T262};
  assign T262 = T263;
  assign T263 = {T942, T264};
  assign T264 = T265;
  assign T265 = {T934, T266};
  assign T266 = T267;
  assign T267 = {T926, T268};
  assign T268 = T269;
  assign T269 = {T918, T270};
  assign T270 = T271;
  assign T271 = {T910, T272};
  assign T272 = T273;
  assign T273 = {T902, T274};
  assign T274 = T275;
  assign T275 = {T894, T276};
  assign T276 = T277;
  assign T277 = {T886, T278};
  assign T278 = T279;
  assign T279 = {T878, T280};
  assign T280 = T281;
  assign T281 = {T870, T282};
  assign T282 = T283;
  assign T283 = {T862, T284};
  assign T284 = T285;
  assign T285 = {T854, T286};
  assign T286 = T287;
  assign T287 = {T846, T288};
  assign T288 = T289;
  assign T289 = {T838, T290};
  assign T290 = T291;
  assign T291 = {T830, T292};
  assign T292 = T293;
  assign T293 = {T822, T294};
  assign T294 = T295;
  assign T295 = {T814, T296};
  assign T296 = T297;
  assign T297 = {T806, T298};
  assign T298 = T299;
  assign T299 = {T798, T300};
  assign T300 = T301;
  assign T301 = {T790, T302};
  assign T302 = T303;
  assign T303 = {T782, T304};
  assign T304 = T305;
  assign T305 = {T774, T306};
  assign T306 = T307;
  assign T307 = {T766, T308};
  assign T308 = T309;
  assign T309 = {T758, T310};
  assign T310 = T311;
  assign T311 = {T750, T312};
  assign T312 = T313;
  assign T313 = {T742, T314};
  assign T314 = T315;
  assign T315 = {T734, T316};
  assign T316 = T317;
  assign T317 = {T726, T318};
  assign T318 = T319;
  assign T319 = {T718, T320};
  assign T320 = T321;
  assign T321 = {T710, T322};
  assign T322 = T323;
  assign T323 = {T702, T324};
  assign T324 = T325;
  assign T325 = {T694, T326};
  assign T326 = T327;
  assign T327 = {T686, T328};
  assign T328 = T329;
  assign T329 = {T678, T330};
  assign T330 = T331;
  assign T331 = {T670, T332};
  assign T332 = T333;
  assign T333 = {T662, T334};
  assign T334 = T335;
  assign T335 = {T654, T336};
  assign T336 = T337;
  assign T337 = {T646, T338};
  assign T338 = T339;
  assign T339 = {T638, T340};
  assign T340 = T341;
  assign T341 = {T630, T342};
  assign T342 = T343;
  assign T343 = {T622, T344};
  assign T344 = T345;
  assign T345 = {T614, T346};
  assign T346 = T347;
  assign T347 = {T606, T348};
  assign T348 = T349;
  assign T349 = {T598, T350};
  assign T350 = T351;
  assign T351 = {T590, T352};
  assign T352 = T353;
  assign T353 = {T582, T354};
  assign T354 = T355;
  assign T355 = {T574, T356};
  assign T356 = T357;
  assign T357 = {T566, T358};
  assign T358 = T359;
  assign T359 = {T558, T360};
  assign T360 = T361;
  assign T361 = {T550, T362};
  assign T362 = T363;
  assign T363 = {T542, T364};
  assign T364 = T365;
  assign T365 = {T534, T366};
  assign T366 = T367;
  assign T367 = {T526, T368};
  assign T368 = T369;
  assign T369 = {T518, T370};
  assign T370 = T371;
  assign T371 = {T510, T372};
  assign T372 = T373;
  assign T373 = {T502, T374};
  assign T374 = T375;
  assign T375 = {T494, T376};
  assign T376 = T377;
  assign T377 = {T486, T378};
  assign T378 = T379;
  assign T379 = {T478, T380};
  assign T380 = T381;
  assign T381 = {T470, T382};
  assign T382 = T383;
  assign T383 = {T462, T384};
  assign T384 = T385;
  assign T385 = {T454, T386};
  assign T386 = T387;
  assign T387 = {T446, T388};
  assign T388 = T389;
  assign T389 = {T438, T390};
  assign T390 = T391;
  assign T391 = {T430, T392};
  assign T392 = T393;
  assign T393 = {T422, T394};
  assign T394 = T395;
  assign T395 = {T414, T396};
  assign T396 = T397;
  assign T397 = {T406, T398};
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[4'he/* 14*/:4'hc/* 12*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[5'h11/* 17*/:4'hf/* 15*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[5'h14/* 20*/:5'h12/* 18*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[5'h17/* 23*/:5'h15/* 21*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[5'h1a/* 26*/:5'h18/* 24*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[5'h1d/* 29*/:5'h1b/* 27*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[6'h34/* 52*/:6'h32/* 50*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[6'h37/* 55*/:6'h35/* 53*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[6'h3a/* 58*/:6'h38/* 56*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[6'h3d/* 61*/:6'h3b/* 59*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h40/* 64*/:6'h3e/* 62*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h43/* 67*/:7'h41/* 65*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h46/* 70*/:7'h44/* 68*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h49/* 73*/:7'h47/* 71*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[7'h4c/* 76*/:7'h4a/* 74*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[7'h4f/* 79*/:7'h4d/* 77*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[6'h34/* 52*/:6'h34/* 52*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h55/* 85*/:7'h54/* 84*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[6'h35/* 53*/:6'h35/* 53*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h57/* 87*/:7'h56/* 86*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[7'h59/* 89*/:7'h58/* 88*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[7'h66/* 102*/:7'h64/* 100*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[7'h69/* 105*/:7'h67/* 103*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[7'h6c/* 108*/:7'h6a/* 106*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[7'h7e/* 126*/:7'h7c/* 124*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'h81/* 129*/:7'h7f/* 127*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'h83/* 131*/:8'h82/* 130*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'h85/* 133*/:8'h84/* 132*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'h87/* 135*/:8'h86/* 134*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h53/* 83*/:7'h53/* 83*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h54/* 84*/:7'h54/* 84*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[7'h55/* 85*/:7'h55/* 85*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[8'h91/* 145*/:8'h90/* 144*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[8'h93/* 147*/:8'h92/* 146*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[8'h95/* 149*/:8'h94/* 148*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[8'ha0/* 160*/:8'h96/* 150*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[8'hae/* 174*/:8'ha4/* 164*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[7'h65/* 101*/:7'h64/* 100*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[8'hb1/* 177*/:8'haf/* 175*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[7'h69/* 105*/:7'h66/* 102*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[8'hbc/* 188*/:8'hb2/* 178*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[8'hbf/* 191*/:8'hbd/* 189*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[7'h71/* 113*/:7'h70/* 112*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[8'hcd/* 205*/:8'hcb/* 203*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[8'hd8/* 216*/:8'hce/* 206*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[7'h77/* 119*/:7'h76/* 118*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[8'hdb/* 219*/:8'hd9/* 217*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[8'he6/* 230*/:8'hdc/* 220*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[8'he9/* 233*/:8'he7/* 231*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'h81/* 129*/:7'h7e/* 126*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[8'hf4/* 244*/:8'hea/* 234*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[8'hf7/* 247*/:8'hf5/* 245*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h102/* 258*/:8'hf8/* 248*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'h89/* 137*/:8'h88/* 136*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h105/* 261*/:9'h103/* 259*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h110/* 272*/:9'h106/* 262*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h113/* 275*/:9'h111/* 273*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h11e/* 286*/:9'h114/* 276*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'h95/* 149*/:8'h94/* 148*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h121/* 289*/:9'h11f/* 287*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h12c/* 300*/:9'h122/* 290*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h13b/* 315*/:9'h13a/* 314*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h146/* 326*/:9'h13c/* 316*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'ha4/* 164*/:8'ha4/* 164*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'ha8/* 168*/:8'ha5/* 165*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h153/* 339*/:9'h149/* 329*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h155/* 341*/:9'h154/* 340*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'had/* 173*/:8'haa/* 170*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h160/* 352*/:9'h156/* 342*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h162/* 354*/:9'h161/* 353*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hb2/* 178*/:8'haf/* 175*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h16d/* 365*/:9'h163/* 355*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h16f/* 367*/:9'h16e/* 366*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h17a/* 378*/:9'h170/* 368*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[9'h17c/* 380*/:9'h17b/* 379*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hbc/* 188*/:8'hb9/* 185*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[9'h187/* 391*/:9'h17d/* 381*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[9'h189/* 393*/:9'h188/* 392*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hc1/* 193*/:8'hbe/* 190*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[9'h194/* 404*/:9'h18a/* 394*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[9'h196/* 406*/:9'h195/* 405*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[9'h1a6/* 422*/:9'h1a4/* 420*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[9'h1a9/* 425*/:9'h1a7/* 423*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[9'h1ac/* 428*/:9'h1aa/* 426*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[8'hd1/* 209*/:8'hce/* 206*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[9'h1b6/* 438*/:9'h1ad/* 429*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[9'h1b9/* 441*/:9'h1b7/* 439*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[8'hd5/* 213*/:8'hd4/* 212*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[9'h1bc/* 444*/:9'h1ba/* 442*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[8'hd7/* 215*/:8'hd6/* 214*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[9'h1bf/* 447*/:9'h1bd/* 445*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[9'h1c2/* 450*/:9'h1c0/* 448*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[8'hdd/* 221*/:8'hda/* 218*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[9'h1cc/* 460*/:9'h1c3/* 451*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[9'h1cf/* 463*/:9'h1cd/* 461*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[9'h1d1/* 465*/:9'h1d0/* 464*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[9'h1d3/* 467*/:9'h1d2/* 466*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[8'he2/* 226*/:8'he2/* 226*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[9'h1d5/* 469*/:9'h1d4/* 468*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[8'he6/* 230*/:8'he3/* 227*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[9'h1df/* 479*/:9'h1d6/* 470*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[8'he7/* 231*/:8'he7/* 231*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[9'h1e1/* 481*/:9'h1e0/* 480*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[8'he8/* 232*/:8'he8/* 232*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[9'h1e3/* 483*/:9'h1e2/* 482*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[8'he9/* 233*/:8'he9/* 233*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[9'h1e5/* 485*/:9'h1e4/* 484*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[8'hea/* 234*/:8'hea/* 234*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[9'h1e7/* 487*/:9'h1e6/* 486*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[8'hee/* 238*/:8'heb/* 235*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[9'h1f1/* 497*/:9'h1e8/* 488*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[8'hef/* 239*/:8'hef/* 239*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[9'h1f3/* 499*/:9'h1f2/* 498*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[9'h1f5/* 501*/:9'h1f4/* 500*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[9'h1f7/* 503*/:9'h1f6/* 502*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[9'h1f9/* 505*/:9'h1f8/* 504*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[8'hf6/* 246*/:8'hf3/* 243*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h203/* 515*/:9'h1fa/* 506*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h205/* 517*/:10'h204/* 516*/];
  assign T1398 = T1399;
  assign T1399 = T1400;
  assign T1400 = T1404[T1401];
  assign T1401 = T1402;
  assign T1402 = T1403;
  assign T1403 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1404 = T1405;
  assign T1405 = io_chanxy_in[10'h207/* 519*/:10'h206/* 518*/];
  assign T1406 = T1407;
  assign T1407 = T1408;
  assign T1408 = T1412[T1409];
  assign T1409 = T1410;
  assign T1410 = T1411;
  assign T1411 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T1412 = T1413;
  assign T1413 = io_chanxy_in[10'h209/* 521*/:10'h208/* 520*/];
  assign T1414 = T1415;
  assign T1415 = T1416;
  assign T1416 = T1420[T1417];
  assign T1417 = T1418;
  assign T1418 = T1419;
  assign T1419 = io_chanxy_config[8'hfa/* 250*/:8'hfa/* 250*/];
  assign T1420 = T1421;
  assign T1421 = io_chanxy_in[10'h20b/* 523*/:10'h20a/* 522*/];
  assign T1422 = T1423;
  assign T1423 = T1424;
  assign T1424 = T1428[T1425];
  assign T1425 = T1426;
  assign T1426 = T1427;
  assign T1427 = io_chanxy_config[8'hfe/* 254*/:8'hfb/* 251*/];
  assign T1428 = T1429;
  assign T1429 = io_chanxy_in[10'h215/* 533*/:10'h20c/* 524*/];
  assign T1430 = T1431;
  assign T1431 = T1432;
  assign T1432 = T1436[T1433];
  assign T1433 = T1434;
  assign T1434 = T1435;
  assign T1435 = io_chanxy_config[8'hff/* 255*/:8'hff/* 255*/];
  assign T1436 = T1437;
  assign T1437 = io_chanxy_in[10'h217/* 535*/:10'h216/* 534*/];
  assign T1438 = T1439;
  assign T1439 = T1440;
  assign T1440 = T1444[T1441];
  assign T1441 = T1442;
  assign T1442 = T1443;
  assign T1443 = io_chanxy_config[9'h100/* 256*/:9'h100/* 256*/];
  assign T1444 = T1445;
  assign T1445 = io_chanxy_in[10'h219/* 537*/:10'h218/* 536*/];
  assign T1446 = T1447;
  assign T1447 = T1448;
  assign T1448 = T1452[T1449];
  assign T1449 = T1450;
  assign T1450 = T1451;
  assign T1451 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1452 = T1453;
  assign T1453 = io_chanxy_in[10'h21b/* 539*/:10'h21a/* 538*/];
  assign T1454 = T1455;
  assign T1455 = T1456;
  assign T1456 = T1460[T1457];
  assign T1457 = T1458;
  assign T1458 = T1459;
  assign T1459 = io_chanxy_config[9'h102/* 258*/:9'h102/* 258*/];
  assign T1460 = T1461;
  assign T1461 = io_chanxy_in[10'h21d/* 541*/:10'h21c/* 540*/];
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_chanxy_config[9'h106/* 262*/:9'h103/* 259*/];
  assign T1468 = T1469;
  assign T1469 = io_chanxy_in[10'h227/* 551*/:10'h21e/* 542*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_chanxy_config[9'h107/* 263*/:9'h107/* 263*/];
  assign T1476 = T1477;
  assign T1477 = io_chanxy_in[10'h229/* 553*/:10'h228/* 552*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_chanxy_config[9'h108/* 264*/:9'h108/* 264*/];
  assign T1484 = T1485;
  assign T1485 = io_chanxy_in[10'h22b/* 555*/:10'h22a/* 554*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_chanxy_config[9'h109/* 265*/:9'h109/* 265*/];
  assign T1492 = T1493;
  assign T1493 = io_chanxy_in[10'h22d/* 557*/:10'h22c/* 556*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_chanxy_config[9'h10a/* 266*/:9'h10a/* 266*/];
  assign T1500 = T1501;
  assign T1501 = io_chanxy_in[10'h22f/* 559*/:10'h22e/* 558*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_chanxy_config[9'h10e/* 270*/:9'h10b/* 267*/];
  assign T1508 = T1509;
  assign T1509 = io_chanxy_in[10'h239/* 569*/:10'h230/* 560*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_chanxy_config[9'h10f/* 271*/:9'h10f/* 271*/];
  assign T1516 = T1517;
  assign T1517 = io_chanxy_in[10'h23b/* 571*/:10'h23a/* 570*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_chanxy_config[9'h110/* 272*/:9'h110/* 272*/];
  assign T1524 = T1525;
  assign T1525 = io_chanxy_in[10'h23d/* 573*/:10'h23c/* 572*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_chanxy_config[9'h111/* 273*/:9'h111/* 273*/];
  assign T1532 = T1533;
  assign T1533 = io_chanxy_in[10'h23f/* 575*/:10'h23e/* 574*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_chanxy_config[9'h112/* 274*/:9'h112/* 274*/];
  assign T1540 = T1541;
  assign T1541 = io_chanxy_in[10'h241/* 577*/:10'h240/* 576*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_chanxy_config[9'h116/* 278*/:9'h113/* 275*/];
  assign T1548 = T1549;
  assign T1549 = io_chanxy_in[10'h24a/* 586*/:10'h242/* 578*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_chanxy_config[9'h117/* 279*/:9'h117/* 279*/];
  assign T1556 = T1557;
  assign T1557 = io_chanxy_in[10'h24c/* 588*/:10'h24b/* 587*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_chanxy_config[9'h118/* 280*/:9'h118/* 280*/];
  assign T1564 = T1565;
  assign T1565 = io_chanxy_in[10'h24e/* 590*/:10'h24d/* 589*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_chanxy_config[9'h119/* 281*/:9'h119/* 281*/];
  assign T1572 = T1573;
  assign T1573 = io_chanxy_in[10'h250/* 592*/:10'h24f/* 591*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_chanxy_config[9'h11a/* 282*/:9'h11a/* 282*/];
  assign T1580 = T1581;
  assign T1581 = io_chanxy_in[10'h252/* 594*/:10'h251/* 593*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_chanxy_config[9'h11e/* 286*/:9'h11b/* 283*/];
  assign T1588 = T1589;
  assign T1589 = io_chanxy_in[10'h25b/* 603*/:10'h253/* 595*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_chanxy_config[9'h11f/* 287*/:9'h11f/* 287*/];
  assign T1596 = T1597;
  assign T1597 = io_chanxy_in[10'h25d/* 605*/:10'h25c/* 604*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_chanxy_config[9'h120/* 288*/:9'h120/* 288*/];
  assign T1604 = T1605;
  assign T1605 = io_chanxy_in[10'h25f/* 607*/:10'h25e/* 606*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_chanxy_config[9'h121/* 289*/:9'h121/* 289*/];
  assign T1612 = T1613;
  assign T1613 = io_chanxy_in[10'h261/* 609*/:10'h260/* 608*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_chanxy_config[9'h122/* 290*/:9'h122/* 290*/];
  assign T1620 = T1621;
  assign T1621 = io_chanxy_in[10'h263/* 611*/:10'h262/* 610*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_chanxy_config[9'h126/* 294*/:9'h123/* 291*/];
  assign T1628 = T1629;
  assign T1629 = io_chanxy_in[10'h26c/* 620*/:10'h264/* 612*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_chanxy_config[9'h127/* 295*/:9'h127/* 295*/];
  assign T1636 = T1637;
  assign T1637 = io_chanxy_in[10'h26e/* 622*/:10'h26d/* 621*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_chanxy_config[9'h128/* 296*/:9'h128/* 296*/];
  assign T1644 = T1645;
  assign T1645 = io_chanxy_in[10'h270/* 624*/:10'h26f/* 623*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_chanxy_config[9'h129/* 297*/:9'h129/* 297*/];
  assign T1652 = T1653;
  assign T1653 = io_chanxy_in[10'h272/* 626*/:10'h271/* 625*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_chanxy_config[9'h12a/* 298*/:9'h12a/* 298*/];
  assign T1660 = T1661;
  assign T1661 = io_chanxy_in[10'h274/* 628*/:10'h273/* 627*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_chanxy_config[9'h12e/* 302*/:9'h12b/* 299*/];
  assign T1668 = T1669;
  assign T1669 = io_chanxy_in[10'h27d/* 637*/:10'h275/* 629*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_chanxy_config[9'h12f/* 303*/:9'h12f/* 303*/];
  assign T1676 = T1677;
  assign T1677 = io_chanxy_in[10'h27f/* 639*/:10'h27e/* 638*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_chanxy_config[9'h130/* 304*/:9'h130/* 304*/];
  assign T1684 = T1685;
  assign T1685 = io_chanxy_in[10'h281/* 641*/:10'h280/* 640*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_chanxy_config[9'h131/* 305*/:9'h131/* 305*/];
  assign T1692 = T1693;
  assign T1693 = io_chanxy_in[10'h283/* 643*/:10'h282/* 642*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_chanxy_config[9'h132/* 306*/:9'h132/* 306*/];
  assign T1700 = T1701;
  assign T1701 = io_chanxy_in[10'h285/* 645*/:10'h284/* 644*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_chanxy_config[9'h136/* 310*/:9'h133/* 307*/];
  assign T1708 = T1709;
  assign T1709 = io_chanxy_in[10'h28e/* 654*/:10'h286/* 646*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_chanxy_config[9'h137/* 311*/:9'h137/* 311*/];
  assign T1716 = T1717;
  assign T1717 = io_chanxy_in[10'h290/* 656*/:10'h28f/* 655*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_chanxy_config[9'h138/* 312*/:9'h138/* 312*/];
  assign T1724 = T1725;
  assign T1725 = io_chanxy_in[10'h292/* 658*/:10'h291/* 657*/];
  assign T1726 = T1727;
  assign T1727 = T1728;
  assign T1728 = T1732[T1729];
  assign T1729 = T1730;
  assign T1730 = T1731;
  assign T1731 = io_chanxy_config[9'h139/* 313*/:9'h139/* 313*/];
  assign T1732 = T1733;
  assign T1733 = io_chanxy_in[10'h294/* 660*/:10'h293/* 659*/];
  assign T1734 = T1735;
  assign T1735 = T1736;
  assign T1736 = T1740[T1737];
  assign T1737 = T1738;
  assign T1738 = T1739;
  assign T1739 = io_chanxy_config[9'h13a/* 314*/:9'h13a/* 314*/];
  assign T1740 = T1741;
  assign T1741 = io_chanxy_in[10'h296/* 662*/:10'h295/* 661*/];
  assign T1742 = T1743;
  assign T1743 = T1744;
  assign T1744 = T1748[T1745];
  assign T1745 = T1746;
  assign T1746 = T1747;
  assign T1747 = io_chanxy_config[9'h13e/* 318*/:9'h13b/* 315*/];
  assign T1748 = T1749;
  assign T1749 = io_chanxy_in[10'h29f/* 671*/:10'h297/* 663*/];
  assign T1750 = T1751;
  assign T1751 = T1752;
  assign T1752 = T1756[T1753];
  assign T1753 = T1754;
  assign T1754 = T1755;
  assign T1755 = io_chanxy_config[9'h13f/* 319*/:9'h13f/* 319*/];
  assign T1756 = T1757;
  assign T1757 = io_chanxy_in[10'h2a1/* 673*/:10'h2a0/* 672*/];
  assign T1758 = T1759;
  assign T1759 = T1760;
  assign T1760 = T1764[T1761];
  assign T1761 = T1762;
  assign T1762 = T1763;
  assign T1763 = io_chanxy_config[9'h140/* 320*/:9'h140/* 320*/];
  assign T1764 = T1765;
  assign T1765 = io_chanxy_in[10'h2a3/* 675*/:10'h2a2/* 674*/];
  assign T1766 = T1767;
  assign T1767 = T1768;
  assign T1768 = T1772[T1769];
  assign T1769 = T1770;
  assign T1770 = T1771;
  assign T1771 = io_chanxy_config[9'h141/* 321*/:9'h141/* 321*/];
  assign T1772 = T1773;
  assign T1773 = io_chanxy_in[10'h2a5/* 677*/:10'h2a4/* 676*/];
  assign T1774 = T1775;
  assign T1775 = T1776;
  assign T1776 = T1780[T1777];
  assign T1777 = T1778;
  assign T1778 = T1779;
  assign T1779 = io_chanxy_config[9'h142/* 322*/:9'h142/* 322*/];
  assign T1780 = T1781;
  assign T1781 = io_chanxy_in[10'h2a7/* 679*/:10'h2a6/* 678*/];
  assign T1782 = T1783;
  assign T1783 = T1784;
  assign T1784 = T1788[T1785];
  assign T1785 = T1786;
  assign T1786 = T1787;
  assign T1787 = io_chanxy_config[9'h146/* 326*/:9'h143/* 323*/];
  assign T1788 = T1789;
  assign T1789 = io_chanxy_in[10'h2b0/* 688*/:10'h2a8/* 680*/];
  assign T1790 = T1791;
  assign T1791 = T1792;
  assign T1792 = T1796[T1793];
  assign T1793 = T1794;
  assign T1794 = T1795;
  assign T1795 = io_chanxy_config[9'h147/* 327*/:9'h147/* 327*/];
  assign T1796 = T1797;
  assign T1797 = io_chanxy_in[10'h2b2/* 690*/:10'h2b1/* 689*/];
  assign T1798 = T1799;
  assign T1799 = T1800;
  assign T1800 = T1804[T1801];
  assign T1801 = T1802;
  assign T1802 = T1803;
  assign T1803 = io_chanxy_config[9'h148/* 328*/:9'h148/* 328*/];
  assign T1804 = T1805;
  assign T1805 = io_chanxy_in[10'h2b4/* 692*/:10'h2b3/* 691*/];
  assign T1806 = T1807;
  assign T1807 = T1808;
  assign T1808 = T1812[T1809];
  assign T1809 = T1810;
  assign T1810 = T1811;
  assign T1811 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1812 = T1813;
  assign T1813 = io_chanxy_in[10'h2b6/* 694*/:10'h2b5/* 693*/];
  assign T1814 = T1815;
  assign T1815 = T1816;
  assign T1816 = T1820[T1817];
  assign T1817 = T1818;
  assign T1818 = T1819;
  assign T1819 = io_chanxy_config[9'h14a/* 330*/:9'h14a/* 330*/];
  assign T1820 = T1821;
  assign T1821 = io_chanxy_in[10'h2b8/* 696*/:10'h2b7/* 695*/];
  assign T1822 = T1823;
  assign T1823 = T1824;
  assign T1824 = T1828[T1825];
  assign T1825 = T1826;
  assign T1826 = T1827;
  assign T1827 = io_chanxy_config[9'h14e/* 334*/:9'h14b/* 331*/];
  assign T1828 = T1829;
  assign T1829 = io_chanxy_in[10'h2c1/* 705*/:10'h2b9/* 697*/];
  assign T1830 = T1831;
  assign T1831 = T1832;
  assign T1832 = T1836[T1833];
  assign T1833 = T1834;
  assign T1834 = T1835;
  assign T1835 = io_chanxy_config[9'h14f/* 335*/:9'h14f/* 335*/];
  assign T1836 = T1837;
  assign T1837 = io_chanxy_in[10'h2c3/* 707*/:10'h2c2/* 706*/];
  assign T1838 = T1839;
  assign T1839 = T1840;
  assign T1840 = T1844[T1841];
  assign T1841 = T1842;
  assign T1842 = T1843;
  assign T1843 = io_chanxy_config[9'h150/* 336*/:9'h150/* 336*/];
  assign T1844 = T1845;
  assign T1845 = io_chanxy_in[10'h2c5/* 709*/:10'h2c4/* 708*/];
  assign T1846 = T1847;
  assign T1847 = T1848;
  assign T1848 = T1852[T1849];
  assign T1849 = T1850;
  assign T1850 = T1851;
  assign T1851 = io_chanxy_config[9'h151/* 337*/:9'h151/* 337*/];
  assign T1852 = T1853;
  assign T1853 = io_chanxy_in[10'h2c7/* 711*/:10'h2c6/* 710*/];
  assign T1854 = T1855;
  assign T1855 = T1856;
  assign T1856 = T1860[T1857];
  assign T1857 = T1858;
  assign T1858 = T1859;
  assign T1859 = io_chanxy_config[9'h152/* 338*/:9'h152/* 338*/];
  assign T1860 = T1861;
  assign T1861 = io_chanxy_in[10'h2c9/* 713*/:10'h2c8/* 712*/];
  assign T1862 = T1863;
  assign T1863 = T1864;
  assign T1864 = T1868[T1865];
  assign T1865 = T1866;
  assign T1866 = T1867;
  assign T1867 = io_chanxy_config[9'h156/* 342*/:9'h153/* 339*/];
  assign T1868 = T1869;
  assign T1869 = io_chanxy_in[10'h2d2/* 722*/:10'h2ca/* 714*/];
  assign T1870 = T1871;
  assign T1871 = T1872;
  assign T1872 = T1876[T1873];
  assign T1873 = T1874;
  assign T1874 = T1875;
  assign T1875 = io_chanxy_config[9'h157/* 343*/:9'h157/* 343*/];
  assign T1876 = T1877;
  assign T1877 = io_chanxy_in[10'h2d4/* 724*/:10'h2d3/* 723*/];
  assign T1878 = T1879;
  assign T1879 = T1880;
  assign T1880 = T1884[T1881];
  assign T1881 = T1882;
  assign T1882 = T1883;
  assign T1883 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1884 = T1885;
  assign T1885 = io_chanxy_in[10'h2d6/* 726*/:10'h2d5/* 725*/];
  assign T1886 = T1887;
  assign T1887 = T1888;
  assign T1888 = T1892[T1889];
  assign T1889 = T1890;
  assign T1890 = T1891;
  assign T1891 = io_chanxy_config[9'h159/* 345*/:9'h159/* 345*/];
  assign T1892 = T1893;
  assign T1893 = io_chanxy_in[10'h2d8/* 728*/:10'h2d7/* 727*/];
  assign T1894 = T1895;
  assign T1895 = T1896;
  assign T1896 = T1900[T1897];
  assign T1897 = T1898;
  assign T1898 = T1899;
  assign T1899 = io_chanxy_config[9'h15a/* 346*/:9'h15a/* 346*/];
  assign T1900 = T1901;
  assign T1901 = io_chanxy_in[10'h2da/* 730*/:10'h2d9/* 729*/];
  assign T1902 = T1903;
  assign T1903 = T1904;
  assign T1904 = T1908[T1905];
  assign T1905 = T1906;
  assign T1906 = T1907;
  assign T1907 = io_chanxy_config[9'h15e/* 350*/:9'h15b/* 347*/];
  assign T1908 = T1909;
  assign T1909 = io_chanxy_in[10'h2e3/* 739*/:10'h2db/* 731*/];
  assign T1910 = T1911;
  assign T1911 = T1912;
  assign T1912 = T1916[T1913];
  assign T1913 = T1914;
  assign T1914 = T1915;
  assign T1915 = io_chanxy_config[9'h15f/* 351*/:9'h15f/* 351*/];
  assign T1916 = T1917;
  assign T1917 = io_chanxy_in[10'h2e5/* 741*/:10'h2e4/* 740*/];
  assign T1918 = T1919;
  assign T1919 = T1920;
  assign T1920 = T1924[T1921];
  assign T1921 = T1922;
  assign T1922 = T1923;
  assign T1923 = io_chanxy_config[9'h160/* 352*/:9'h160/* 352*/];
  assign T1924 = T1925;
  assign T1925 = io_chanxy_in[10'h2e7/* 743*/:10'h2e6/* 742*/];
  assign T1926 = T1927;
  assign T1927 = T1928;
  assign T1928 = T1932[T1929];
  assign T1929 = T1930;
  assign T1930 = T1931;
  assign T1931 = io_chanxy_config[9'h161/* 353*/:9'h161/* 353*/];
  assign T1932 = T1933;
  assign T1933 = io_chanxy_in[10'h2e9/* 745*/:10'h2e8/* 744*/];
  assign T1934 = T1935;
  assign T1935 = T1936;
  assign T1936 = T1940[T1937];
  assign T1937 = T1938;
  assign T1938 = T1939;
  assign T1939 = io_chanxy_config[9'h162/* 354*/:9'h162/* 354*/];
  assign T1940 = T1941;
  assign T1941 = io_chanxy_in[10'h2eb/* 747*/:10'h2ea/* 746*/];
  assign T1942 = T1943;
  assign T1943 = T1944;
  assign T1944 = T1948[T1945];
  assign T1945 = T1946;
  assign T1946 = T1947;
  assign T1947 = io_chanxy_config[9'h166/* 358*/:9'h163/* 355*/];
  assign T1948 = T1949;
  assign T1949 = io_chanxy_in[10'h2f4/* 756*/:10'h2ec/* 748*/];
  assign T1950 = T1951;
  assign T1951 = T1952;
  assign T1952 = T1956[T1953];
  assign T1953 = T1954;
  assign T1954 = T1955;
  assign T1955 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1956 = T1957;
  assign T1957 = io_chanxy_in[10'h2f6/* 758*/:10'h2f5/* 757*/];
  assign T1958 = T1959;
  assign T1959 = T1960;
  assign T1960 = T1964[T1961];
  assign T1961 = T1962;
  assign T1962 = T1963;
  assign T1963 = io_chanxy_config[9'h168/* 360*/:9'h168/* 360*/];
  assign T1964 = T1965;
  assign T1965 = io_chanxy_in[10'h2f8/* 760*/:10'h2f7/* 759*/];
  assign T1966 = T1967;
  assign T1967 = T1968;
  assign T1968 = T1972[T1969];
  assign T1969 = T1970;
  assign T1970 = T1971;
  assign T1971 = io_chanxy_config[9'h169/* 361*/:9'h169/* 361*/];
  assign T1972 = T1973;
  assign T1973 = io_chanxy_in[10'h2fa/* 762*/:10'h2f9/* 761*/];
  assign T1974 = T1975;
  assign T1975 = T1976;
  assign T1976 = T1980[T1977];
  assign T1977 = T1978;
  assign T1978 = T1979;
  assign T1979 = io_chanxy_config[9'h16a/* 362*/:9'h16a/* 362*/];
  assign T1980 = T1981;
  assign T1981 = io_chanxy_in[10'h2fc/* 764*/:10'h2fb/* 763*/];
  assign T1982 = T1983;
  assign T1983 = T1984;
  assign T1984 = T1988[T1985];
  assign T1985 = T1986;
  assign T1986 = T1987;
  assign T1987 = io_chanxy_config[9'h16e/* 366*/:9'h16b/* 363*/];
  assign T1988 = T1989;
  assign T1989 = io_chanxy_in[10'h305/* 773*/:10'h2fd/* 765*/];
  assign T1990 = T1991;
  assign T1991 = T1992;
  assign T1992 = T1996[T1993];
  assign T1993 = T1994;
  assign T1994 = T1995;
  assign T1995 = io_chanxy_config[9'h16f/* 367*/:9'h16f/* 367*/];
  assign T1996 = T1997;
  assign T1997 = io_chanxy_in[10'h307/* 775*/:10'h306/* 774*/];
  assign io_ipin_out = T1998;
  assign T1998 = T1999;
  assign T1999 = {T2318, T2000};
  assign T2000 = T2001;
  assign T2001 = {T2310, T2002};
  assign T2002 = T2003;
  assign T2003 = {T2302, T2004};
  assign T2004 = T2005;
  assign T2005 = {T2294, T2006};
  assign T2006 = T2007;
  assign T2007 = {T2286, T2008};
  assign T2008 = T2009;
  assign T2009 = {T2278, T2010};
  assign T2010 = T2011;
  assign T2011 = {T2270, T2012};
  assign T2012 = T2013;
  assign T2013 = {T2262, T2014};
  assign T2014 = T2015;
  assign T2015 = {T2254, T2016};
  assign T2016 = T2017;
  assign T2017 = {T2246, T2018};
  assign T2018 = T2019;
  assign T2019 = {T2238, T2020};
  assign T2020 = T2021;
  assign T2021 = {T2230, T2022};
  assign T2022 = T2023;
  assign T2023 = {T2222, T2024};
  assign T2024 = T2025;
  assign T2025 = {T2214, T2026};
  assign T2026 = T2027;
  assign T2027 = {T2206, T2028};
  assign T2028 = T2029;
  assign T2029 = {T2198, T2030};
  assign T2030 = T2031;
  assign T2031 = {T2190, T2032};
  assign T2032 = T2033;
  assign T2033 = {T2182, T2034};
  assign T2034 = T2035;
  assign T2035 = {T2174, T2036};
  assign T2036 = T2037;
  assign T2037 = {T2166, T2038};
  assign T2038 = T2039;
  assign T2039 = {T2158, T2040};
  assign T2040 = T2041;
  assign T2041 = {T2150, T2042};
  assign T2042 = T2043;
  assign T2043 = {T2142, T2044};
  assign T2044 = T2045;
  assign T2045 = {T2134, T2046};
  assign T2046 = T2047;
  assign T2047 = {T2126, T2048};
  assign T2048 = T2049;
  assign T2049 = {T2118, T2050};
  assign T2050 = T2051;
  assign T2051 = {T2110, T2052};
  assign T2052 = T2053;
  assign T2053 = {T2102, T2054};
  assign T2054 = T2055;
  assign T2055 = {T2094, T2056};
  assign T2056 = T2057;
  assign T2057 = {T2086, T2058};
  assign T2058 = T2059;
  assign T2059 = {T2078, T2060};
  assign T2060 = T2061;
  assign T2061 = {T2070, T2062};
  assign T2062 = T2063;
  assign T2063 = T2064;
  assign T2064 = T2068[T2065];
  assign T2065 = T2066;
  assign T2066 = T2067;
  assign T2067 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T2068 = T2069;
  assign T2069 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T2070 = T2071;
  assign T2071 = T2072;
  assign T2072 = T2076[T2073];
  assign T2073 = T2074;
  assign T2074 = T2075;
  assign T2075 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T2076 = T2077;
  assign T2077 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T2078 = T2079;
  assign T2079 = T2080;
  assign T2080 = T2084[T2081];
  assign T2081 = T2082;
  assign T2082 = T2083;
  assign T2083 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T2084 = T2085;
  assign T2085 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T2086 = T2087;
  assign T2087 = T2088;
  assign T2088 = T2092[T2089];
  assign T2089 = T2090;
  assign T2090 = T2091;
  assign T2091 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T2092 = T2093;
  assign T2093 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T2094 = T2095;
  assign T2095 = T2096;
  assign T2096 = T2100[T2097];
  assign T2097 = T2098;
  assign T2098 = T2099;
  assign T2099 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T2100 = T2101;
  assign T2101 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T2102 = T2103;
  assign T2103 = T2104;
  assign T2104 = T2108[T2105];
  assign T2105 = T2106;
  assign T2106 = T2107;
  assign T2107 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T2108 = T2109;
  assign T2109 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T2110 = T2111;
  assign T2111 = T2112;
  assign T2112 = T2116[T2113];
  assign T2113 = T2114;
  assign T2114 = T2115;
  assign T2115 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T2116 = T2117;
  assign T2117 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T2118 = T2119;
  assign T2119 = T2120;
  assign T2120 = T2124[T2121];
  assign T2121 = T2122;
  assign T2122 = T2123;
  assign T2123 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T2124 = T2125;
  assign T2125 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T2126 = T2127;
  assign T2127 = T2128;
  assign T2128 = T2132[T2129];
  assign T2129 = T2130;
  assign T2130 = T2131;
  assign T2131 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T2132 = T2133;
  assign T2133 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T2134 = T2135;
  assign T2135 = T2136;
  assign T2136 = T2140[T2137];
  assign T2137 = T2138;
  assign T2138 = T2139;
  assign T2139 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T2140 = T2141;
  assign T2141 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T2142 = T2143;
  assign T2143 = T2144;
  assign T2144 = T2148[T2145];
  assign T2145 = T2146;
  assign T2146 = T2147;
  assign T2147 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T2148 = T2149;
  assign T2149 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T2150 = T2151;
  assign T2151 = T2152;
  assign T2152 = T2156[T2153];
  assign T2153 = T2154;
  assign T2154 = T2155;
  assign T2155 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T2156 = T2157;
  assign T2157 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T2158 = T2159;
  assign T2159 = T2160;
  assign T2160 = T2164[T2161];
  assign T2161 = T2162;
  assign T2162 = T2163;
  assign T2163 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T2164 = T2165;
  assign T2165 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T2166 = T2167;
  assign T2167 = T2168;
  assign T2168 = T2172[T2169];
  assign T2169 = T2170;
  assign T2170 = T2171;
  assign T2171 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T2172 = T2173;
  assign T2173 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T2174 = T2175;
  assign T2175 = T2176;
  assign T2176 = T2180[T2177];
  assign T2177 = T2178;
  assign T2178 = T2179;
  assign T2179 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T2180 = T2181;
  assign T2181 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T2182 = T2183;
  assign T2183 = T2184;
  assign T2184 = T2188[T2185];
  assign T2185 = T2186;
  assign T2186 = T2187;
  assign T2187 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T2188 = T2189;
  assign T2189 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T2190 = T2191;
  assign T2191 = T2192;
  assign T2192 = T2196[T2193];
  assign T2193 = T2194;
  assign T2194 = T2195;
  assign T2195 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T2196 = T2197;
  assign T2197 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T2198 = T2199;
  assign T2199 = T2200;
  assign T2200 = T2204[T2201];
  assign T2201 = T2202;
  assign T2202 = T2203;
  assign T2203 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T2204 = T2205;
  assign T2205 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T2206 = T2207;
  assign T2207 = T2208;
  assign T2208 = T2212[T2209];
  assign T2209 = T2210;
  assign T2210 = T2211;
  assign T2211 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T2212 = T2213;
  assign T2213 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T2214 = T2215;
  assign T2215 = T2216;
  assign T2216 = T2220[T2217];
  assign T2217 = T2218;
  assign T2218 = T2219;
  assign T2219 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T2220 = T2221;
  assign T2221 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T2222 = T2223;
  assign T2223 = T2224;
  assign T2224 = T2228[T2225];
  assign T2225 = T2226;
  assign T2226 = T2227;
  assign T2227 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T2228 = T2229;
  assign T2229 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T2230 = T2231;
  assign T2231 = T2232;
  assign T2232 = T2236[T2233];
  assign T2233 = T2234;
  assign T2234 = T2235;
  assign T2235 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T2236 = T2237;
  assign T2237 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T2238 = T2239;
  assign T2239 = T2240;
  assign T2240 = T2244[T2241];
  assign T2241 = T2242;
  assign T2242 = T2243;
  assign T2243 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T2244 = T2245;
  assign T2245 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T2246 = T2247;
  assign T2247 = T2248;
  assign T2248 = T2252[T2249];
  assign T2249 = T2250;
  assign T2250 = T2251;
  assign T2251 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T2252 = T2253;
  assign T2253 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T2254 = T2255;
  assign T2255 = T2256;
  assign T2256 = T2260[T2257];
  assign T2257 = T2258;
  assign T2258 = T2259;
  assign T2259 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T2260 = T2261;
  assign T2261 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T2262 = T2263;
  assign T2263 = T2264;
  assign T2264 = T2268[T2265];
  assign T2265 = T2266;
  assign T2266 = T2267;
  assign T2267 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T2268 = T2269;
  assign T2269 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T2270 = T2271;
  assign T2271 = T2272;
  assign T2272 = T2276[T2273];
  assign T2273 = T2274;
  assign T2274 = T2275;
  assign T2275 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T2276 = T2277;
  assign T2277 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T2278 = T2279;
  assign T2279 = T2280;
  assign T2280 = T2284[T2281];
  assign T2281 = T2282;
  assign T2282 = T2283;
  assign T2283 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T2284 = T2285;
  assign T2285 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T2286 = T2287;
  assign T2287 = T2288;
  assign T2288 = T2292[T2289];
  assign T2289 = T2290;
  assign T2290 = T2291;
  assign T2291 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T2292 = T2293;
  assign T2293 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T2294 = T2295;
  assign T2295 = T2296;
  assign T2296 = T2300[T2297];
  assign T2297 = T2298;
  assign T2298 = T2299;
  assign T2299 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T2300 = T2301;
  assign T2301 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T2302 = T2303;
  assign T2303 = T2304;
  assign T2304 = T2308[T2305];
  assign T2305 = T2306;
  assign T2306 = T2307;
  assign T2307 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T2308 = T2309;
  assign T2309 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T2310 = T2311;
  assign T2311 = T2312;
  assign T2312 = T2316[T2313];
  assign T2313 = T2314;
  assign T2314 = T2315;
  assign T2315 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T2316 = T2317;
  assign T2317 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T2318 = T2319;
  assign T2319 = T2320;
  assign T2320 = T2324[T2321];
  assign T2321 = T2322;
  assign T2322 = T2323;
  assign T2323 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T2324 = T2325;
  assign T2325 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_5(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [47:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [775:0] io_chanxy_in,
    output[199:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[367:0] T0;
  wire[1535:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[199:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5e5/* 1509*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_48 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_5 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_6(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [795:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[1:0] T281;
  wire[1:0] T282;
  wire[1:0] T283;
  wire[2:0] T284;
  wire[2:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[1:0] T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[2:0] T292;
  wire[2:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[1:0] T297;
  wire[1:0] T298;
  wire[1:0] T299;
  wire[2:0] T300;
  wire[2:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[1:0] T305;
  wire[1:0] T306;
  wire[1:0] T307;
  wire[2:0] T308;
  wire[2:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[1:0] T313;
  wire[1:0] T314;
  wire[1:0] T315;
  wire[2:0] T316;
  wire[2:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[1:0] T321;
  wire[1:0] T322;
  wire[1:0] T323;
  wire[2:0] T324;
  wire[2:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[1:0] T329;
  wire[1:0] T330;
  wire[1:0] T331;
  wire[2:0] T332;
  wire[2:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[1:0] T337;
  wire[1:0] T338;
  wire[1:0] T339;
  wire[2:0] T340;
  wire[2:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[1:0] T345;
  wire[1:0] T346;
  wire[1:0] T347;
  wire[2:0] T348;
  wire[2:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[2:0] T356;
  wire[2:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire[1:0] T364;
  wire[1:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire[1:0] T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire[1:0] T380;
  wire[1:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[1:0] T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  wire T394;
  wire T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[1:0] T441;
  wire[1:0] T442;
  wire[1:0] T443;
  wire[2:0] T444;
  wire[2:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[1:0] T449;
  wire[1:0] T450;
  wire[1:0] T451;
  wire[2:0] T452;
  wire[2:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[1:0] T457;
  wire[1:0] T458;
  wire[1:0] T459;
  wire[2:0] T460;
  wire[2:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[1:0] T465;
  wire[1:0] T466;
  wire[1:0] T467;
  wire[2:0] T468;
  wire[2:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[1:0] T473;
  wire[1:0] T474;
  wire[1:0] T475;
  wire[2:0] T476;
  wire[2:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[1:0] T481;
  wire[1:0] T482;
  wire[1:0] T483;
  wire[2:0] T484;
  wire[2:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[1:0] T489;
  wire[1:0] T490;
  wire[1:0] T491;
  wire[2:0] T492;
  wire[2:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[2:0] T500;
  wire[2:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[1:0] T505;
  wire[1:0] T506;
  wire[1:0] T507;
  wire[2:0] T508;
  wire[2:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[1:0] T513;
  wire[1:0] T514;
  wire[1:0] T515;
  wire[2:0] T516;
  wire[2:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[3:0] T761;
  wire[3:0] T762;
  wire[3:0] T763;
  wire[10:0] T764;
  wire[10:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[10:0] T780;
  wire[10:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[3:0] T793;
  wire[3:0] T794;
  wire[3:0] T795;
  wire[10:0] T796;
  wire[10:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire[1:0] T801;
  wire[1:0] T802;
  wire[1:0] T803;
  wire[2:0] T804;
  wire[2:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[3:0] T809;
  wire[3:0] T810;
  wire[3:0] T811;
  wire[10:0] T812;
  wire[10:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[1:0] T817;
  wire[1:0] T818;
  wire[1:0] T819;
  wire[2:0] T820;
  wire[2:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[3:0] T825;
  wire[3:0] T826;
  wire[3:0] T827;
  wire[10:0] T828;
  wire[10:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[1:0] T833;
  wire[1:0] T834;
  wire[1:0] T835;
  wire[2:0] T836;
  wire[2:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[3:0] T841;
  wire[3:0] T842;
  wire[3:0] T843;
  wire[10:0] T844;
  wire[10:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire[1:0] T849;
  wire[1:0] T850;
  wire[1:0] T851;
  wire[2:0] T852;
  wire[2:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[10:0] T860;
  wire[10:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[1:0] T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[2:0] T868;
  wire[2:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T875;
  wire[10:0] T876;
  wire[10:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[1:0] T881;
  wire[1:0] T882;
  wire[1:0] T883;
  wire[2:0] T884;
  wire[2:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[3:0] T890;
  wire[3:0] T891;
  wire[10:0] T892;
  wire[10:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[1:0] T897;
  wire[1:0] T898;
  wire[1:0] T899;
  wire[2:0] T900;
  wire[2:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[3:0] T905;
  wire[3:0] T906;
  wire[3:0] T907;
  wire[10:0] T908;
  wire[10:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[1:0] T913;
  wire[1:0] T914;
  wire[1:0] T915;
  wire[2:0] T916;
  wire[2:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[3:0] T921;
  wire[3:0] T922;
  wire[3:0] T923;
  wire[10:0] T924;
  wire[10:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire T929;
  wire T930;
  wire T931;
  wire[1:0] T932;
  wire[1:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[10:0] T940;
  wire[10:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire[1:0] T948;
  wire[1:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[3:0] T953;
  wire[3:0] T954;
  wire[3:0] T955;
  wire[10:0] T956;
  wire[10:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[1:0] T964;
  wire[1:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[3:0] T969;
  wire[3:0] T970;
  wire[3:0] T971;
  wire[10:0] T972;
  wire[10:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[1:0] T980;
  wire[1:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[3:0] T985;
  wire[3:0] T986;
  wire[3:0] T987;
  wire[10:0] T988;
  wire[10:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire[1:0] T996;
  wire[1:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire[3:0] T1001;
  wire[3:0] T1002;
  wire[3:0] T1003;
  wire[10:0] T1004;
  wire[10:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire[3:0] T1017;
  wire[3:0] T1018;
  wire[3:0] T1019;
  wire[10:0] T1020;
  wire[10:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[3:0] T1033;
  wire[3:0] T1034;
  wire[3:0] T1035;
  wire[10:0] T1036;
  wire[10:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire[3:0] T1049;
  wire[3:0] T1050;
  wire[3:0] T1051;
  wire[10:0] T1052;
  wire[10:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire[3:0] T1065;
  wire[3:0] T1066;
  wire[3:0] T1067;
  wire[10:0] T1068;
  wire[10:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire[3:0] T1081;
  wire[3:0] T1082;
  wire[3:0] T1083;
  wire[9:0] T1084;
  wire[9:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[9:0] T1092;
  wire[9:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[9:0] T1100;
  wire[9:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[9:0] T1108;
  wire[9:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[9:0] T1116;
  wire[9:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[9:0] T1124;
  wire[9:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[9:0] T1132;
  wire[9:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[9:0] T1140;
  wire[9:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[8:0] T1148;
  wire[8:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[8:0] T1156;
  wire[8:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire[3:0] T1161;
  wire[3:0] T1162;
  wire[3:0] T1163;
  wire[8:0] T1164;
  wire[8:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[8:0] T1172;
  wire[8:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[8:0] T1180;
  wire[8:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[8:0] T1188;
  wire[8:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[8:0] T1196;
  wire[8:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[3:0] T1201;
  wire[3:0] T1202;
  wire[3:0] T1203;
  wire[8:0] T1204;
  wire[8:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[8:0] T1212;
  wire[8:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[3:0] T1217;
  wire[3:0] T1218;
  wire[3:0] T1219;
  wire[8:0] T1220;
  wire[8:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[8:0] T1228;
  wire[8:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire[3:0] T1235;
  wire[8:0] T1236;
  wire[8:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[3:0] T1241;
  wire[3:0] T1242;
  wire[3:0] T1243;
  wire[9:0] T1244;
  wire[9:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[3:0] T1249;
  wire[3:0] T1250;
  wire[3:0] T1251;
  wire[9:0] T1252;
  wire[9:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[9:0] T1260;
  wire[9:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire[3:0] T1265;
  wire[3:0] T1266;
  wire[3:0] T1267;
  wire[9:0] T1268;
  wire[9:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[9:0] T1276;
  wire[9:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire[3:0] T1281;
  wire[3:0] T1282;
  wire[3:0] T1283;
  wire[9:0] T1284;
  wire[9:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[9:0] T1292;
  wire[9:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[3:0] T1297;
  wire[3:0] T1298;
  wire[3:0] T1299;
  wire[9:0] T1300;
  wire[9:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[8:0] T1308;
  wire[8:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[3:0] T1313;
  wire[3:0] T1314;
  wire[3:0] T1315;
  wire[8:0] T1316;
  wire[8:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[3:0] T1321;
  wire[3:0] T1322;
  wire[3:0] T1323;
  wire[8:0] T1324;
  wire[8:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[3:0] T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[8:0] T1332;
  wire[8:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[8:0] T1340;
  wire[8:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire[3:0] T1345;
  wire[3:0] T1346;
  wire[3:0] T1347;
  wire[8:0] T1348;
  wire[8:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[8:0] T1356;
  wire[8:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[3:0] T1361;
  wire[3:0] T1362;
  wire[3:0] T1363;
  wire[8:0] T1364;
  wire[8:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[8:0] T1372;
  wire[8:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire[3:0] T1379;
  wire[8:0] T1380;
  wire[8:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[8:0] T1388;
  wire[8:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[3:0] T1393;
  wire[3:0] T1394;
  wire[3:0] T1395;
  wire[8:0] T1396;
  wire[8:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[1'h1/* 1*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[2'h2/* 2*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[2'h3/* 3*/:2'h2/* 2*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[3'h5/* 5*/:2'h3/* 3*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[3'h5/* 5*/:3'h4/* 4*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[4'h8/* 8*/:3'h6/* 6*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[3'h7/* 7*/:3'h6/* 6*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[4'hb/* 11*/:4'h9/* 9*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[4'h9/* 9*/:4'h8/* 8*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[4'he/* 14*/:4'hc/* 12*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[4'hb/* 11*/:4'ha/* 10*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[5'h11/* 17*/:4'hf/* 15*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[4'hd/* 13*/:4'hc/* 12*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[5'h14/* 20*/:5'h12/* 18*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[4'hf/* 15*/:4'he/* 14*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[5'h17/* 23*/:5'h15/* 21*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[5'h11/* 17*/:5'h10/* 16*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[5'h1a/* 26*/:5'h18/* 24*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[5'h13/* 19*/:5'h12/* 18*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[5'h1d/* 29*/:5'h1b/* 27*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[6'h34/* 52*/:6'h32/* 50*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[6'h21/* 33*/:6'h20/* 32*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[6'h37/* 55*/:6'h35/* 53*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[6'h23/* 35*/:6'h22/* 34*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[6'h3a/* 58*/:6'h38/* 56*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[6'h25/* 37*/:6'h24/* 36*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[6'h3d/* 61*/:6'h3b/* 59*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[6'h27/* 39*/:6'h26/* 38*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[7'h40/* 64*/:6'h3e/* 62*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[6'h29/* 41*/:6'h28/* 40*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[7'h43/* 67*/:7'h41/* 65*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[7'h46/* 70*/:7'h44/* 68*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[7'h49/* 73*/:7'h47/* 71*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[7'h4c/* 76*/:7'h4a/* 74*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[6'h31/* 49*/:6'h30/* 48*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[7'h4f/* 79*/:7'h4d/* 77*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[6'h34/* 52*/:6'h34/* 52*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[7'h55/* 85*/:7'h54/* 84*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[6'h35/* 53*/:6'h35/* 53*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[7'h57/* 87*/:7'h56/* 86*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[7'h59/* 89*/:7'h58/* 88*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[7'h66/* 102*/:7'h64/* 100*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[7'h69/* 105*/:7'h67/* 103*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[7'h41/* 65*/:7'h40/* 64*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[7'h6c/* 108*/:7'h6a/* 106*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[7'h43/* 67*/:7'h42/* 66*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[7'h6f/* 111*/:7'h6d/* 109*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[7'h45/* 69*/:7'h44/* 68*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[7'h72/* 114*/:7'h70/* 112*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[7'h47/* 71*/:7'h46/* 70*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[7'h75/* 117*/:7'h73/* 115*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[7'h49/* 73*/:7'h48/* 72*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[7'h78/* 120*/:7'h76/* 118*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h7b/* 123*/:7'h79/* 121*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h7e/* 126*/:7'h7c/* 124*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[8'h81/* 129*/:7'h7f/* 127*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[7'h50/* 80*/:7'h50/* 80*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[8'h83/* 131*/:8'h82/* 130*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[7'h51/* 81*/:7'h51/* 81*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[8'h85/* 133*/:8'h84/* 132*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[7'h52/* 82*/:7'h52/* 82*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[8'h87/* 135*/:8'h86/* 134*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[7'h53/* 83*/:7'h53/* 83*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[8'h89/* 137*/:8'h88/* 136*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[7'h54/* 84*/:7'h54/* 84*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[8'h8b/* 139*/:8'h8a/* 138*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[7'h55/* 85*/:7'h55/* 85*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[7'h56/* 86*/:7'h56/* 86*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[7'h57/* 87*/:7'h57/* 87*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[8'h91/* 145*/:8'h90/* 144*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[7'h58/* 88*/:7'h58/* 88*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[8'h93/* 147*/:8'h92/* 146*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[8'h95/* 149*/:8'h94/* 148*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[8'ha0/* 160*/:8'h96/* 150*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[8'ha3/* 163*/:8'ha1/* 161*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[8'hae/* 174*/:8'ha4/* 164*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[7'h65/* 101*/:7'h64/* 100*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[8'hb1/* 177*/:8'haf/* 175*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[7'h69/* 105*/:7'h66/* 102*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[8'hbc/* 188*/:8'hb2/* 178*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[8'hbf/* 191*/:8'hbd/* 189*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[8'hca/* 202*/:8'hc0/* 192*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[7'h71/* 113*/:7'h70/* 112*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[8'hcd/* 205*/:8'hcb/* 203*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[7'h75/* 117*/:7'h72/* 114*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[8'hd8/* 216*/:8'hce/* 206*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[7'h77/* 119*/:7'h76/* 118*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[8'hdb/* 219*/:8'hd9/* 217*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[8'he6/* 230*/:8'hdc/* 220*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[7'h7d/* 125*/:7'h7c/* 124*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[8'he9/* 233*/:8'he7/* 231*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'h81/* 129*/:7'h7e/* 126*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[8'hf4/* 244*/:8'hea/* 234*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'h83/* 131*/:8'h82/* 130*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[8'hf7/* 247*/:8'hf5/* 245*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h102/* 258*/:8'hf8/* 248*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'h89/* 137*/:8'h88/* 136*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h105/* 261*/:9'h103/* 259*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'h8d/* 141*/:8'h8a/* 138*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h110/* 272*/:9'h106/* 262*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'h8f/* 143*/:8'h8e/* 142*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h113/* 275*/:9'h111/* 273*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h11e/* 286*/:9'h114/* 276*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'h95/* 149*/:8'h94/* 148*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h121/* 289*/:9'h11f/* 287*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h12c/* 300*/:9'h122/* 290*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h12e/* 302*/:9'h12d/* 301*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h139/* 313*/:9'h12f/* 303*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h13b/* 315*/:9'h13a/* 314*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'ha3/* 163*/:8'ha0/* 160*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h146/* 326*/:9'h13c/* 316*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'ha4/* 164*/:8'ha4/* 164*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'ha8/* 168*/:8'ha5/* 165*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h153/* 339*/:9'h149/* 329*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h155/* 341*/:9'h154/* 340*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'had/* 173*/:8'haa/* 170*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h160/* 352*/:9'h156/* 342*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h162/* 354*/:9'h161/* 353*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'hb2/* 178*/:8'haf/* 175*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h16d/* 365*/:9'h163/* 355*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h16f/* 367*/:9'h16e/* 366*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h17a/* 378*/:9'h170/* 368*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h17c/* 380*/:9'h17b/* 379*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'hbc/* 188*/:8'hb9/* 185*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h187/* 391*/:9'h17d/* 381*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h189/* 393*/:9'h188/* 392*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'hc1/* 193*/:8'hbe/* 190*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h194/* 404*/:9'h18a/* 394*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h196/* 406*/:9'h195/* 405*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hc6/* 198*/:8'hc3/* 195*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h1ad/* 429*/:9'h1a4/* 420*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h1b7/* 439*/:9'h1ae/* 430*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'hd3/* 211*/:8'hd0/* 208*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h1c1/* 449*/:9'h1b8/* 440*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h1cb/* 459*/:9'h1c2/* 450*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h1d5/* 469*/:9'h1cc/* 460*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'hdf/* 223*/:8'hdc/* 220*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h1df/* 479*/:9'h1d6/* 470*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h1e9/* 489*/:9'h1e0/* 480*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h1f3/* 499*/:9'h1ea/* 490*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[9'h1fc/* 508*/:9'h1f4/* 500*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h205/* 517*/:9'h1fd/* 509*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h20e/* 526*/:10'h206/* 518*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'hf7/* 247*/:8'hf4/* 244*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h217/* 535*/:10'h20f/* 527*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h220/* 544*/:10'h218/* 536*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h229/* 553*/:10'h221/* 545*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h232/* 562*/:10'h22a/* 554*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h23b/* 571*/:10'h233/* 563*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h10b/* 267*/:9'h108/* 264*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h244/* 580*/:10'h23c/* 572*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h24d/* 589*/:10'h245/* 581*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h113/* 275*/:9'h110/* 272*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h256/* 598*/:10'h24e/* 590*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h117/* 279*/:9'h114/* 276*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h25f/* 607*/:10'h257/* 599*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h269/* 617*/:10'h260/* 608*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h11f/* 287*/:9'h11c/* 284*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h273/* 627*/:10'h26a/* 618*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h123/* 291*/:9'h120/* 288*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h27d/* 637*/:10'h274/* 628*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h287/* 647*/:10'h27e/* 638*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h12b/* 299*/:9'h128/* 296*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h291/* 657*/:10'h288/* 648*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h12f/* 303*/:9'h12c/* 300*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h29b/* 667*/:10'h292/* 658*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h2a5/* 677*/:10'h29c/* 668*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h2af/* 687*/:10'h2a6/* 678*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h13b/* 315*/:9'h138/* 312*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h2b8/* 696*/:10'h2b0/* 688*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h13f/* 319*/:9'h13c/* 316*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h2c1/* 705*/:10'h2b9/* 697*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h2ca/* 714*/:10'h2c2/* 706*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h147/* 327*/:9'h144/* 324*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h2d3/* 723*/:10'h2cb/* 715*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h14b/* 331*/:9'h148/* 328*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h2dc/* 732*/:10'h2d4/* 724*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h14f/* 335*/:9'h14c/* 332*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h2e5/* 741*/:10'h2dd/* 733*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h153/* 339*/:9'h150/* 336*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h2ee/* 750*/:10'h2e6/* 742*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h2f7/* 759*/:10'h2ef/* 751*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h15b/* 347*/:9'h158/* 344*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h300/* 768*/:10'h2f8/* 760*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h15f/* 351*/:9'h15c/* 348*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h309/* 777*/:10'h301/* 769*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h163/* 355*/:9'h160/* 352*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h312/* 786*/:10'h30a/* 778*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h164/* 356*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h31b/* 795*/:10'h313/* 787*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_6(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [795:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_6 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_7(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [795:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_6 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_8(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [795:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_6 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


module sbcb_sp_7(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [695:0] io_chanxy_in,
    input [327:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[199:0] io_chanxy_out);

  wire[199:0] T0;
  wire[199:0] T1;
  wire[198:0] T2;
  wire[198:0] T3;
  wire[197:0] T4;
  wire[197:0] T5;
  wire[196:0] T6;
  wire[196:0] T7;
  wire[195:0] T8;
  wire[195:0] T9;
  wire[194:0] T10;
  wire[194:0] T11;
  wire[193:0] T12;
  wire[193:0] T13;
  wire[192:0] T14;
  wire[192:0] T15;
  wire[191:0] T16;
  wire[191:0] T17;
  wire[190:0] T18;
  wire[190:0] T19;
  wire[189:0] T20;
  wire[189:0] T21;
  wire[188:0] T22;
  wire[188:0] T23;
  wire[187:0] T24;
  wire[187:0] T25;
  wire[186:0] T26;
  wire[186:0] T27;
  wire[185:0] T28;
  wire[185:0] T29;
  wire[184:0] T30;
  wire[184:0] T31;
  wire[183:0] T32;
  wire[183:0] T33;
  wire[182:0] T34;
  wire[182:0] T35;
  wire[181:0] T36;
  wire[181:0] T37;
  wire[180:0] T38;
  wire[180:0] T39;
  wire[179:0] T40;
  wire[179:0] T41;
  wire[178:0] T42;
  wire[178:0] T43;
  wire[177:0] T44;
  wire[177:0] T45;
  wire[176:0] T46;
  wire[176:0] T47;
  wire[175:0] T48;
  wire[175:0] T49;
  wire[174:0] T50;
  wire[174:0] T51;
  wire[173:0] T52;
  wire[173:0] T53;
  wire[172:0] T54;
  wire[172:0] T55;
  wire[171:0] T56;
  wire[171:0] T57;
  wire[170:0] T58;
  wire[170:0] T59;
  wire[169:0] T60;
  wire[169:0] T61;
  wire[168:0] T62;
  wire[168:0] T63;
  wire[167:0] T64;
  wire[167:0] T65;
  wire[166:0] T66;
  wire[166:0] T67;
  wire[165:0] T68;
  wire[165:0] T69;
  wire[164:0] T70;
  wire[164:0] T71;
  wire[163:0] T72;
  wire[163:0] T73;
  wire[162:0] T74;
  wire[162:0] T75;
  wire[161:0] T76;
  wire[161:0] T77;
  wire[160:0] T78;
  wire[160:0] T79;
  wire[159:0] T80;
  wire[159:0] T81;
  wire[158:0] T82;
  wire[158:0] T83;
  wire[157:0] T84;
  wire[157:0] T85;
  wire[156:0] T86;
  wire[156:0] T87;
  wire[155:0] T88;
  wire[155:0] T89;
  wire[154:0] T90;
  wire[154:0] T91;
  wire[153:0] T92;
  wire[153:0] T93;
  wire[152:0] T94;
  wire[152:0] T95;
  wire[151:0] T96;
  wire[151:0] T97;
  wire[150:0] T98;
  wire[150:0] T99;
  wire[149:0] T100;
  wire[149:0] T101;
  wire[148:0] T102;
  wire[148:0] T103;
  wire[147:0] T104;
  wire[147:0] T105;
  wire[146:0] T106;
  wire[146:0] T107;
  wire[145:0] T108;
  wire[145:0] T109;
  wire[144:0] T110;
  wire[144:0] T111;
  wire[143:0] T112;
  wire[143:0] T113;
  wire[142:0] T114;
  wire[142:0] T115;
  wire[141:0] T116;
  wire[141:0] T117;
  wire[140:0] T118;
  wire[140:0] T119;
  wire[139:0] T120;
  wire[139:0] T121;
  wire[138:0] T122;
  wire[138:0] T123;
  wire[137:0] T124;
  wire[137:0] T125;
  wire[136:0] T126;
  wire[136:0] T127;
  wire[135:0] T128;
  wire[135:0] T129;
  wire[134:0] T130;
  wire[134:0] T131;
  wire[133:0] T132;
  wire[133:0] T133;
  wire[132:0] T134;
  wire[132:0] T135;
  wire[131:0] T136;
  wire[131:0] T137;
  wire[130:0] T138;
  wire[130:0] T139;
  wire[129:0] T140;
  wire[129:0] T141;
  wire[128:0] T142;
  wire[128:0] T143;
  wire[127:0] T144;
  wire[127:0] T145;
  wire[126:0] T146;
  wire[126:0] T147;
  wire[125:0] T148;
  wire[125:0] T149;
  wire[124:0] T150;
  wire[124:0] T151;
  wire[123:0] T152;
  wire[123:0] T153;
  wire[122:0] T154;
  wire[122:0] T155;
  wire[121:0] T156;
  wire[121:0] T157;
  wire[120:0] T158;
  wire[120:0] T159;
  wire[119:0] T160;
  wire[119:0] T161;
  wire[118:0] T162;
  wire[118:0] T163;
  wire[117:0] T164;
  wire[117:0] T165;
  wire[116:0] T166;
  wire[116:0] T167;
  wire[115:0] T168;
  wire[115:0] T169;
  wire[114:0] T170;
  wire[114:0] T171;
  wire[113:0] T172;
  wire[113:0] T173;
  wire[112:0] T174;
  wire[112:0] T175;
  wire[111:0] T176;
  wire[111:0] T177;
  wire[110:0] T178;
  wire[110:0] T179;
  wire[109:0] T180;
  wire[109:0] T181;
  wire[108:0] T182;
  wire[108:0] T183;
  wire[107:0] T184;
  wire[107:0] T185;
  wire[106:0] T186;
  wire[106:0] T187;
  wire[105:0] T188;
  wire[105:0] T189;
  wire[104:0] T190;
  wire[104:0] T191;
  wire[103:0] T192;
  wire[103:0] T193;
  wire[102:0] T194;
  wire[102:0] T195;
  wire[101:0] T196;
  wire[101:0] T197;
  wire[100:0] T198;
  wire[100:0] T199;
  wire[99:0] T200;
  wire[99:0] T201;
  wire[98:0] T202;
  wire[98:0] T203;
  wire[97:0] T204;
  wire[97:0] T205;
  wire[96:0] T206;
  wire[96:0] T207;
  wire[95:0] T208;
  wire[95:0] T209;
  wire[94:0] T210;
  wire[94:0] T211;
  wire[93:0] T212;
  wire[93:0] T213;
  wire[92:0] T214;
  wire[92:0] T215;
  wire[91:0] T216;
  wire[91:0] T217;
  wire[90:0] T218;
  wire[90:0] T219;
  wire[89:0] T220;
  wire[89:0] T221;
  wire[88:0] T222;
  wire[88:0] T223;
  wire[87:0] T224;
  wire[87:0] T225;
  wire[86:0] T226;
  wire[86:0] T227;
  wire[85:0] T228;
  wire[85:0] T229;
  wire[84:0] T230;
  wire[84:0] T231;
  wire[83:0] T232;
  wire[83:0] T233;
  wire[82:0] T234;
  wire[82:0] T235;
  wire[81:0] T236;
  wire[81:0] T237;
  wire[80:0] T238;
  wire[80:0] T239;
  wire[79:0] T240;
  wire[79:0] T241;
  wire[78:0] T242;
  wire[78:0] T243;
  wire[77:0] T244;
  wire[77:0] T245;
  wire[76:0] T246;
  wire[76:0] T247;
  wire[75:0] T248;
  wire[75:0] T249;
  wire[74:0] T250;
  wire[74:0] T251;
  wire[73:0] T252;
  wire[73:0] T253;
  wire[72:0] T254;
  wire[72:0] T255;
  wire[71:0] T256;
  wire[71:0] T257;
  wire[70:0] T258;
  wire[70:0] T259;
  wire[69:0] T260;
  wire[69:0] T261;
  wire[68:0] T262;
  wire[68:0] T263;
  wire[67:0] T264;
  wire[67:0] T265;
  wire[66:0] T266;
  wire[66:0] T267;
  wire[65:0] T268;
  wire[65:0] T269;
  wire[64:0] T270;
  wire[64:0] T271;
  wire[63:0] T272;
  wire[63:0] T273;
  wire[62:0] T274;
  wire[62:0] T275;
  wire[61:0] T276;
  wire[61:0] T277;
  wire[60:0] T278;
  wire[60:0] T279;
  wire[59:0] T280;
  wire[59:0] T281;
  wire[58:0] T282;
  wire[58:0] T283;
  wire[57:0] T284;
  wire[57:0] T285;
  wire[56:0] T286;
  wire[56:0] T287;
  wire[55:0] T288;
  wire[55:0] T289;
  wire[54:0] T290;
  wire[54:0] T291;
  wire[53:0] T292;
  wire[53:0] T293;
  wire[52:0] T294;
  wire[52:0] T295;
  wire[51:0] T296;
  wire[51:0] T297;
  wire[50:0] T298;
  wire[50:0] T299;
  wire[49:0] T300;
  wire[49:0] T301;
  wire[48:0] T302;
  wire[48:0] T303;
  wire[47:0] T304;
  wire[47:0] T305;
  wire[46:0] T306;
  wire[46:0] T307;
  wire[45:0] T308;
  wire[45:0] T309;
  wire[44:0] T310;
  wire[44:0] T311;
  wire[43:0] T312;
  wire[43:0] T313;
  wire[42:0] T314;
  wire[42:0] T315;
  wire[41:0] T316;
  wire[41:0] T317;
  wire[40:0] T318;
  wire[40:0] T319;
  wire[39:0] T320;
  wire[39:0] T321;
  wire[38:0] T322;
  wire[38:0] T323;
  wire[37:0] T324;
  wire[37:0] T325;
  wire[36:0] T326;
  wire[36:0] T327;
  wire[35:0] T328;
  wire[35:0] T329;
  wire[34:0] T330;
  wire[34:0] T331;
  wire[33:0] T332;
  wire[33:0] T333;
  wire[32:0] T334;
  wire[32:0] T335;
  wire[31:0] T336;
  wire[31:0] T337;
  wire[30:0] T338;
  wire[30:0] T339;
  wire[29:0] T340;
  wire[29:0] T341;
  wire[28:0] T342;
  wire[28:0] T343;
  wire[27:0] T344;
  wire[27:0] T345;
  wire[26:0] T346;
  wire[26:0] T347;
  wire[25:0] T348;
  wire[25:0] T349;
  wire[24:0] T350;
  wire[24:0] T351;
  wire[23:0] T352;
  wire[23:0] T353;
  wire[22:0] T354;
  wire[22:0] T355;
  wire[21:0] T356;
  wire[21:0] T357;
  wire[20:0] T358;
  wire[20:0] T359;
  wire[19:0] T360;
  wire[19:0] T361;
  wire[18:0] T362;
  wire[18:0] T363;
  wire[17:0] T364;
  wire[17:0] T365;
  wire[16:0] T366;
  wire[16:0] T367;
  wire[15:0] T368;
  wire[15:0] T369;
  wire[14:0] T370;
  wire[14:0] T371;
  wire[13:0] T372;
  wire[13:0] T373;
  wire[12:0] T374;
  wire[12:0] T375;
  wire[11:0] T376;
  wire[11:0] T377;
  wire[10:0] T378;
  wire[10:0] T379;
  wire[9:0] T380;
  wire[9:0] T381;
  wire[8:0] T382;
  wire[8:0] T383;
  wire[7:0] T384;
  wire[7:0] T385;
  wire[6:0] T386;
  wire[6:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[4:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[3:0] T393;
  wire[2:0] T394;
  wire[2:0] T395;
  wire[1:0] T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[1:0] T404;
  wire[1:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[1:0] T412;
  wire[1:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire[1:0] T420;
  wire[1:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire[1:0] T428;
  wire[1:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire[1:0] T436;
  wire[1:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire[1:0] T444;
  wire[1:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire[1:0] T452;
  wire[1:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire[1:0] T460;
  wire[1:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire[1:0] T468;
  wire[1:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire[1:0] T476;
  wire[1:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire[1:0] T484;
  wire[1:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire[1:0] T492;
  wire[1:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire T499;
  wire[1:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire[1:0] T508;
  wire[1:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire[1:0] T516;
  wire[1:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire[1:0] T524;
  wire[1:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[1:0] T532;
  wire[1:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire[1:0] T540;
  wire[1:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[1:0] T548;
  wire[1:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[1:0] T556;
  wire[1:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire[1:0] T564;
  wire[1:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire[1:0] T572;
  wire[1:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire T577;
  wire T578;
  wire T579;
  wire[1:0] T580;
  wire[1:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire T585;
  wire T586;
  wire T587;
  wire[1:0] T588;
  wire[1:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire T595;
  wire[1:0] T596;
  wire[1:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire[1:0] T604;
  wire[1:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire[1:0] T612;
  wire[1:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire[1:0] T620;
  wire[1:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire[1:0] T628;
  wire[1:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire[1:0] T636;
  wire[1:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire[1:0] T644;
  wire[1:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire[1:0] T652;
  wire[1:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire[1:0] T668;
  wire[1:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[1:0] T676;
  wire[1:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire[1:0] T764;
  wire[1:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire[1:0] T772;
  wire[1:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire[1:0] T780;
  wire[1:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire[1:0] T788;
  wire[1:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire[1:0] T796;
  wire[1:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire[1:0] T804;
  wire[1:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire[1:0] T812;
  wire[1:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[1:0] T820;
  wire[1:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire T825;
  wire T826;
  wire T827;
  wire[1:0] T828;
  wire[1:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[1:0] T836;
  wire[1:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[3:0] T881;
  wire[3:0] T882;
  wire[3:0] T883;
  wire[8:0] T884;
  wire[8:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[8:0] T900;
  wire[8:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[3:0] T913;
  wire[3:0] T914;
  wire[3:0] T915;
  wire[8:0] T916;
  wire[8:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire T921;
  wire T922;
  wire T923;
  wire[1:0] T924;
  wire[1:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[3:0] T929;
  wire[3:0] T930;
  wire[3:0] T931;
  wire[8:0] T932;
  wire[8:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire[1:0] T940;
  wire[1:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[3:0] T945;
  wire[3:0] T946;
  wire[3:0] T947;
  wire[8:0] T948;
  wire[8:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire[1:0] T956;
  wire[1:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[3:0] T961;
  wire[3:0] T962;
  wire[3:0] T963;
  wire[8:0] T964;
  wire[8:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire T969;
  wire T970;
  wire T971;
  wire[1:0] T972;
  wire[1:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[8:0] T980;
  wire[8:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[1:0] T988;
  wire[1:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[3:0] T993;
  wire[3:0] T994;
  wire[3:0] T995;
  wire[8:0] T996;
  wire[8:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire[3:0] T1009;
  wire[3:0] T1010;
  wire[3:0] T1011;
  wire[8:0] T1012;
  wire[8:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire[3:0] T1025;
  wire[3:0] T1026;
  wire[3:0] T1027;
  wire[8:0] T1028;
  wire[8:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire[3:0] T1041;
  wire[3:0] T1042;
  wire[3:0] T1043;
  wire[8:0] T1044;
  wire[8:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire[3:0] T1057;
  wire[3:0] T1058;
  wire[3:0] T1059;
  wire[8:0] T1060;
  wire[8:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire[3:0] T1073;
  wire[3:0] T1074;
  wire[3:0] T1075;
  wire[8:0] T1076;
  wire[8:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[8:0] T1092;
  wire[8:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[3:0] T1105;
  wire[3:0] T1106;
  wire[3:0] T1107;
  wire[8:0] T1108;
  wire[8:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[3:0] T1121;
  wire[3:0] T1122;
  wire[3:0] T1123;
  wire[8:0] T1124;
  wire[8:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[8:0] T1140;
  wire[8:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire[1:0] T1148;
  wire[1:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[8:0] T1156;
  wire[8:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[8:0] T1172;
  wire[8:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[3:0] T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[8:0] T1188;
  wire[8:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[1:0] T1201;
  wire[1:0] T1202;
  wire[1:0] T1203;
  wire[2:0] T1204;
  wire[2:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[1:0] T1209;
  wire[1:0] T1210;
  wire[1:0] T1211;
  wire[2:0] T1212;
  wire[2:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire[1:0] T1220;
  wire[1:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire[1:0] T1228;
  wire[1:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire[1:0] T1236;
  wire[1:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire[1:0] T1244;
  wire[1:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[1:0] T1252;
  wire[1:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire[1:0] T1260;
  wire[1:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[1:0] T1268;
  wire[1:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[1:0] T1276;
  wire[1:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire[1:0] T1292;
  wire[1:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire[1:0] T1308;
  wire[1:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire[1:0] T1340;
  wire[1:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire[1:0] T1356;
  wire[1:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[2:0] T1364;
  wire[2:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[1:0] T1369;
  wire[1:0] T1370;
  wire[1:0] T1371;
  wire[2:0] T1372;
  wire[2:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire[1:0] T1380;
  wire[1:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire[1:0] T1388;
  wire[1:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[1:0] T1396;
  wire[1:0] T1397;
  wire T1398;
  wire T1399;
  wire T1400;
  wire T1401;
  wire T1402;
  wire T1403;
  wire[1:0] T1404;
  wire[1:0] T1405;
  wire T1406;
  wire T1407;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire[1:0] T1412;
  wire[1:0] T1413;
  wire T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire[1:0] T1420;
  wire[1:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire[1:0] T1428;
  wire[1:0] T1429;
  wire T1430;
  wire T1431;
  wire T1432;
  wire T1433;
  wire T1434;
  wire T1435;
  wire[1:0] T1436;
  wire[1:0] T1437;
  wire T1438;
  wire T1439;
  wire T1440;
  wire T1441;
  wire T1442;
  wire T1443;
  wire[1:0] T1444;
  wire[1:0] T1445;
  wire T1446;
  wire T1447;
  wire T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire[1:0] T1452;
  wire[1:0] T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire T1458;
  wire T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire[1:0] T1468;
  wire[1:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire T1473;
  wire T1474;
  wire T1475;
  wire[1:0] T1476;
  wire[1:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire[1:0] T1484;
  wire[1:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire[1:0] T1492;
  wire[1:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire T1497;
  wire T1498;
  wire T1499;
  wire[1:0] T1500;
  wire[1:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire T1505;
  wire T1506;
  wire T1507;
  wire[1:0] T1508;
  wire[1:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire[1:0] T1516;
  wire[1:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[1:0] T1521;
  wire[1:0] T1522;
  wire[1:0] T1523;
  wire[2:0] T1524;
  wire[2:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[1:0] T1529;
  wire[1:0] T1530;
  wire[1:0] T1531;
  wire[2:0] T1532;
  wire[2:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire[1:0] T1540;
  wire[1:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire T1545;
  wire T1546;
  wire T1547;
  wire[1:0] T1548;
  wire[1:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire[1:0] T1556;
  wire[1:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire[1:0] T1564;
  wire[1:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire[1:0] T1572;
  wire[1:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire T1577;
  wire T1578;
  wire T1579;
  wire[1:0] T1580;
  wire[1:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire T1585;
  wire T1586;
  wire T1587;
  wire[1:0] T1588;
  wire[1:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire[1:0] T1596;
  wire[1:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire T1602;
  wire T1603;
  wire[1:0] T1604;
  wire[1:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire[1:0] T1612;
  wire[1:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire T1617;
  wire T1618;
  wire T1619;
  wire[1:0] T1620;
  wire[1:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire[1:0] T1628;
  wire[1:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire[1:0] T1636;
  wire[1:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire T1641;
  wire T1642;
  wire T1643;
  wire[1:0] T1644;
  wire[1:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire T1649;
  wire T1650;
  wire T1651;
  wire[1:0] T1652;
  wire[1:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire[1:0] T1660;
  wire[1:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire T1665;
  wire T1666;
  wire T1667;
  wire[1:0] T1668;
  wire[1:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire[1:0] T1676;
  wire[1:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[9:0] T1684;
  wire[9:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[1:0] T1689;
  wire[1:0] T1690;
  wire[1:0] T1691;
  wire[2:0] T1692;
  wire[2:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[9:0] T1700;
  wire[9:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[1:0] T1705;
  wire[1:0] T1706;
  wire[1:0] T1707;
  wire[2:0] T1708;
  wire[2:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[9:0] T1716;
  wire[9:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire T1723;
  wire[1:0] T1724;
  wire[1:0] T1725;
  wire T1726;
  wire T1727;
  wire T1728;
  wire[3:0] T1729;
  wire[3:0] T1730;
  wire[3:0] T1731;
  wire[9:0] T1732;
  wire[9:0] T1733;
  wire T1734;
  wire T1735;
  wire T1736;
  wire T1737;
  wire T1738;
  wire T1739;
  wire[1:0] T1740;
  wire[1:0] T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire[3:0] T1745;
  wire[3:0] T1746;
  wire[3:0] T1747;
  wire[9:0] T1748;
  wire[9:0] T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire T1753;
  wire T1754;
  wire T1755;
  wire[1:0] T1756;
  wire[1:0] T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire[3:0] T1761;
  wire[3:0] T1762;
  wire[3:0] T1763;
  wire[9:0] T1764;
  wire[9:0] T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire T1770;
  wire T1771;
  wire[1:0] T1772;
  wire[1:0] T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire[3:0] T1777;
  wire[3:0] T1778;
  wire[3:0] T1779;
  wire[9:0] T1780;
  wire[9:0] T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire[1:0] T1788;
  wire[1:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire[3:0] T1793;
  wire[3:0] T1794;
  wire[3:0] T1795;
  wire[9:0] T1796;
  wire[9:0] T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire[1:0] T1804;
  wire[1:0] T1805;
  wire T1806;
  wire T1807;
  wire T1808;
  wire[3:0] T1809;
  wire[3:0] T1810;
  wire[3:0] T1811;
  wire[8:0] T1812;
  wire[8:0] T1813;
  wire T1814;
  wire T1815;
  wire T1816;
  wire T1817;
  wire T1818;
  wire T1819;
  wire[1:0] T1820;
  wire[1:0] T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[3:0] T1825;
  wire[3:0] T1826;
  wire[3:0] T1827;
  wire[8:0] T1828;
  wire[8:0] T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire T1834;
  wire T1835;
  wire[1:0] T1836;
  wire[1:0] T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire[3:0] T1841;
  wire[3:0] T1842;
  wire[3:0] T1843;
  wire[8:0] T1844;
  wire[8:0] T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire T1851;
  wire[1:0] T1852;
  wire[1:0] T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire[3:0] T1857;
  wire[3:0] T1858;
  wire[3:0] T1859;
  wire[8:0] T1860;
  wire[8:0] T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[1:0] T1868;
  wire[1:0] T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire[3:0] T1873;
  wire[3:0] T1874;
  wire[3:0] T1875;
  wire[8:0] T1876;
  wire[8:0] T1877;
  wire T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire[1:0] T1884;
  wire[1:0] T1885;
  wire T1886;
  wire T1887;
  wire T1888;
  wire[3:0] T1889;
  wire[3:0] T1890;
  wire[3:0] T1891;
  wire[8:0] T1892;
  wire[8:0] T1893;
  wire T1894;
  wire T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire[1:0] T1900;
  wire[1:0] T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire[3:0] T1905;
  wire[3:0] T1906;
  wire[3:0] T1907;
  wire[8:0] T1908;
  wire[8:0] T1909;
  wire T1910;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire[1:0] T1916;
  wire[1:0] T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire[3:0] T1921;
  wire[3:0] T1922;
  wire[3:0] T1923;
  wire[8:0] T1924;
  wire[8:0] T1925;
  wire T1926;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire[1:0] T1932;
  wire[1:0] T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire[3:0] T1937;
  wire[3:0] T1938;
  wire[3:0] T1939;
  wire[8:0] T1940;
  wire[8:0] T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire T1945;
  wire T1946;
  wire T1947;
  wire[1:0] T1948;
  wire[1:0] T1949;
  wire T1950;
  wire T1951;
  wire T1952;
  wire[3:0] T1953;
  wire[3:0] T1954;
  wire[3:0] T1955;
  wire[8:0] T1956;
  wire[8:0] T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire T1961;
  wire T1962;
  wire T1963;
  wire[1:0] T1964;
  wire[1:0] T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire[3:0] T1969;
  wire[3:0] T1970;
  wire[3:0] T1971;
  wire[8:0] T1972;
  wire[8:0] T1973;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire T1979;
  wire[1:0] T1980;
  wire[1:0] T1981;
  wire T1982;
  wire T1983;
  wire T1984;
  wire[3:0] T1985;
  wire[3:0] T1986;
  wire[3:0] T1987;
  wire[8:0] T1988;
  wire[8:0] T1989;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire T1995;
  wire[1:0] T1996;
  wire[1:0] T1997;
  wire[32:0] T1998;
  wire[32:0] T1999;
  wire[31:0] T2000;
  wire[31:0] T2001;
  wire[30:0] T2002;
  wire[30:0] T2003;
  wire[29:0] T2004;
  wire[29:0] T2005;
  wire[28:0] T2006;
  wire[28:0] T2007;
  wire[27:0] T2008;
  wire[27:0] T2009;
  wire[26:0] T2010;
  wire[26:0] T2011;
  wire[25:0] T2012;
  wire[25:0] T2013;
  wire[24:0] T2014;
  wire[24:0] T2015;
  wire[23:0] T2016;
  wire[23:0] T2017;
  wire[22:0] T2018;
  wire[22:0] T2019;
  wire[21:0] T2020;
  wire[21:0] T2021;
  wire[20:0] T2022;
  wire[20:0] T2023;
  wire[19:0] T2024;
  wire[19:0] T2025;
  wire[18:0] T2026;
  wire[18:0] T2027;
  wire[17:0] T2028;
  wire[17:0] T2029;
  wire[16:0] T2030;
  wire[16:0] T2031;
  wire[15:0] T2032;
  wire[15:0] T2033;
  wire[14:0] T2034;
  wire[14:0] T2035;
  wire[13:0] T2036;
  wire[13:0] T2037;
  wire[12:0] T2038;
  wire[12:0] T2039;
  wire[11:0] T2040;
  wire[11:0] T2041;
  wire[10:0] T2042;
  wire[10:0] T2043;
  wire[9:0] T2044;
  wire[9:0] T2045;
  wire[8:0] T2046;
  wire[8:0] T2047;
  wire[7:0] T2048;
  wire[7:0] T2049;
  wire[6:0] T2050;
  wire[6:0] T2051;
  wire[5:0] T2052;
  wire[5:0] T2053;
  wire[4:0] T2054;
  wire[4:0] T2055;
  wire[3:0] T2056;
  wire[3:0] T2057;
  wire[2:0] T2058;
  wire[2:0] T2059;
  wire[1:0] T2060;
  wire[1:0] T2061;
  wire T2062;
  wire T2063;
  wire T2064;
  wire[3:0] T2065;
  wire[3:0] T2066;
  wire[3:0] T2067;
  wire[15:0] T2068;
  wire[15:0] T2069;
  wire T2070;
  wire T2071;
  wire T2072;
  wire[3:0] T2073;
  wire[3:0] T2074;
  wire[3:0] T2075;
  wire[15:0] T2076;
  wire[15:0] T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[3:0] T2081;
  wire[3:0] T2082;
  wire[3:0] T2083;
  wire[15:0] T2084;
  wire[15:0] T2085;
  wire T2086;
  wire T2087;
  wire T2088;
  wire[3:0] T2089;
  wire[3:0] T2090;
  wire[3:0] T2091;
  wire[15:0] T2092;
  wire[15:0] T2093;
  wire T2094;
  wire T2095;
  wire T2096;
  wire[3:0] T2097;
  wire[3:0] T2098;
  wire[3:0] T2099;
  wire[15:0] T2100;
  wire[15:0] T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire[3:0] T2105;
  wire[3:0] T2106;
  wire[3:0] T2107;
  wire[15:0] T2108;
  wire[15:0] T2109;
  wire T2110;
  wire T2111;
  wire T2112;
  wire[3:0] T2113;
  wire[3:0] T2114;
  wire[3:0] T2115;
  wire[15:0] T2116;
  wire[15:0] T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire[3:0] T2121;
  wire[3:0] T2122;
  wire[3:0] T2123;
  wire[15:0] T2124;
  wire[15:0] T2125;
  wire T2126;
  wire T2127;
  wire T2128;
  wire[3:0] T2129;
  wire[3:0] T2130;
  wire[3:0] T2131;
  wire[15:0] T2132;
  wire[15:0] T2133;
  wire T2134;
  wire T2135;
  wire T2136;
  wire[3:0] T2137;
  wire[3:0] T2138;
  wire[3:0] T2139;
  wire[15:0] T2140;
  wire[15:0] T2141;
  wire T2142;
  wire T2143;
  wire T2144;
  wire[3:0] T2145;
  wire[3:0] T2146;
  wire[3:0] T2147;
  wire[15:0] T2148;
  wire[15:0] T2149;
  wire T2150;
  wire T2151;
  wire T2152;
  wire[3:0] T2153;
  wire[3:0] T2154;
  wire[3:0] T2155;
  wire[15:0] T2156;
  wire[15:0] T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire[3:0] T2161;
  wire[3:0] T2162;
  wire[3:0] T2163;
  wire[15:0] T2164;
  wire[15:0] T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire[3:0] T2169;
  wire[3:0] T2170;
  wire[3:0] T2171;
  wire[15:0] T2172;
  wire[15:0] T2173;
  wire T2174;
  wire T2175;
  wire T2176;
  wire[3:0] T2177;
  wire[3:0] T2178;
  wire[3:0] T2179;
  wire[15:0] T2180;
  wire[15:0] T2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire[3:0] T2185;
  wire[3:0] T2186;
  wire[3:0] T2187;
  wire[15:0] T2188;
  wire[15:0] T2189;
  wire T2190;
  wire T2191;
  wire T2192;
  wire[3:0] T2193;
  wire[3:0] T2194;
  wire[3:0] T2195;
  wire[15:0] T2196;
  wire[15:0] T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  wire[3:0] T2201;
  wire[3:0] T2202;
  wire[3:0] T2203;
  wire[15:0] T2204;
  wire[15:0] T2205;
  wire T2206;
  wire T2207;
  wire T2208;
  wire[3:0] T2209;
  wire[3:0] T2210;
  wire[3:0] T2211;
  wire[15:0] T2212;
  wire[15:0] T2213;
  wire T2214;
  wire T2215;
  wire T2216;
  wire[3:0] T2217;
  wire[3:0] T2218;
  wire[3:0] T2219;
  wire[15:0] T2220;
  wire[15:0] T2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire[3:0] T2225;
  wire[3:0] T2226;
  wire[3:0] T2227;
  wire[15:0] T2228;
  wire[15:0] T2229;
  wire T2230;
  wire T2231;
  wire T2232;
  wire[3:0] T2233;
  wire[3:0] T2234;
  wire[3:0] T2235;
  wire[15:0] T2236;
  wire[15:0] T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  wire[3:0] T2241;
  wire[3:0] T2242;
  wire[3:0] T2243;
  wire[15:0] T2244;
  wire[15:0] T2245;
  wire T2246;
  wire T2247;
  wire T2248;
  wire[3:0] T2249;
  wire[3:0] T2250;
  wire[3:0] T2251;
  wire[15:0] T2252;
  wire[15:0] T2253;
  wire T2254;
  wire T2255;
  wire T2256;
  wire[3:0] T2257;
  wire[3:0] T2258;
  wire[3:0] T2259;
  wire[15:0] T2260;
  wire[15:0] T2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire[3:0] T2265;
  wire[3:0] T2266;
  wire[3:0] T2267;
  wire[15:0] T2268;
  wire[15:0] T2269;
  wire T2270;
  wire T2271;
  wire T2272;
  wire[3:0] T2273;
  wire[3:0] T2274;
  wire[3:0] T2275;
  wire[15:0] T2276;
  wire[15:0] T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  wire[3:0] T2281;
  wire[3:0] T2282;
  wire[3:0] T2283;
  wire[15:0] T2284;
  wire[15:0] T2285;
  wire T2286;
  wire T2287;
  wire T2288;
  wire[3:0] T2289;
  wire[3:0] T2290;
  wire[3:0] T2291;
  wire[15:0] T2292;
  wire[15:0] T2293;
  wire T2294;
  wire T2295;
  wire T2296;
  wire[3:0] T2297;
  wire[3:0] T2298;
  wire[3:0] T2299;
  wire[15:0] T2300;
  wire[15:0] T2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire[3:0] T2305;
  wire[3:0] T2306;
  wire[3:0] T2307;
  wire[15:0] T2308;
  wire[15:0] T2309;
  wire T2310;
  wire T2311;
  wire T2312;
  wire[3:0] T2313;
  wire[3:0] T2314;
  wire[3:0] T2315;
  wire[15:0] T2316;
  wire[15:0] T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  wire[3:0] T2321;
  wire[3:0] T2322;
  wire[3:0] T2323;
  wire[15:0] T2324;
  wire[15:0] T2325;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1990, T2};
  assign T2 = T3;
  assign T3 = {T1982, T4};
  assign T4 = T5;
  assign T5 = {T1974, T6};
  assign T6 = T7;
  assign T7 = {T1966, T8};
  assign T8 = T9;
  assign T9 = {T1958, T10};
  assign T10 = T11;
  assign T11 = {T1950, T12};
  assign T12 = T13;
  assign T13 = {T1942, T14};
  assign T14 = T15;
  assign T15 = {T1934, T16};
  assign T16 = T17;
  assign T17 = {T1926, T18};
  assign T18 = T19;
  assign T19 = {T1918, T20};
  assign T20 = T21;
  assign T21 = {T1910, T22};
  assign T22 = T23;
  assign T23 = {T1902, T24};
  assign T24 = T25;
  assign T25 = {T1894, T26};
  assign T26 = T27;
  assign T27 = {T1886, T28};
  assign T28 = T29;
  assign T29 = {T1878, T30};
  assign T30 = T31;
  assign T31 = {T1870, T32};
  assign T32 = T33;
  assign T33 = {T1862, T34};
  assign T34 = T35;
  assign T35 = {T1854, T36};
  assign T36 = T37;
  assign T37 = {T1846, T38};
  assign T38 = T39;
  assign T39 = {T1838, T40};
  assign T40 = T41;
  assign T41 = {T1830, T42};
  assign T42 = T43;
  assign T43 = {T1822, T44};
  assign T44 = T45;
  assign T45 = {T1814, T46};
  assign T46 = T47;
  assign T47 = {T1806, T48};
  assign T48 = T49;
  assign T49 = {T1798, T50};
  assign T50 = T51;
  assign T51 = {T1790, T52};
  assign T52 = T53;
  assign T53 = {T1782, T54};
  assign T54 = T55;
  assign T55 = {T1774, T56};
  assign T56 = T57;
  assign T57 = {T1766, T58};
  assign T58 = T59;
  assign T59 = {T1758, T60};
  assign T60 = T61;
  assign T61 = {T1750, T62};
  assign T62 = T63;
  assign T63 = {T1742, T64};
  assign T64 = T65;
  assign T65 = {T1734, T66};
  assign T66 = T67;
  assign T67 = {T1726, T68};
  assign T68 = T69;
  assign T69 = {T1718, T70};
  assign T70 = T71;
  assign T71 = {T1710, T72};
  assign T72 = T73;
  assign T73 = {T1702, T74};
  assign T74 = T75;
  assign T75 = {T1694, T76};
  assign T76 = T77;
  assign T77 = {T1686, T78};
  assign T78 = T79;
  assign T79 = {T1678, T80};
  assign T80 = T81;
  assign T81 = {T1670, T82};
  assign T82 = T83;
  assign T83 = {T1662, T84};
  assign T84 = T85;
  assign T85 = {T1654, T86};
  assign T86 = T87;
  assign T87 = {T1646, T88};
  assign T88 = T89;
  assign T89 = {T1638, T90};
  assign T90 = T91;
  assign T91 = {T1630, T92};
  assign T92 = T93;
  assign T93 = {T1622, T94};
  assign T94 = T95;
  assign T95 = {T1614, T96};
  assign T96 = T97;
  assign T97 = {T1606, T98};
  assign T98 = T99;
  assign T99 = {T1598, T100};
  assign T100 = T101;
  assign T101 = {T1590, T102};
  assign T102 = T103;
  assign T103 = {T1582, T104};
  assign T104 = T105;
  assign T105 = {T1574, T106};
  assign T106 = T107;
  assign T107 = {T1566, T108};
  assign T108 = T109;
  assign T109 = {T1558, T110};
  assign T110 = T111;
  assign T111 = {T1550, T112};
  assign T112 = T113;
  assign T113 = {T1542, T114};
  assign T114 = T115;
  assign T115 = {T1534, T116};
  assign T116 = T117;
  assign T117 = {T1526, T118};
  assign T118 = T119;
  assign T119 = {T1518, T120};
  assign T120 = T121;
  assign T121 = {T1510, T122};
  assign T122 = T123;
  assign T123 = {T1502, T124};
  assign T124 = T125;
  assign T125 = {T1494, T126};
  assign T126 = T127;
  assign T127 = {T1486, T128};
  assign T128 = T129;
  assign T129 = {T1478, T130};
  assign T130 = T131;
  assign T131 = {T1470, T132};
  assign T132 = T133;
  assign T133 = {T1462, T134};
  assign T134 = T135;
  assign T135 = {T1454, T136};
  assign T136 = T137;
  assign T137 = {T1446, T138};
  assign T138 = T139;
  assign T139 = {T1438, T140};
  assign T140 = T141;
  assign T141 = {T1430, T142};
  assign T142 = T143;
  assign T143 = {T1422, T144};
  assign T144 = T145;
  assign T145 = {T1414, T146};
  assign T146 = T147;
  assign T147 = {T1406, T148};
  assign T148 = T149;
  assign T149 = {T1398, T150};
  assign T150 = T151;
  assign T151 = {T1390, T152};
  assign T152 = T153;
  assign T153 = {T1382, T154};
  assign T154 = T155;
  assign T155 = {T1374, T156};
  assign T156 = T157;
  assign T157 = {T1366, T158};
  assign T158 = T159;
  assign T159 = {T1358, T160};
  assign T160 = T161;
  assign T161 = {T1350, T162};
  assign T162 = T163;
  assign T163 = {T1342, T164};
  assign T164 = T165;
  assign T165 = {T1334, T166};
  assign T166 = T167;
  assign T167 = {T1326, T168};
  assign T168 = T169;
  assign T169 = {T1318, T170};
  assign T170 = T171;
  assign T171 = {T1310, T172};
  assign T172 = T173;
  assign T173 = {T1302, T174};
  assign T174 = T175;
  assign T175 = {T1294, T176};
  assign T176 = T177;
  assign T177 = {T1286, T178};
  assign T178 = T179;
  assign T179 = {T1278, T180};
  assign T180 = T181;
  assign T181 = {T1270, T182};
  assign T182 = T183;
  assign T183 = {T1262, T184};
  assign T184 = T185;
  assign T185 = {T1254, T186};
  assign T186 = T187;
  assign T187 = {T1246, T188};
  assign T188 = T189;
  assign T189 = {T1238, T190};
  assign T190 = T191;
  assign T191 = {T1230, T192};
  assign T192 = T193;
  assign T193 = {T1222, T194};
  assign T194 = T195;
  assign T195 = {T1214, T196};
  assign T196 = T197;
  assign T197 = {T1206, T198};
  assign T198 = T199;
  assign T199 = {T1198, T200};
  assign T200 = T201;
  assign T201 = {T1190, T202};
  assign T202 = T203;
  assign T203 = {T1182, T204};
  assign T204 = T205;
  assign T205 = {T1174, T206};
  assign T206 = T207;
  assign T207 = {T1166, T208};
  assign T208 = T209;
  assign T209 = {T1158, T210};
  assign T210 = T211;
  assign T211 = {T1150, T212};
  assign T212 = T213;
  assign T213 = {T1142, T214};
  assign T214 = T215;
  assign T215 = {T1134, T216};
  assign T216 = T217;
  assign T217 = {T1126, T218};
  assign T218 = T219;
  assign T219 = {T1118, T220};
  assign T220 = T221;
  assign T221 = {T1110, T222};
  assign T222 = T223;
  assign T223 = {T1102, T224};
  assign T224 = T225;
  assign T225 = {T1094, T226};
  assign T226 = T227;
  assign T227 = {T1086, T228};
  assign T228 = T229;
  assign T229 = {T1078, T230};
  assign T230 = T231;
  assign T231 = {T1070, T232};
  assign T232 = T233;
  assign T233 = {T1062, T234};
  assign T234 = T235;
  assign T235 = {T1054, T236};
  assign T236 = T237;
  assign T237 = {T1046, T238};
  assign T238 = T239;
  assign T239 = {T1038, T240};
  assign T240 = T241;
  assign T241 = {T1030, T242};
  assign T242 = T243;
  assign T243 = {T1022, T244};
  assign T244 = T245;
  assign T245 = {T1014, T246};
  assign T246 = T247;
  assign T247 = {T1006, T248};
  assign T248 = T249;
  assign T249 = {T998, T250};
  assign T250 = T251;
  assign T251 = {T990, T252};
  assign T252 = T253;
  assign T253 = {T982, T254};
  assign T254 = T255;
  assign T255 = {T974, T256};
  assign T256 = T257;
  assign T257 = {T966, T258};
  assign T258 = T259;
  assign T259 = {T958, T260};
  assign T260 = T261;
  assign T261 = {T950, T262};
  assign T262 = T263;
  assign T263 = {T942, T264};
  assign T264 = T265;
  assign T265 = {T934, T266};
  assign T266 = T267;
  assign T267 = {T926, T268};
  assign T268 = T269;
  assign T269 = {T918, T270};
  assign T270 = T271;
  assign T271 = {T910, T272};
  assign T272 = T273;
  assign T273 = {T902, T274};
  assign T274 = T275;
  assign T275 = {T894, T276};
  assign T276 = T277;
  assign T277 = {T886, T278};
  assign T278 = T279;
  assign T279 = {T878, T280};
  assign T280 = T281;
  assign T281 = {T870, T282};
  assign T282 = T283;
  assign T283 = {T862, T284};
  assign T284 = T285;
  assign T285 = {T854, T286};
  assign T286 = T287;
  assign T287 = {T846, T288};
  assign T288 = T289;
  assign T289 = {T838, T290};
  assign T290 = T291;
  assign T291 = {T830, T292};
  assign T292 = T293;
  assign T293 = {T822, T294};
  assign T294 = T295;
  assign T295 = {T814, T296};
  assign T296 = T297;
  assign T297 = {T806, T298};
  assign T298 = T299;
  assign T299 = {T798, T300};
  assign T300 = T301;
  assign T301 = {T790, T302};
  assign T302 = T303;
  assign T303 = {T782, T304};
  assign T304 = T305;
  assign T305 = {T774, T306};
  assign T306 = T307;
  assign T307 = {T766, T308};
  assign T308 = T309;
  assign T309 = {T758, T310};
  assign T310 = T311;
  assign T311 = {T750, T312};
  assign T312 = T313;
  assign T313 = {T742, T314};
  assign T314 = T315;
  assign T315 = {T734, T316};
  assign T316 = T317;
  assign T317 = {T726, T318};
  assign T318 = T319;
  assign T319 = {T718, T320};
  assign T320 = T321;
  assign T321 = {T710, T322};
  assign T322 = T323;
  assign T323 = {T702, T324};
  assign T324 = T325;
  assign T325 = {T694, T326};
  assign T326 = T327;
  assign T327 = {T686, T328};
  assign T328 = T329;
  assign T329 = {T678, T330};
  assign T330 = T331;
  assign T331 = {T670, T332};
  assign T332 = T333;
  assign T333 = {T662, T334};
  assign T334 = T335;
  assign T335 = {T654, T336};
  assign T336 = T337;
  assign T337 = {T646, T338};
  assign T338 = T339;
  assign T339 = {T638, T340};
  assign T340 = T341;
  assign T341 = {T630, T342};
  assign T342 = T343;
  assign T343 = {T622, T344};
  assign T344 = T345;
  assign T345 = {T614, T346};
  assign T346 = T347;
  assign T347 = {T606, T348};
  assign T348 = T349;
  assign T349 = {T598, T350};
  assign T350 = T351;
  assign T351 = {T590, T352};
  assign T352 = T353;
  assign T353 = {T582, T354};
  assign T354 = T355;
  assign T355 = {T574, T356};
  assign T356 = T357;
  assign T357 = {T566, T358};
  assign T358 = T359;
  assign T359 = {T558, T360};
  assign T360 = T361;
  assign T361 = {T550, T362};
  assign T362 = T363;
  assign T363 = {T542, T364};
  assign T364 = T365;
  assign T365 = {T534, T366};
  assign T366 = T367;
  assign T367 = {T526, T368};
  assign T368 = T369;
  assign T369 = {T518, T370};
  assign T370 = T371;
  assign T371 = {T510, T372};
  assign T372 = T373;
  assign T373 = {T502, T374};
  assign T374 = T375;
  assign T375 = {T494, T376};
  assign T376 = T377;
  assign T377 = {T486, T378};
  assign T378 = T379;
  assign T379 = {T478, T380};
  assign T380 = T381;
  assign T381 = {T470, T382};
  assign T382 = T383;
  assign T383 = {T462, T384};
  assign T384 = T385;
  assign T385 = {T454, T386};
  assign T386 = T387;
  assign T387 = {T446, T388};
  assign T388 = T389;
  assign T389 = {T438, T390};
  assign T390 = T391;
  assign T391 = {T430, T392};
  assign T392 = T393;
  assign T393 = {T422, T394};
  assign T394 = T395;
  assign T395 = {T414, T396};
  assign T396 = T397;
  assign T397 = {T406, T398};
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[1'h0/* 0*/:1'h0/* 0*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[1'h1/* 1*/:1'h0/* 0*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[1'h1/* 1*/:1'h1/* 1*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[2'h3/* 3*/:2'h2/* 2*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[2'h2/* 2*/:2'h2/* 2*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[3'h5/* 5*/:3'h4/* 4*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[2'h3/* 3*/:2'h3/* 3*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[3'h7/* 7*/:3'h6/* 6*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[3'h4/* 4*/:3'h4/* 4*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[4'h9/* 9*/:4'h8/* 8*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[3'h5/* 5*/:3'h5/* 5*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[4'hb/* 11*/:4'ha/* 10*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[3'h6/* 6*/:3'h6/* 6*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[4'hd/* 13*/:4'hc/* 12*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[3'h7/* 7*/:3'h7/* 7*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[4'hf/* 15*/:4'he/* 14*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[4'h8/* 8*/:4'h8/* 8*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[5'h11/* 17*/:5'h10/* 16*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[4'h9/* 9*/:4'h9/* 9*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[5'h13/* 19*/:5'h12/* 18*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[4'ha/* 10*/:4'ha/* 10*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[5'h15/* 21*/:5'h14/* 20*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[4'hb/* 11*/:4'hb/* 11*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[5'h17/* 23*/:5'h16/* 22*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[4'hc/* 12*/:4'hc/* 12*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[5'h19/* 25*/:5'h18/* 24*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[4'hd/* 13*/:4'hd/* 13*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[5'h1b/* 27*/:5'h1a/* 26*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[4'he/* 14*/:4'he/* 14*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[5'h1d/* 29*/:5'h1c/* 28*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[4'hf/* 15*/:4'hf/* 15*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[5'h1f/* 31*/:5'h1e/* 30*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[5'h10/* 16*/:5'h10/* 16*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[6'h21/* 33*/:6'h20/* 32*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[5'h11/* 17*/:5'h11/* 17*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[6'h23/* 35*/:6'h22/* 34*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[5'h12/* 18*/:5'h12/* 18*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[6'h25/* 37*/:6'h24/* 36*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[5'h13/* 19*/:5'h13/* 19*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[6'h27/* 39*/:6'h26/* 38*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[5'h14/* 20*/:5'h14/* 20*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[6'h29/* 41*/:6'h28/* 40*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[5'h15/* 21*/:5'h15/* 21*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[6'h2b/* 43*/:6'h2a/* 42*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[5'h16/* 22*/:5'h16/* 22*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[6'h2d/* 45*/:6'h2c/* 44*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[5'h17/* 23*/:5'h17/* 23*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[6'h2f/* 47*/:6'h2e/* 46*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[5'h18/* 24*/:5'h18/* 24*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[6'h31/* 49*/:6'h30/* 48*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[5'h19/* 25*/:5'h19/* 25*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[6'h33/* 51*/:6'h32/* 50*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[5'h1a/* 26*/:5'h1a/* 26*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[6'h35/* 53*/:6'h34/* 52*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[5'h1b/* 27*/:5'h1b/* 27*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[6'h37/* 55*/:6'h36/* 54*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[5'h1c/* 28*/:5'h1c/* 28*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[6'h39/* 57*/:6'h38/* 56*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[5'h1d/* 29*/:5'h1d/* 29*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[6'h3b/* 59*/:6'h3a/* 58*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[5'h1e/* 30*/:5'h1e/* 30*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[6'h3d/* 61*/:6'h3c/* 60*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[5'h1f/* 31*/:5'h1f/* 31*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[6'h3f/* 63*/:6'h3e/* 62*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[6'h20/* 32*/:6'h20/* 32*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[7'h41/* 65*/:7'h40/* 64*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[6'h21/* 33*/:6'h21/* 33*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[7'h43/* 67*/:7'h42/* 66*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[6'h22/* 34*/:6'h22/* 34*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[7'h45/* 69*/:7'h44/* 68*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[6'h23/* 35*/:6'h23/* 35*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[7'h47/* 71*/:7'h46/* 70*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[6'h24/* 36*/:6'h24/* 36*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[7'h49/* 73*/:7'h48/* 72*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[6'h25/* 37*/:6'h25/* 37*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[7'h4b/* 75*/:7'h4a/* 74*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[6'h26/* 38*/:6'h26/* 38*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[7'h4d/* 77*/:7'h4c/* 76*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[6'h27/* 39*/:6'h27/* 39*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[7'h4f/* 79*/:7'h4e/* 78*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[6'h28/* 40*/:6'h28/* 40*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[7'h51/* 81*/:7'h50/* 80*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[6'h29/* 41*/:6'h29/* 41*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[7'h53/* 83*/:7'h52/* 82*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[6'h2a/* 42*/:6'h2a/* 42*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[7'h55/* 85*/:7'h54/* 84*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[6'h2b/* 43*/:6'h2b/* 43*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[7'h57/* 87*/:7'h56/* 86*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[6'h2c/* 44*/:6'h2c/* 44*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[7'h59/* 89*/:7'h58/* 88*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[6'h2d/* 45*/:6'h2d/* 45*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[7'h5b/* 91*/:7'h5a/* 90*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[6'h2e/* 46*/:6'h2e/* 46*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[7'h5d/* 93*/:7'h5c/* 92*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[6'h2f/* 47*/:6'h2f/* 47*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[7'h5f/* 95*/:7'h5e/* 94*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[6'h30/* 48*/:6'h30/* 48*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[7'h61/* 97*/:7'h60/* 96*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[6'h31/* 49*/:6'h31/* 49*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[7'h63/* 99*/:7'h62/* 98*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[6'h32/* 50*/:6'h32/* 50*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[7'h65/* 101*/:7'h64/* 100*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[6'h33/* 51*/:6'h33/* 51*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[7'h67/* 103*/:7'h66/* 102*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[6'h34/* 52*/:6'h34/* 52*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[7'h69/* 105*/:7'h68/* 104*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[6'h35/* 53*/:6'h35/* 53*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[7'h6b/* 107*/:7'h6a/* 106*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[6'h36/* 54*/:6'h36/* 54*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[7'h6d/* 109*/:7'h6c/* 108*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[6'h37/* 55*/:6'h37/* 55*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[7'h6f/* 111*/:7'h6e/* 110*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[6'h38/* 56*/:6'h38/* 56*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[7'h71/* 113*/:7'h70/* 112*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[6'h39/* 57*/:6'h39/* 57*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[7'h73/* 115*/:7'h72/* 114*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[6'h3a/* 58*/:6'h3a/* 58*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[7'h75/* 117*/:7'h74/* 116*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[6'h3b/* 59*/:6'h3b/* 59*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[7'h77/* 119*/:7'h76/* 118*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[8'h80/* 128*/:7'h78/* 120*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[7'h40/* 64*/:7'h40/* 64*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[8'h82/* 130*/:8'h81/* 129*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[7'h44/* 68*/:7'h41/* 65*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[8'h8b/* 139*/:8'h83/* 131*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[7'h45/* 69*/:7'h45/* 69*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[8'h8d/* 141*/:8'h8c/* 140*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[7'h49/* 73*/:7'h46/* 70*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[8'h96/* 150*/:8'h8e/* 142*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[7'h4a/* 74*/:7'h4a/* 74*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[8'h98/* 152*/:8'h97/* 151*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[7'h4e/* 78*/:7'h4b/* 75*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[8'ha1/* 161*/:8'h99/* 153*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[7'h4f/* 79*/:7'h4f/* 79*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[8'hac/* 172*/:8'ha4/* 164*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[7'h54/* 84*/:7'h54/* 84*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[8'hae/* 174*/:8'had/* 173*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[7'h58/* 88*/:7'h55/* 85*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[8'hb7/* 183*/:8'haf/* 175*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[7'h59/* 89*/:7'h59/* 89*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[7'h5d/* 93*/:7'h5a/* 90*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[8'hc2/* 194*/:8'hba/* 186*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[7'h5e/* 94*/:7'h5e/* 94*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[8'hc4/* 196*/:8'hc3/* 195*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[7'h62/* 98*/:7'h5f/* 95*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[8'hcd/* 205*/:8'hc5/* 197*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[7'h63/* 99*/:7'h63/* 99*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[8'hcf/* 207*/:8'hce/* 206*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[8'hd8/* 216*/:8'hd0/* 208*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[7'h68/* 104*/:7'h68/* 104*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[8'hda/* 218*/:8'hd9/* 217*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[7'h6c/* 108*/:7'h69/* 105*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[8'he3/* 227*/:8'hdb/* 219*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[7'h6d/* 109*/:7'h6d/* 109*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[8'he5/* 229*/:8'he4/* 228*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[7'h71/* 113*/:7'h6e/* 110*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[8'hee/* 238*/:8'he6/* 230*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[7'h72/* 114*/:7'h72/* 114*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[8'hf0/* 240*/:8'hef/* 239*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[7'h76/* 118*/:7'h73/* 115*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[8'hf9/* 249*/:8'hf1/* 241*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[7'h77/* 119*/:7'h77/* 119*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h104/* 260*/:8'hfc/* 252*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[7'h7c/* 124*/:7'h7c/* 124*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[9'h106/* 262*/:9'h105/* 261*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'h80/* 128*/:7'h7d/* 125*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[9'h10f/* 271*/:9'h107/* 263*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[8'h81/* 129*/:8'h81/* 129*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[9'h111/* 273*/:9'h110/* 272*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[8'h85/* 133*/:8'h82/* 130*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[9'h11a/* 282*/:9'h112/* 274*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[8'h86/* 134*/:8'h86/* 134*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[9'h11c/* 284*/:9'h11b/* 283*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[8'h8a/* 138*/:8'h87/* 135*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[9'h125/* 293*/:9'h11d/* 285*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[8'h8b/* 139*/:8'h8b/* 139*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[9'h127/* 295*/:9'h126/* 294*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[9'h130/* 304*/:9'h128/* 296*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[8'h90/* 144*/:8'h90/* 144*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[9'h132/* 306*/:9'h131/* 305*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[8'h94/* 148*/:8'h91/* 145*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[9'h13b/* 315*/:9'h133/* 307*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[8'h95/* 149*/:8'h95/* 149*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[9'h13d/* 317*/:9'h13c/* 316*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[8'h99/* 153*/:8'h96/* 150*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[9'h146/* 326*/:9'h13e/* 318*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[8'h9a/* 154*/:8'h9a/* 154*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[9'h148/* 328*/:9'h147/* 327*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[8'h9e/* 158*/:8'h9b/* 155*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[9'h151/* 337*/:9'h149/* 329*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[8'h9f/* 159*/:8'h9f/* 159*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[9'h153/* 339*/:9'h152/* 338*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[9'h156/* 342*/:9'h154/* 340*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[9'h159/* 345*/:9'h157/* 343*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[8'ha4/* 164*/:8'ha4/* 164*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[9'h15b/* 347*/:9'h15a/* 346*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[8'ha5/* 165*/:8'ha5/* 165*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[9'h15d/* 349*/:9'h15c/* 348*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[8'ha6/* 166*/:8'ha6/* 166*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[9'h15f/* 351*/:9'h15e/* 350*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[8'ha7/* 167*/:8'ha7/* 167*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[9'h161/* 353*/:9'h160/* 352*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[8'ha8/* 168*/:8'ha8/* 168*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[9'h163/* 355*/:9'h162/* 354*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[8'ha9/* 169*/:8'ha9/* 169*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[9'h165/* 357*/:9'h164/* 356*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[8'haa/* 170*/:8'haa/* 170*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[9'h167/* 359*/:9'h166/* 358*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[8'hab/* 171*/:8'hab/* 171*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[9'h169/* 361*/:9'h168/* 360*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[8'hac/* 172*/:8'hac/* 172*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[9'h16b/* 363*/:9'h16a/* 362*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[8'had/* 173*/:8'had/* 173*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[9'h16d/* 365*/:9'h16c/* 364*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[8'hae/* 174*/:8'hae/* 174*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[9'h16f/* 367*/:9'h16e/* 366*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[8'haf/* 175*/:8'haf/* 175*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[9'h171/* 369*/:9'h170/* 368*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[8'hb0/* 176*/:8'hb0/* 176*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[9'h173/* 371*/:9'h172/* 370*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[8'hb1/* 177*/:8'hb1/* 177*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[9'h175/* 373*/:9'h174/* 372*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[8'hb2/* 178*/:8'hb2/* 178*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[9'h177/* 375*/:9'h176/* 374*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[8'hb3/* 179*/:8'hb3/* 179*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[9'h179/* 377*/:9'h178/* 376*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[8'hb4/* 180*/:8'hb4/* 180*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[9'h17b/* 379*/:9'h17a/* 378*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[9'h17d/* 381*/:9'h17c/* 380*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[9'h180/* 384*/:9'h17e/* 382*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[9'h183/* 387*/:9'h181/* 385*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[9'h185/* 389*/:9'h184/* 388*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[8'hbb/* 187*/:8'hbb/* 187*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[9'h187/* 391*/:9'h186/* 390*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[8'hbc/* 188*/:8'hbc/* 188*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[9'h189/* 393*/:9'h188/* 392*/];
  assign T1398 = T1399;
  assign T1399 = T1400;
  assign T1400 = T1404[T1401];
  assign T1401 = T1402;
  assign T1402 = T1403;
  assign T1403 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T1404 = T1405;
  assign T1405 = io_chanxy_in[9'h18b/* 395*/:9'h18a/* 394*/];
  assign T1406 = T1407;
  assign T1407 = T1408;
  assign T1408 = T1412[T1409];
  assign T1409 = T1410;
  assign T1410 = T1411;
  assign T1411 = io_chanxy_config[8'hbe/* 190*/:8'hbe/* 190*/];
  assign T1412 = T1413;
  assign T1413 = io_chanxy_in[9'h18d/* 397*/:9'h18c/* 396*/];
  assign T1414 = T1415;
  assign T1415 = T1416;
  assign T1416 = T1420[T1417];
  assign T1417 = T1418;
  assign T1418 = T1419;
  assign T1419 = io_chanxy_config[8'hbf/* 191*/:8'hbf/* 191*/];
  assign T1420 = T1421;
  assign T1421 = io_chanxy_in[9'h18f/* 399*/:9'h18e/* 398*/];
  assign T1422 = T1423;
  assign T1423 = T1424;
  assign T1424 = T1428[T1425];
  assign T1425 = T1426;
  assign T1426 = T1427;
  assign T1427 = io_chanxy_config[8'hc0/* 192*/:8'hc0/* 192*/];
  assign T1428 = T1429;
  assign T1429 = io_chanxy_in[9'h191/* 401*/:9'h190/* 400*/];
  assign T1430 = T1431;
  assign T1431 = T1432;
  assign T1432 = T1436[T1433];
  assign T1433 = T1434;
  assign T1434 = T1435;
  assign T1435 = io_chanxy_config[8'hc1/* 193*/:8'hc1/* 193*/];
  assign T1436 = T1437;
  assign T1437 = io_chanxy_in[9'h193/* 403*/:9'h192/* 402*/];
  assign T1438 = T1439;
  assign T1439 = T1440;
  assign T1440 = T1444[T1441];
  assign T1441 = T1442;
  assign T1442 = T1443;
  assign T1443 = io_chanxy_config[8'hc2/* 194*/:8'hc2/* 194*/];
  assign T1444 = T1445;
  assign T1445 = io_chanxy_in[9'h195/* 405*/:9'h194/* 404*/];
  assign T1446 = T1447;
  assign T1447 = T1448;
  assign T1448 = T1452[T1449];
  assign T1449 = T1450;
  assign T1450 = T1451;
  assign T1451 = io_chanxy_config[8'hc3/* 195*/:8'hc3/* 195*/];
  assign T1452 = T1453;
  assign T1453 = io_chanxy_in[9'h197/* 407*/:9'h196/* 406*/];
  assign T1454 = T1455;
  assign T1455 = T1456;
  assign T1456 = T1460[T1457];
  assign T1457 = T1458;
  assign T1458 = T1459;
  assign T1459 = io_chanxy_config[8'hc4/* 196*/:8'hc4/* 196*/];
  assign T1460 = T1461;
  assign T1461 = io_chanxy_in[9'h199/* 409*/:9'h198/* 408*/];
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_chanxy_config[8'hc5/* 197*/:8'hc5/* 197*/];
  assign T1468 = T1469;
  assign T1469 = io_chanxy_in[9'h19b/* 411*/:9'h19a/* 410*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_chanxy_config[8'hc6/* 198*/:8'hc6/* 198*/];
  assign T1476 = T1477;
  assign T1477 = io_chanxy_in[9'h19d/* 413*/:9'h19c/* 412*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_chanxy_config[8'hc7/* 199*/:8'hc7/* 199*/];
  assign T1484 = T1485;
  assign T1485 = io_chanxy_in[9'h19f/* 415*/:9'h19e/* 414*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_chanxy_config[8'hc8/* 200*/:8'hc8/* 200*/];
  assign T1492 = T1493;
  assign T1493 = io_chanxy_in[9'h1a1/* 417*/:9'h1a0/* 416*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_chanxy_config[8'hc9/* 201*/:8'hc9/* 201*/];
  assign T1500 = T1501;
  assign T1501 = io_chanxy_in[9'h1a3/* 419*/:9'h1a2/* 418*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_chanxy_config[8'hca/* 202*/:8'hca/* 202*/];
  assign T1508 = T1509;
  assign T1509 = io_chanxy_in[9'h1a5/* 421*/:9'h1a4/* 420*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_chanxy_config[8'hcb/* 203*/:8'hcb/* 203*/];
  assign T1516 = T1517;
  assign T1517 = io_chanxy_in[9'h1a7/* 423*/:9'h1a6/* 422*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T1524 = T1525;
  assign T1525 = io_chanxy_in[9'h1aa/* 426*/:9'h1a8/* 424*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T1532 = T1533;
  assign T1533 = io_chanxy_in[9'h1ad/* 429*/:9'h1ab/* 427*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_chanxy_config[8'hd0/* 208*/:8'hd0/* 208*/];
  assign T1540 = T1541;
  assign T1541 = io_chanxy_in[9'h1af/* 431*/:9'h1ae/* 430*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_chanxy_config[8'hd1/* 209*/:8'hd1/* 209*/];
  assign T1548 = T1549;
  assign T1549 = io_chanxy_in[9'h1b1/* 433*/:9'h1b0/* 432*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T1556 = T1557;
  assign T1557 = io_chanxy_in[9'h1b3/* 435*/:9'h1b2/* 434*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_chanxy_config[8'hd3/* 211*/:8'hd3/* 211*/];
  assign T1564 = T1565;
  assign T1565 = io_chanxy_in[9'h1b5/* 437*/:9'h1b4/* 436*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_chanxy_config[8'hd4/* 212*/:8'hd4/* 212*/];
  assign T1572 = T1573;
  assign T1573 = io_chanxy_in[9'h1b7/* 439*/:9'h1b6/* 438*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_chanxy_config[8'hd5/* 213*/:8'hd5/* 213*/];
  assign T1580 = T1581;
  assign T1581 = io_chanxy_in[9'h1b9/* 441*/:9'h1b8/* 440*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T1588 = T1589;
  assign T1589 = io_chanxy_in[9'h1bb/* 443*/:9'h1ba/* 442*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T1596 = T1597;
  assign T1597 = io_chanxy_in[9'h1bd/* 445*/:9'h1bc/* 444*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T1604 = T1605;
  assign T1605 = io_chanxy_in[9'h1bf/* 447*/:9'h1be/* 446*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T1612 = T1613;
  assign T1613 = io_chanxy_in[9'h1c1/* 449*/:9'h1c0/* 448*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T1620 = T1621;
  assign T1621 = io_chanxy_in[9'h1c3/* 451*/:9'h1c2/* 450*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T1628 = T1629;
  assign T1629 = io_chanxy_in[9'h1c5/* 453*/:9'h1c4/* 452*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_chanxy_config[8'hdc/* 220*/:8'hdc/* 220*/];
  assign T1636 = T1637;
  assign T1637 = io_chanxy_in[9'h1c7/* 455*/:9'h1c6/* 454*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_chanxy_config[8'hdd/* 221*/:8'hdd/* 221*/];
  assign T1644 = T1645;
  assign T1645 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_chanxy_config[8'hde/* 222*/:8'hde/* 222*/];
  assign T1652 = T1653;
  assign T1653 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_chanxy_config[8'hdf/* 223*/:8'hdf/* 223*/];
  assign T1660 = T1661;
  assign T1661 = io_chanxy_in[9'h1cd/* 461*/:9'h1cc/* 460*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_chanxy_config[8'he0/* 224*/:8'he0/* 224*/];
  assign T1668 = T1669;
  assign T1669 = io_chanxy_in[9'h1cf/* 463*/:9'h1ce/* 462*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_chanxy_config[8'he1/* 225*/:8'he1/* 225*/];
  assign T1676 = T1677;
  assign T1677 = io_chanxy_in[9'h1d1/* 465*/:9'h1d0/* 464*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_chanxy_config[8'he5/* 229*/:8'he2/* 226*/];
  assign T1684 = T1685;
  assign T1685 = io_chanxy_in[9'h1db/* 475*/:9'h1d2/* 466*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_chanxy_config[8'he7/* 231*/:8'he6/* 230*/];
  assign T1692 = T1693;
  assign T1693 = io_chanxy_in[9'h1de/* 478*/:9'h1dc/* 476*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_chanxy_config[8'heb/* 235*/:8'he8/* 232*/];
  assign T1700 = T1701;
  assign T1701 = io_chanxy_in[9'h1e8/* 488*/:9'h1df/* 479*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_chanxy_config[8'hed/* 237*/:8'hec/* 236*/];
  assign T1708 = T1709;
  assign T1709 = io_chanxy_in[9'h1eb/* 491*/:9'h1e9/* 489*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_chanxy_config[8'hf1/* 241*/:8'hee/* 238*/];
  assign T1716 = T1717;
  assign T1717 = io_chanxy_in[9'h1f5/* 501*/:9'h1ec/* 492*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1724 = T1725;
  assign T1725 = io_chanxy_in[9'h1f7/* 503*/:9'h1f6/* 502*/];
  assign T1726 = T1727;
  assign T1727 = T1728;
  assign T1728 = T1732[T1729];
  assign T1729 = T1730;
  assign T1730 = T1731;
  assign T1731 = io_chanxy_config[8'hf6/* 246*/:8'hf3/* 243*/];
  assign T1732 = T1733;
  assign T1733 = io_chanxy_in[10'h201/* 513*/:9'h1f8/* 504*/];
  assign T1734 = T1735;
  assign T1735 = T1736;
  assign T1736 = T1740[T1737];
  assign T1737 = T1738;
  assign T1738 = T1739;
  assign T1739 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T1740 = T1741;
  assign T1741 = io_chanxy_in[10'h203/* 515*/:10'h202/* 514*/];
  assign T1742 = T1743;
  assign T1743 = T1744;
  assign T1744 = T1748[T1745];
  assign T1745 = T1746;
  assign T1746 = T1747;
  assign T1747 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T1748 = T1749;
  assign T1749 = io_chanxy_in[10'h20d/* 525*/:10'h204/* 516*/];
  assign T1750 = T1751;
  assign T1751 = T1752;
  assign T1752 = T1756[T1753];
  assign T1753 = T1754;
  assign T1754 = T1755;
  assign T1755 = io_chanxy_config[8'hfc/* 252*/:8'hfc/* 252*/];
  assign T1756 = T1757;
  assign T1757 = io_chanxy_in[10'h20f/* 527*/:10'h20e/* 526*/];
  assign T1758 = T1759;
  assign T1759 = T1760;
  assign T1760 = T1764[T1761];
  assign T1761 = T1762;
  assign T1762 = T1763;
  assign T1763 = io_chanxy_config[9'h100/* 256*/:8'hfd/* 253*/];
  assign T1764 = T1765;
  assign T1765 = io_chanxy_in[10'h219/* 537*/:10'h210/* 528*/];
  assign T1766 = T1767;
  assign T1767 = T1768;
  assign T1768 = T1772[T1769];
  assign T1769 = T1770;
  assign T1770 = T1771;
  assign T1771 = io_chanxy_config[9'h101/* 257*/:9'h101/* 257*/];
  assign T1772 = T1773;
  assign T1773 = io_chanxy_in[10'h21b/* 539*/:10'h21a/* 538*/];
  assign T1774 = T1775;
  assign T1775 = T1776;
  assign T1776 = T1780[T1777];
  assign T1777 = T1778;
  assign T1778 = T1779;
  assign T1779 = io_chanxy_config[9'h105/* 261*/:9'h102/* 258*/];
  assign T1780 = T1781;
  assign T1781 = io_chanxy_in[10'h225/* 549*/:10'h21c/* 540*/];
  assign T1782 = T1783;
  assign T1783 = T1784;
  assign T1784 = T1788[T1785];
  assign T1785 = T1786;
  assign T1786 = T1787;
  assign T1787 = io_chanxy_config[9'h106/* 262*/:9'h106/* 262*/];
  assign T1788 = T1789;
  assign T1789 = io_chanxy_in[10'h227/* 551*/:10'h226/* 550*/];
  assign T1790 = T1791;
  assign T1791 = T1792;
  assign T1792 = T1796[T1793];
  assign T1793 = T1794;
  assign T1794 = T1795;
  assign T1795 = io_chanxy_config[9'h10a/* 266*/:9'h107/* 263*/];
  assign T1796 = T1797;
  assign T1797 = io_chanxy_in[10'h231/* 561*/:10'h228/* 552*/];
  assign T1798 = T1799;
  assign T1799 = T1800;
  assign T1800 = T1804[T1801];
  assign T1801 = T1802;
  assign T1802 = T1803;
  assign T1803 = io_chanxy_config[9'h10b/* 267*/:9'h10b/* 267*/];
  assign T1804 = T1805;
  assign T1805 = io_chanxy_in[10'h233/* 563*/:10'h232/* 562*/];
  assign T1806 = T1807;
  assign T1807 = T1808;
  assign T1808 = T1812[T1809];
  assign T1809 = T1810;
  assign T1810 = T1811;
  assign T1811 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1812 = T1813;
  assign T1813 = io_chanxy_in[10'h23c/* 572*/:10'h234/* 564*/];
  assign T1814 = T1815;
  assign T1815 = T1816;
  assign T1816 = T1820[T1817];
  assign T1817 = T1818;
  assign T1818 = T1819;
  assign T1819 = io_chanxy_config[9'h110/* 272*/:9'h110/* 272*/];
  assign T1820 = T1821;
  assign T1821 = io_chanxy_in[10'h23e/* 574*/:10'h23d/* 573*/];
  assign T1822 = T1823;
  assign T1823 = T1824;
  assign T1824 = T1828[T1825];
  assign T1825 = T1826;
  assign T1826 = T1827;
  assign T1827 = io_chanxy_config[9'h114/* 276*/:9'h111/* 273*/];
  assign T1828 = T1829;
  assign T1829 = io_chanxy_in[10'h247/* 583*/:10'h23f/* 575*/];
  assign T1830 = T1831;
  assign T1831 = T1832;
  assign T1832 = T1836[T1833];
  assign T1833 = T1834;
  assign T1834 = T1835;
  assign T1835 = io_chanxy_config[9'h115/* 277*/:9'h115/* 277*/];
  assign T1836 = T1837;
  assign T1837 = io_chanxy_in[10'h249/* 585*/:10'h248/* 584*/];
  assign T1838 = T1839;
  assign T1839 = T1840;
  assign T1840 = T1844[T1841];
  assign T1841 = T1842;
  assign T1842 = T1843;
  assign T1843 = io_chanxy_config[9'h119/* 281*/:9'h116/* 278*/];
  assign T1844 = T1845;
  assign T1845 = io_chanxy_in[10'h252/* 594*/:10'h24a/* 586*/];
  assign T1846 = T1847;
  assign T1847 = T1848;
  assign T1848 = T1852[T1849];
  assign T1849 = T1850;
  assign T1850 = T1851;
  assign T1851 = io_chanxy_config[9'h11a/* 282*/:9'h11a/* 282*/];
  assign T1852 = T1853;
  assign T1853 = io_chanxy_in[10'h254/* 596*/:10'h253/* 595*/];
  assign T1854 = T1855;
  assign T1855 = T1856;
  assign T1856 = T1860[T1857];
  assign T1857 = T1858;
  assign T1858 = T1859;
  assign T1859 = io_chanxy_config[9'h11e/* 286*/:9'h11b/* 283*/];
  assign T1860 = T1861;
  assign T1861 = io_chanxy_in[10'h25d/* 605*/:10'h255/* 597*/];
  assign T1862 = T1863;
  assign T1863 = T1864;
  assign T1864 = T1868[T1865];
  assign T1865 = T1866;
  assign T1866 = T1867;
  assign T1867 = io_chanxy_config[9'h11f/* 287*/:9'h11f/* 287*/];
  assign T1868 = T1869;
  assign T1869 = io_chanxy_in[10'h25f/* 607*/:10'h25e/* 606*/];
  assign T1870 = T1871;
  assign T1871 = T1872;
  assign T1872 = T1876[T1873];
  assign T1873 = T1874;
  assign T1874 = T1875;
  assign T1875 = io_chanxy_config[9'h123/* 291*/:9'h120/* 288*/];
  assign T1876 = T1877;
  assign T1877 = io_chanxy_in[10'h268/* 616*/:10'h260/* 608*/];
  assign T1878 = T1879;
  assign T1879 = T1880;
  assign T1880 = T1884[T1881];
  assign T1881 = T1882;
  assign T1882 = T1883;
  assign T1883 = io_chanxy_config[9'h124/* 292*/:9'h124/* 292*/];
  assign T1884 = T1885;
  assign T1885 = io_chanxy_in[10'h26a/* 618*/:10'h269/* 617*/];
  assign T1886 = T1887;
  assign T1887 = T1888;
  assign T1888 = T1892[T1889];
  assign T1889 = T1890;
  assign T1890 = T1891;
  assign T1891 = io_chanxy_config[9'h128/* 296*/:9'h125/* 293*/];
  assign T1892 = T1893;
  assign T1893 = io_chanxy_in[10'h273/* 627*/:10'h26b/* 619*/];
  assign T1894 = T1895;
  assign T1895 = T1896;
  assign T1896 = T1900[T1897];
  assign T1897 = T1898;
  assign T1898 = T1899;
  assign T1899 = io_chanxy_config[9'h129/* 297*/:9'h129/* 297*/];
  assign T1900 = T1901;
  assign T1901 = io_chanxy_in[10'h275/* 629*/:10'h274/* 628*/];
  assign T1902 = T1903;
  assign T1903 = T1904;
  assign T1904 = T1908[T1905];
  assign T1905 = T1906;
  assign T1906 = T1907;
  assign T1907 = io_chanxy_config[9'h12d/* 301*/:9'h12a/* 298*/];
  assign T1908 = T1909;
  assign T1909 = io_chanxy_in[10'h27e/* 638*/:10'h276/* 630*/];
  assign T1910 = T1911;
  assign T1911 = T1912;
  assign T1912 = T1916[T1913];
  assign T1913 = T1914;
  assign T1914 = T1915;
  assign T1915 = io_chanxy_config[9'h12e/* 302*/:9'h12e/* 302*/];
  assign T1916 = T1917;
  assign T1917 = io_chanxy_in[10'h280/* 640*/:10'h27f/* 639*/];
  assign T1918 = T1919;
  assign T1919 = T1920;
  assign T1920 = T1924[T1921];
  assign T1921 = T1922;
  assign T1922 = T1923;
  assign T1923 = io_chanxy_config[9'h132/* 306*/:9'h12f/* 303*/];
  assign T1924 = T1925;
  assign T1925 = io_chanxy_in[10'h289/* 649*/:10'h281/* 641*/];
  assign T1926 = T1927;
  assign T1927 = T1928;
  assign T1928 = T1932[T1929];
  assign T1929 = T1930;
  assign T1930 = T1931;
  assign T1931 = io_chanxy_config[9'h133/* 307*/:9'h133/* 307*/];
  assign T1932 = T1933;
  assign T1933 = io_chanxy_in[10'h28b/* 651*/:10'h28a/* 650*/];
  assign T1934 = T1935;
  assign T1935 = T1936;
  assign T1936 = T1940[T1937];
  assign T1937 = T1938;
  assign T1938 = T1939;
  assign T1939 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1940 = T1941;
  assign T1941 = io_chanxy_in[10'h294/* 660*/:10'h28c/* 652*/];
  assign T1942 = T1943;
  assign T1943 = T1944;
  assign T1944 = T1948[T1945];
  assign T1945 = T1946;
  assign T1946 = T1947;
  assign T1947 = io_chanxy_config[9'h138/* 312*/:9'h138/* 312*/];
  assign T1948 = T1949;
  assign T1949 = io_chanxy_in[10'h296/* 662*/:10'h295/* 661*/];
  assign T1950 = T1951;
  assign T1951 = T1952;
  assign T1952 = T1956[T1953];
  assign T1953 = T1954;
  assign T1954 = T1955;
  assign T1955 = io_chanxy_config[9'h13c/* 316*/:9'h139/* 313*/];
  assign T1956 = T1957;
  assign T1957 = io_chanxy_in[10'h29f/* 671*/:10'h297/* 663*/];
  assign T1958 = T1959;
  assign T1959 = T1960;
  assign T1960 = T1964[T1961];
  assign T1961 = T1962;
  assign T1962 = T1963;
  assign T1963 = io_chanxy_config[9'h13d/* 317*/:9'h13d/* 317*/];
  assign T1964 = T1965;
  assign T1965 = io_chanxy_in[10'h2a1/* 673*/:10'h2a0/* 672*/];
  assign T1966 = T1967;
  assign T1967 = T1968;
  assign T1968 = T1972[T1969];
  assign T1969 = T1970;
  assign T1970 = T1971;
  assign T1971 = io_chanxy_config[9'h141/* 321*/:9'h13e/* 318*/];
  assign T1972 = T1973;
  assign T1973 = io_chanxy_in[10'h2aa/* 682*/:10'h2a2/* 674*/];
  assign T1974 = T1975;
  assign T1975 = T1976;
  assign T1976 = T1980[T1977];
  assign T1977 = T1978;
  assign T1978 = T1979;
  assign T1979 = io_chanxy_config[9'h142/* 322*/:9'h142/* 322*/];
  assign T1980 = T1981;
  assign T1981 = io_chanxy_in[10'h2ac/* 684*/:10'h2ab/* 683*/];
  assign T1982 = T1983;
  assign T1983 = T1984;
  assign T1984 = T1988[T1985];
  assign T1985 = T1986;
  assign T1986 = T1987;
  assign T1987 = io_chanxy_config[9'h146/* 326*/:9'h143/* 323*/];
  assign T1988 = T1989;
  assign T1989 = io_chanxy_in[10'h2b5/* 693*/:10'h2ad/* 685*/];
  assign T1990 = T1991;
  assign T1991 = T1992;
  assign T1992 = T1996[T1993];
  assign T1993 = T1994;
  assign T1994 = T1995;
  assign T1995 = io_chanxy_config[9'h147/* 327*/:9'h147/* 327*/];
  assign T1996 = T1997;
  assign T1997 = io_chanxy_in[10'h2b7/* 695*/:10'h2b6/* 694*/];
  assign io_ipin_out = T1998;
  assign T1998 = T1999;
  assign T1999 = {T2318, T2000};
  assign T2000 = T2001;
  assign T2001 = {T2310, T2002};
  assign T2002 = T2003;
  assign T2003 = {T2302, T2004};
  assign T2004 = T2005;
  assign T2005 = {T2294, T2006};
  assign T2006 = T2007;
  assign T2007 = {T2286, T2008};
  assign T2008 = T2009;
  assign T2009 = {T2278, T2010};
  assign T2010 = T2011;
  assign T2011 = {T2270, T2012};
  assign T2012 = T2013;
  assign T2013 = {T2262, T2014};
  assign T2014 = T2015;
  assign T2015 = {T2254, T2016};
  assign T2016 = T2017;
  assign T2017 = {T2246, T2018};
  assign T2018 = T2019;
  assign T2019 = {T2238, T2020};
  assign T2020 = T2021;
  assign T2021 = {T2230, T2022};
  assign T2022 = T2023;
  assign T2023 = {T2222, T2024};
  assign T2024 = T2025;
  assign T2025 = {T2214, T2026};
  assign T2026 = T2027;
  assign T2027 = {T2206, T2028};
  assign T2028 = T2029;
  assign T2029 = {T2198, T2030};
  assign T2030 = T2031;
  assign T2031 = {T2190, T2032};
  assign T2032 = T2033;
  assign T2033 = {T2182, T2034};
  assign T2034 = T2035;
  assign T2035 = {T2174, T2036};
  assign T2036 = T2037;
  assign T2037 = {T2166, T2038};
  assign T2038 = T2039;
  assign T2039 = {T2158, T2040};
  assign T2040 = T2041;
  assign T2041 = {T2150, T2042};
  assign T2042 = T2043;
  assign T2043 = {T2142, T2044};
  assign T2044 = T2045;
  assign T2045 = {T2134, T2046};
  assign T2046 = T2047;
  assign T2047 = {T2126, T2048};
  assign T2048 = T2049;
  assign T2049 = {T2118, T2050};
  assign T2050 = T2051;
  assign T2051 = {T2110, T2052};
  assign T2052 = T2053;
  assign T2053 = {T2102, T2054};
  assign T2054 = T2055;
  assign T2055 = {T2094, T2056};
  assign T2056 = T2057;
  assign T2057 = {T2086, T2058};
  assign T2058 = T2059;
  assign T2059 = {T2078, T2060};
  assign T2060 = T2061;
  assign T2061 = {T2070, T2062};
  assign T2062 = T2063;
  assign T2063 = T2064;
  assign T2064 = T2068[T2065];
  assign T2065 = T2066;
  assign T2066 = T2067;
  assign T2067 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T2068 = T2069;
  assign T2069 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T2070 = T2071;
  assign T2071 = T2072;
  assign T2072 = T2076[T2073];
  assign T2073 = T2074;
  assign T2074 = T2075;
  assign T2075 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T2076 = T2077;
  assign T2077 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T2078 = T2079;
  assign T2079 = T2080;
  assign T2080 = T2084[T2081];
  assign T2081 = T2082;
  assign T2082 = T2083;
  assign T2083 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T2084 = T2085;
  assign T2085 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T2086 = T2087;
  assign T2087 = T2088;
  assign T2088 = T2092[T2089];
  assign T2089 = T2090;
  assign T2090 = T2091;
  assign T2091 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T2092 = T2093;
  assign T2093 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T2094 = T2095;
  assign T2095 = T2096;
  assign T2096 = T2100[T2097];
  assign T2097 = T2098;
  assign T2098 = T2099;
  assign T2099 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T2100 = T2101;
  assign T2101 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T2102 = T2103;
  assign T2103 = T2104;
  assign T2104 = T2108[T2105];
  assign T2105 = T2106;
  assign T2106 = T2107;
  assign T2107 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T2108 = T2109;
  assign T2109 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T2110 = T2111;
  assign T2111 = T2112;
  assign T2112 = T2116[T2113];
  assign T2113 = T2114;
  assign T2114 = T2115;
  assign T2115 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T2116 = T2117;
  assign T2117 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T2118 = T2119;
  assign T2119 = T2120;
  assign T2120 = T2124[T2121];
  assign T2121 = T2122;
  assign T2122 = T2123;
  assign T2123 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T2124 = T2125;
  assign T2125 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T2126 = T2127;
  assign T2127 = T2128;
  assign T2128 = T2132[T2129];
  assign T2129 = T2130;
  assign T2130 = T2131;
  assign T2131 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T2132 = T2133;
  assign T2133 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T2134 = T2135;
  assign T2135 = T2136;
  assign T2136 = T2140[T2137];
  assign T2137 = T2138;
  assign T2138 = T2139;
  assign T2139 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T2140 = T2141;
  assign T2141 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T2142 = T2143;
  assign T2143 = T2144;
  assign T2144 = T2148[T2145];
  assign T2145 = T2146;
  assign T2146 = T2147;
  assign T2147 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T2148 = T2149;
  assign T2149 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T2150 = T2151;
  assign T2151 = T2152;
  assign T2152 = T2156[T2153];
  assign T2153 = T2154;
  assign T2154 = T2155;
  assign T2155 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T2156 = T2157;
  assign T2157 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T2158 = T2159;
  assign T2159 = T2160;
  assign T2160 = T2164[T2161];
  assign T2161 = T2162;
  assign T2162 = T2163;
  assign T2163 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T2164 = T2165;
  assign T2165 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T2166 = T2167;
  assign T2167 = T2168;
  assign T2168 = T2172[T2169];
  assign T2169 = T2170;
  assign T2170 = T2171;
  assign T2171 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T2172 = T2173;
  assign T2173 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T2174 = T2175;
  assign T2175 = T2176;
  assign T2176 = T2180[T2177];
  assign T2177 = T2178;
  assign T2178 = T2179;
  assign T2179 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T2180 = T2181;
  assign T2181 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T2182 = T2183;
  assign T2183 = T2184;
  assign T2184 = T2188[T2185];
  assign T2185 = T2186;
  assign T2186 = T2187;
  assign T2187 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T2188 = T2189;
  assign T2189 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T2190 = T2191;
  assign T2191 = T2192;
  assign T2192 = T2196[T2193];
  assign T2193 = T2194;
  assign T2194 = T2195;
  assign T2195 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T2196 = T2197;
  assign T2197 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T2198 = T2199;
  assign T2199 = T2200;
  assign T2200 = T2204[T2201];
  assign T2201 = T2202;
  assign T2202 = T2203;
  assign T2203 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T2204 = T2205;
  assign T2205 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T2206 = T2207;
  assign T2207 = T2208;
  assign T2208 = T2212[T2209];
  assign T2209 = T2210;
  assign T2210 = T2211;
  assign T2211 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T2212 = T2213;
  assign T2213 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T2214 = T2215;
  assign T2215 = T2216;
  assign T2216 = T2220[T2217];
  assign T2217 = T2218;
  assign T2218 = T2219;
  assign T2219 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T2220 = T2221;
  assign T2221 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T2222 = T2223;
  assign T2223 = T2224;
  assign T2224 = T2228[T2225];
  assign T2225 = T2226;
  assign T2226 = T2227;
  assign T2227 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T2228 = T2229;
  assign T2229 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T2230 = T2231;
  assign T2231 = T2232;
  assign T2232 = T2236[T2233];
  assign T2233 = T2234;
  assign T2234 = T2235;
  assign T2235 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T2236 = T2237;
  assign T2237 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T2238 = T2239;
  assign T2239 = T2240;
  assign T2240 = T2244[T2241];
  assign T2241 = T2242;
  assign T2242 = T2243;
  assign T2243 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T2244 = T2245;
  assign T2245 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T2246 = T2247;
  assign T2247 = T2248;
  assign T2248 = T2252[T2249];
  assign T2249 = T2250;
  assign T2250 = T2251;
  assign T2251 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T2252 = T2253;
  assign T2253 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T2254 = T2255;
  assign T2255 = T2256;
  assign T2256 = T2260[T2257];
  assign T2257 = T2258;
  assign T2258 = T2259;
  assign T2259 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T2260 = T2261;
  assign T2261 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T2262 = T2263;
  assign T2263 = T2264;
  assign T2264 = T2268[T2265];
  assign T2265 = T2266;
  assign T2266 = T2267;
  assign T2267 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T2268 = T2269;
  assign T2269 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T2270 = T2271;
  assign T2271 = T2272;
  assign T2272 = T2276[T2273];
  assign T2273 = T2274;
  assign T2274 = T2275;
  assign T2275 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T2276 = T2277;
  assign T2277 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T2278 = T2279;
  assign T2279 = T2280;
  assign T2280 = T2284[T2281];
  assign T2281 = T2282;
  assign T2282 = T2283;
  assign T2283 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T2284 = T2285;
  assign T2285 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T2286 = T2287;
  assign T2287 = T2288;
  assign T2288 = T2292[T2289];
  assign T2289 = T2290;
  assign T2290 = T2291;
  assign T2291 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T2292 = T2293;
  assign T2293 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T2294 = T2295;
  assign T2295 = T2296;
  assign T2296 = T2300[T2297];
  assign T2297 = T2298;
  assign T2298 = T2299;
  assign T2299 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T2300 = T2301;
  assign T2301 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T2302 = T2303;
  assign T2303 = T2304;
  assign T2304 = T2308[T2305];
  assign T2305 = T2306;
  assign T2306 = T2307;
  assign T2307 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T2308 = T2309;
  assign T2309 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T2310 = T2311;
  assign T2311 = T2312;
  assign T2312 = T2316[T2313];
  assign T2313 = T2314;
  assign T2314 = T2315;
  assign T2315 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T2316 = T2317;
  assign T2317 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T2318 = T2319;
  assign T2319 = T2320;
  assign T2320 = T2324[T2321];
  assign T2321 = T2322;
  assign T2322 = T2323;
  assign T2323 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T2324 = T2325;
  assign T2325 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_9(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [45:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [695:0] io_chanxy_in,
    output[199:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[327:0] T0;
  wire[1471:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[199:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5bd/* 1469*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_46 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_7 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_8(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[10:0] T284;
  wire[10:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[10:0] T292;
  wire[10:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[10:0] T300;
  wire[10:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[10:0] T308;
  wire[10:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[10:0] T316;
  wire[10:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[10:0] T324;
  wire[10:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[10:0] T332;
  wire[10:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[10:0] T340;
  wire[10:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[10:0] T348;
  wire[10:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[10:0] T356;
  wire[10:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[10:0] T364;
  wire[10:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[10:0] T372;
  wire[10:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[10:0] T380;
  wire[10:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[10:0] T388;
  wire[10:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[10:0] T396;
  wire[10:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[10:0] T404;
  wire[10:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[10:0] T412;
  wire[10:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[10:0] T420;
  wire[10:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[10:0] T428;
  wire[10:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[3:0] T433;
  wire[3:0] T434;
  wire[3:0] T435;
  wire[10:0] T436;
  wire[10:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[3:0] T441;
  wire[3:0] T442;
  wire[3:0] T443;
  wire[10:0] T444;
  wire[10:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[3:0] T449;
  wire[3:0] T450;
  wire[3:0] T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[10:0] T460;
  wire[10:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[10:0] T468;
  wire[10:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[3:0] T473;
  wire[3:0] T474;
  wire[3:0] T475;
  wire[10:0] T476;
  wire[10:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[3:0] T481;
  wire[3:0] T482;
  wire[3:0] T483;
  wire[10:0] T484;
  wire[10:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[10:0] T492;
  wire[10:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[10:0] T500;
  wire[10:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[10:0] T508;
  wire[10:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[10:0] T516;
  wire[10:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[3:0] T521;
  wire[3:0] T522;
  wire[3:0] T523;
  wire[10:0] T524;
  wire[10:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[10:0] T532;
  wire[10:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[10:0] T540;
  wire[10:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[10:0] T548;
  wire[10:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[3:0] T553;
  wire[3:0] T554;
  wire[3:0] T555;
  wire[10:0] T556;
  wire[10:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[3:0] T561;
  wire[3:0] T562;
  wire[3:0] T563;
  wire[10:0] T564;
  wire[10:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[3:0] T569;
  wire[3:0] T570;
  wire[3:0] T571;
  wire[10:0] T572;
  wire[10:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[10:0] T580;
  wire[10:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[10:0] T588;
  wire[10:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[3:0] T593;
  wire[3:0] T594;
  wire[3:0] T595;
  wire[10:0] T596;
  wire[10:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[3:0] T633;
  wire[3:0] T634;
  wire[3:0] T635;
  wire[10:0] T636;
  wire[10:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[3:0] T673;
  wire[3:0] T674;
  wire[3:0] T675;
  wire[10:0] T676;
  wire[10:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire[1:0] T683;
  wire[2:0] T684;
  wire[2:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[1:0] T689;
  wire[1:0] T690;
  wire[1:0] T691;
  wire[2:0] T692;
  wire[2:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[1:0] T697;
  wire[1:0] T698;
  wire[1:0] T699;
  wire[2:0] T700;
  wire[2:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[1:0] T705;
  wire[1:0] T706;
  wire[1:0] T707;
  wire[2:0] T708;
  wire[2:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[3:0] T713;
  wire[3:0] T714;
  wire[3:0] T715;
  wire[10:0] T716;
  wire[10:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[2:0] T724;
  wire[2:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[1:0] T729;
  wire[1:0] T730;
  wire[1:0] T731;
  wire[2:0] T732;
  wire[2:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[1:0] T737;
  wire[1:0] T738;
  wire[1:0] T739;
  wire[2:0] T740;
  wire[2:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[1:0] T745;
  wire[1:0] T746;
  wire[1:0] T747;
  wire[2:0] T748;
  wire[2:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[3:0] T753;
  wire[3:0] T754;
  wire[3:0] T755;
  wire[10:0] T756;
  wire[10:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[1:0] T777;
  wire[1:0] T778;
  wire[1:0] T779;
  wire[2:0] T780;
  wire[2:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[3:0] T793;
  wire[3:0] T794;
  wire[3:0] T795;
  wire[10:0] T796;
  wire[10:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire[1:0] T801;
  wire[1:0] T802;
  wire[1:0] T803;
  wire[2:0] T804;
  wire[2:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[1:0] T809;
  wire[1:0] T810;
  wire[1:0] T811;
  wire[2:0] T812;
  wire[2:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[1:0] T817;
  wire[1:0] T818;
  wire[1:0] T819;
  wire[2:0] T820;
  wire[2:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[1:0] T825;
  wire[1:0] T826;
  wire[1:0] T827;
  wire[2:0] T828;
  wire[2:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[3:0] T833;
  wire[3:0] T834;
  wire[3:0] T835;
  wire[10:0] T836;
  wire[10:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[1:0] T841;
  wire[1:0] T842;
  wire[1:0] T843;
  wire[2:0] T844;
  wire[2:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire[1:0] T849;
  wire[1:0] T850;
  wire[1:0] T851;
  wire[2:0] T852;
  wire[2:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[1:0] T857;
  wire[1:0] T858;
  wire[1:0] T859;
  wire[2:0] T860;
  wire[2:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[1:0] T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[2:0] T868;
  wire[2:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[3:0] T873;
  wire[3:0] T874;
  wire[3:0] T875;
  wire[10:0] T876;
  wire[10:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[1:0] T881;
  wire[1:0] T882;
  wire[1:0] T883;
  wire[2:0] T884;
  wire[2:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[1:0] T889;
  wire[1:0] T890;
  wire[1:0] T891;
  wire[2:0] T892;
  wire[2:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[1:0] T897;
  wire[1:0] T898;
  wire[1:0] T899;
  wire[2:0] T900;
  wire[2:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[1:0] T905;
  wire[1:0] T906;
  wire[1:0] T907;
  wire[2:0] T908;
  wire[2:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[3:0] T913;
  wire[3:0] T914;
  wire[3:0] T915;
  wire[10:0] T916;
  wire[10:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire[1:0] T922;
  wire[1:0] T923;
  wire[2:0] T924;
  wire[2:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[2:0] T932;
  wire[2:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[1:0] T937;
  wire[1:0] T938;
  wire[1:0] T939;
  wire[2:0] T940;
  wire[2:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[1:0] T945;
  wire[1:0] T946;
  wire[1:0] T947;
  wire[2:0] T948;
  wire[2:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[3:0] T953;
  wire[3:0] T954;
  wire[3:0] T955;
  wire[10:0] T956;
  wire[10:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[1:0] T961;
  wire[1:0] T962;
  wire[1:0] T963;
  wire[2:0] T964;
  wire[2:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[1:0] T969;
  wire[1:0] T970;
  wire[1:0] T971;
  wire[2:0] T972;
  wire[2:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[1:0] T977;
  wire[1:0] T978;
  wire[1:0] T979;
  wire[2:0] T980;
  wire[2:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[1:0] T985;
  wire[1:0] T986;
  wire[1:0] T987;
  wire[2:0] T988;
  wire[2:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[3:0] T993;
  wire[3:0] T994;
  wire[3:0] T995;
  wire[10:0] T996;
  wire[10:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire[3:0] T1033;
  wire[3:0] T1034;
  wire[3:0] T1035;
  wire[10:0] T1036;
  wire[10:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire[3:0] T1073;
  wire[3:0] T1074;
  wire[3:0] T1075;
  wire[10:0] T1076;
  wire[10:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire[1:0] T1092;
  wire[1:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[1:0] T1108;
  wire[1:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[10:0] T1116;
  wire[10:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire[1:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire[1:0] T1140;
  wire[1:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire[1:0] T1148;
  wire[1:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[3:0] T1153;
  wire[3:0] T1154;
  wire[3:0] T1155;
  wire[10:0] T1156;
  wire[10:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire[1:0] T1172;
  wire[1:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire[1:0] T1188;
  wire[1:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[10:0] T1196;
  wire[10:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire[1:0] T1204;
  wire[1:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire T1211;
  wire[1:0] T1212;
  wire[1:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire[1:0] T1220;
  wire[1:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire[1:0] T1228;
  wire[1:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[3:0] T1233;
  wire[3:0] T1234;
  wire[3:0] T1235;
  wire[10:0] T1236;
  wire[10:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire[1:0] T1244;
  wire[1:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[1:0] T1252;
  wire[1:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire[1:0] T1260;
  wire[1:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[1:0] T1268;
  wire[1:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[10:0] T1276;
  wire[10:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire[1:0] T1292;
  wire[1:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire[1:0] T1308;
  wire[1:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire[3:0] T1313;
  wire[3:0] T1314;
  wire[3:0] T1315;
  wire[10:0] T1316;
  wire[10:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire[1:0] T1340;
  wire[1:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[10:0] T1356;
  wire[10:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire[1:0] T1364;
  wire[1:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire[1:0] T1372;
  wire[1:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire[1:0] T1380;
  wire[1:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire[1:0] T1388;
  wire[1:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire[3:0] T1393;
  wire[3:0] T1394;
  wire[3:0] T1395;
  wire[10:0] T1396;
  wire[10:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h6d/* 109*/:7'h63/* 99*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h78/* 120*/:7'h6e/* 110*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[8'h83/* 131*/:7'h79/* 121*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[8'h8e/* 142*/:8'h84/* 132*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[8'h99/* 153*/:8'h8f/* 143*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[8'ha4/* 164*/:8'h9a/* 154*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[8'haf/* 175*/:8'ha5/* 165*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[8'hba/* 186*/:8'hb0/* 176*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[8'hc5/* 197*/:8'hbb/* 187*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[8'hd0/* 208*/:8'hc6/* 198*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[8'hdb/* 219*/:8'hd1/* 209*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[8'he6/* 230*/:8'hdc/* 220*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[8'hf1/* 241*/:8'he7/* 231*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[8'hfc/* 252*/:8'hf2/* 242*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[9'h107/* 263*/:8'hfd/* 253*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[9'h112/* 274*/:9'h108/* 264*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[9'h11d/* 285*/:9'h113/* 275*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[9'h128/* 296*/:9'h11e/* 286*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[9'h133/* 307*/:9'h129/* 297*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[9'h13e/* 318*/:9'h134/* 308*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[9'h149/* 329*/:9'h13f/* 319*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[9'h154/* 340*/:9'h14a/* 330*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[9'h15f/* 351*/:9'h155/* 341*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[9'h16a/* 362*/:9'h160/* 352*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[9'h175/* 373*/:9'h16b/* 363*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[9'h180/* 384*/:9'h176/* 374*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[9'h18b/* 395*/:9'h181/* 385*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[9'h196/* 406*/:9'h18c/* 396*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[9'h1ac/* 428*/:9'h1a2/* 418*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[9'h1b7/* 439*/:9'h1ad/* 429*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[9'h1ba/* 442*/:9'h1b8/* 440*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[9'h1bd/* 445*/:9'h1bb/* 443*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[9'h1c0/* 448*/:9'h1be/* 446*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[9'h1c3/* 451*/:9'h1c1/* 449*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[8'hab/* 171*/:8'ha8/* 168*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[9'h1ce/* 462*/:9'h1c4/* 452*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[9'h1d1/* 465*/:9'h1cf/* 463*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[9'h1d4/* 468*/:9'h1d2/* 466*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[9'h1d7/* 471*/:9'h1d5/* 469*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[9'h1da/* 474*/:9'h1d8/* 472*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[8'hb7/* 183*/:8'hb4/* 180*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[9'h1e5/* 485*/:9'h1db/* 475*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[9'h1e8/* 488*/:9'h1e6/* 486*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[8'hbb/* 187*/:8'hba/* 186*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[9'h1eb/* 491*/:9'h1e9/* 489*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[8'hbd/* 189*/:8'hbc/* 188*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[9'h1ee/* 494*/:9'h1ec/* 492*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[9'h1f1/* 497*/:9'h1ef/* 495*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[8'hc3/* 195*/:8'hc0/* 192*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[9'h1fc/* 508*/:9'h1f2/* 498*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[9'h1ff/* 511*/:9'h1fd/* 509*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[10'h202/* 514*/:10'h200/* 512*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[10'h205/* 517*/:10'h203/* 515*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[10'h208/* 520*/:10'h206/* 518*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'hcf/* 207*/:8'hcc/* 204*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[10'h213/* 531*/:10'h209/* 521*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[10'h216/* 534*/:10'h214/* 532*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[10'h219/* 537*/:10'h217/* 535*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'hd5/* 213*/:8'hd4/* 212*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[10'h21c/* 540*/:10'h21a/* 538*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'hd7/* 215*/:8'hd6/* 214*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[10'h21f/* 543*/:10'h21d/* 541*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'hdb/* 219*/:8'hd8/* 216*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[10'h22a/* 554*/:10'h220/* 544*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[10'h22d/* 557*/:10'h22b/* 555*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[10'h230/* 560*/:10'h22e/* 558*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'he1/* 225*/:8'he0/* 224*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[10'h233/* 563*/:10'h231/* 561*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'he3/* 227*/:8'he2/* 226*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[10'h236/* 566*/:10'h234/* 564*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'he7/* 231*/:8'he4/* 228*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[10'h241/* 577*/:10'h237/* 567*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'he9/* 233*/:8'he8/* 232*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[10'h244/* 580*/:10'h242/* 578*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'heb/* 235*/:8'hea/* 234*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[10'h247/* 583*/:10'h245/* 581*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'hed/* 237*/:8'hec/* 236*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[10'h24a/* 586*/:10'h248/* 584*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'hef/* 239*/:8'hee/* 238*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[10'h24d/* 589*/:10'h24b/* 587*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'hf3/* 243*/:8'hf0/* 240*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[10'h258/* 600*/:10'h24e/* 590*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'hf5/* 245*/:8'hf4/* 244*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[10'h25b/* 603*/:10'h259/* 601*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'hf7/* 247*/:8'hf6/* 246*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[10'h25e/* 606*/:10'h25c/* 604*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'hf9/* 249*/:8'hf8/* 248*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[10'h261/* 609*/:10'h25f/* 607*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[10'h264/* 612*/:10'h262/* 610*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'hff/* 255*/:8'hfc/* 252*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[10'h26f/* 623*/:10'h265/* 613*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[9'h101/* 257*/:9'h100/* 256*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[10'h272/* 626*/:10'h270/* 624*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[9'h103/* 259*/:9'h102/* 258*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[10'h275/* 629*/:10'h273/* 627*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[9'h105/* 261*/:9'h104/* 260*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[10'h278/* 632*/:10'h276/* 630*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[9'h107/* 263*/:9'h106/* 262*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[10'h27b/* 635*/:10'h279/* 633*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[9'h10b/* 267*/:9'h108/* 264*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[10'h286/* 646*/:10'h27c/* 636*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[10'h289/* 649*/:10'h287/* 647*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[10'h28c/* 652*/:10'h28a/* 650*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[9'h111/* 273*/:9'h110/* 272*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[10'h28f/* 655*/:10'h28d/* 653*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[9'h113/* 275*/:9'h112/* 274*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[10'h292/* 658*/:10'h290/* 656*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[9'h117/* 279*/:9'h114/* 276*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[10'h29d/* 669*/:10'h293/* 659*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[9'h118/* 280*/:9'h118/* 280*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[10'h29f/* 671*/:10'h29e/* 670*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[9'h119/* 281*/:9'h119/* 281*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[10'h2a1/* 673*/:10'h2a0/* 672*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[9'h11a/* 282*/:9'h11a/* 282*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[10'h2a3/* 675*/:10'h2a2/* 674*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[9'h11b/* 283*/:9'h11b/* 283*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[10'h2a5/* 677*/:10'h2a4/* 676*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[9'h11f/* 287*/:9'h11c/* 284*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[10'h2b0/* 688*/:10'h2a6/* 678*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[9'h120/* 288*/:9'h120/* 288*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[10'h2b2/* 690*/:10'h2b1/* 689*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[9'h121/* 289*/:9'h121/* 289*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[10'h2b4/* 692*/:10'h2b3/* 691*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[9'h122/* 290*/:9'h122/* 290*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[10'h2b6/* 694*/:10'h2b5/* 693*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[9'h123/* 291*/:9'h123/* 291*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[10'h2b8/* 696*/:10'h2b7/* 695*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[10'h2c3/* 707*/:10'h2b9/* 697*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[9'h128/* 296*/:9'h128/* 296*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[10'h2c5/* 709*/:10'h2c4/* 708*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[9'h129/* 297*/:9'h129/* 297*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[10'h2c7/* 711*/:10'h2c6/* 710*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[9'h12a/* 298*/:9'h12a/* 298*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[10'h2c9/* 713*/:10'h2c8/* 712*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[9'h12b/* 299*/:9'h12b/* 299*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[10'h2cb/* 715*/:10'h2ca/* 714*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[9'h12f/* 303*/:9'h12c/* 300*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[10'h2d6/* 726*/:10'h2cc/* 716*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[9'h130/* 304*/:9'h130/* 304*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[10'h2d8/* 728*/:10'h2d7/* 727*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[9'h131/* 305*/:9'h131/* 305*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[10'h2da/* 730*/:10'h2d9/* 729*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[9'h132/* 306*/:9'h132/* 306*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[10'h2dc/* 732*/:10'h2db/* 731*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[9'h133/* 307*/:9'h133/* 307*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h2de/* 734*/:10'h2dd/* 733*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[9'h137/* 311*/:9'h134/* 308*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h2e9/* 745*/:10'h2df/* 735*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[9'h138/* 312*/:9'h138/* 312*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h2eb/* 747*/:10'h2ea/* 746*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[9'h139/* 313*/:9'h139/* 313*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h2ed/* 749*/:10'h2ec/* 748*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[9'h13a/* 314*/:9'h13a/* 314*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h2ef/* 751*/:10'h2ee/* 750*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[9'h13b/* 315*/:9'h13b/* 315*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h2f1/* 753*/:10'h2f0/* 752*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h13f/* 319*/:9'h13c/* 316*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h2fc/* 764*/:10'h2f2/* 754*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h140/* 320*/:9'h140/* 320*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h2fe/* 766*/:10'h2fd/* 765*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h141/* 321*/:9'h141/* 321*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h300/* 768*/:10'h2ff/* 767*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h142/* 322*/:9'h142/* 322*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h302/* 770*/:10'h301/* 769*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h143/* 323*/:9'h143/* 323*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h304/* 772*/:10'h303/* 771*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h147/* 327*/:9'h144/* 324*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h30f/* 783*/:10'h305/* 773*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h148/* 328*/:9'h148/* 328*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h311/* 785*/:10'h310/* 784*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h313/* 787*/:10'h312/* 786*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h14a/* 330*/:9'h14a/* 330*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h315/* 789*/:10'h314/* 788*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h14b/* 331*/:9'h14b/* 331*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h317/* 791*/:10'h316/* 790*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h14f/* 335*/:9'h14c/* 332*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h322/* 802*/:10'h318/* 792*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h150/* 336*/:9'h150/* 336*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h324/* 804*/:10'h323/* 803*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h151/* 337*/:9'h151/* 337*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h326/* 806*/:10'h325/* 805*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h152/* 338*/:9'h152/* 338*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h328/* 808*/:10'h327/* 807*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h153/* 339*/:9'h153/* 339*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h32a/* 810*/:10'h329/* 809*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h335/* 821*/:10'h32b/* 811*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h337/* 823*/:10'h336/* 822*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h159/* 345*/:9'h159/* 345*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h339/* 825*/:10'h338/* 824*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h15a/* 346*/:9'h15a/* 346*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h33b/* 827*/:10'h33a/* 826*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h15b/* 347*/:9'h15b/* 347*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h33d/* 829*/:10'h33c/* 828*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h15f/* 351*/:9'h15c/* 348*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h348/* 840*/:10'h33e/* 830*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h160/* 352*/:9'h160/* 352*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h34a/* 842*/:10'h349/* 841*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h161/* 353*/:9'h161/* 353*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h34c/* 844*/:10'h34b/* 843*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h162/* 354*/:9'h162/* 354*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h34e/* 846*/:10'h34d/* 845*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h163/* 355*/:9'h163/* 355*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h350/* 848*/:10'h34f/* 847*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h164/* 356*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h351/* 849*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_10(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_8 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_9(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[10:0] T284;
  wire[10:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[10:0] T292;
  wire[10:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[10:0] T300;
  wire[10:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[10:0] T308;
  wire[10:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[10:0] T316;
  wire[10:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[10:0] T324;
  wire[10:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[10:0] T332;
  wire[10:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[10:0] T340;
  wire[10:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[10:0] T348;
  wire[10:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[10:0] T356;
  wire[10:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[10:0] T364;
  wire[10:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[10:0] T372;
  wire[10:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[10:0] T380;
  wire[10:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[10:0] T388;
  wire[10:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[10:0] T396;
  wire[10:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[10:0] T404;
  wire[10:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[10:0] T412;
  wire[10:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[10:0] T420;
  wire[10:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[10:0] T428;
  wire[10:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[3:0] T433;
  wire[3:0] T434;
  wire[3:0] T435;
  wire[10:0] T436;
  wire[10:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[3:0] T441;
  wire[3:0] T442;
  wire[3:0] T443;
  wire[10:0] T444;
  wire[10:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[3:0] T449;
  wire[3:0] T450;
  wire[3:0] T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[10:0] T460;
  wire[10:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[10:0] T468;
  wire[10:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[3:0] T473;
  wire[3:0] T474;
  wire[3:0] T475;
  wire[10:0] T476;
  wire[10:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[3:0] T481;
  wire[3:0] T482;
  wire[3:0] T483;
  wire[10:0] T484;
  wire[10:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[10:0] T492;
  wire[10:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[10:0] T500;
  wire[10:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[10:0] T508;
  wire[10:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[10:0] T516;
  wire[10:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[3:0] T521;
  wire[3:0] T522;
  wire[3:0] T523;
  wire[10:0] T524;
  wire[10:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[10:0] T532;
  wire[10:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[10:0] T540;
  wire[10:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[10:0] T548;
  wire[10:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[3:0] T553;
  wire[3:0] T554;
  wire[3:0] T555;
  wire[10:0] T556;
  wire[10:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[3:0] T561;
  wire[3:0] T562;
  wire[3:0] T563;
  wire[10:0] T564;
  wire[10:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[3:0] T569;
  wire[3:0] T570;
  wire[3:0] T571;
  wire[10:0] T572;
  wire[10:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[10:0] T580;
  wire[10:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[10:0] T588;
  wire[10:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[3:0] T593;
  wire[3:0] T594;
  wire[3:0] T595;
  wire[10:0] T596;
  wire[10:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[3:0] T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[10:0] T612;
  wire[10:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[3:0] T649;
  wire[3:0] T650;
  wire[3:0] T651;
  wire[10:0] T652;
  wire[10:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire[1:0] T683;
  wire[2:0] T684;
  wire[2:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[3:0] T689;
  wire[3:0] T690;
  wire[3:0] T691;
  wire[10:0] T692;
  wire[10:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[1:0] T697;
  wire[1:0] T698;
  wire[1:0] T699;
  wire[2:0] T700;
  wire[2:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[1:0] T705;
  wire[1:0] T706;
  wire[1:0] T707;
  wire[2:0] T708;
  wire[2:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[1:0] T713;
  wire[1:0] T714;
  wire[1:0] T715;
  wire[2:0] T716;
  wire[2:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[2:0] T724;
  wire[2:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[3:0] T729;
  wire[3:0] T730;
  wire[3:0] T731;
  wire[10:0] T732;
  wire[10:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[1:0] T737;
  wire[1:0] T738;
  wire[1:0] T739;
  wire[2:0] T740;
  wire[2:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[1:0] T745;
  wire[1:0] T746;
  wire[1:0] T747;
  wire[2:0] T748;
  wire[2:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[1:0] T753;
  wire[1:0] T754;
  wire[1:0] T755;
  wire[2:0] T756;
  wire[2:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[3:0] T769;
  wire[3:0] T770;
  wire[3:0] T771;
  wire[10:0] T772;
  wire[10:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[1:0] T777;
  wire[1:0] T778;
  wire[1:0] T779;
  wire[2:0] T780;
  wire[2:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[1:0] T793;
  wire[1:0] T794;
  wire[1:0] T795;
  wire[2:0] T796;
  wire[2:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire[1:0] T801;
  wire[1:0] T802;
  wire[1:0] T803;
  wire[2:0] T804;
  wire[2:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[3:0] T809;
  wire[3:0] T810;
  wire[3:0] T811;
  wire[10:0] T812;
  wire[10:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[1:0] T817;
  wire[1:0] T818;
  wire[1:0] T819;
  wire[2:0] T820;
  wire[2:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[1:0] T825;
  wire[1:0] T826;
  wire[1:0] T827;
  wire[2:0] T828;
  wire[2:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[1:0] T833;
  wire[1:0] T834;
  wire[1:0] T835;
  wire[2:0] T836;
  wire[2:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[1:0] T841;
  wire[1:0] T842;
  wire[1:0] T843;
  wire[2:0] T844;
  wire[2:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire[3:0] T849;
  wire[3:0] T850;
  wire[3:0] T851;
  wire[10:0] T852;
  wire[10:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[1:0] T857;
  wire[1:0] T858;
  wire[1:0] T859;
  wire[2:0] T860;
  wire[2:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[1:0] T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[2:0] T868;
  wire[2:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[1:0] T873;
  wire[1:0] T874;
  wire[1:0] T875;
  wire[2:0] T876;
  wire[2:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[1:0] T881;
  wire[1:0] T882;
  wire[1:0] T883;
  wire[2:0] T884;
  wire[2:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[3:0] T889;
  wire[3:0] T890;
  wire[3:0] T891;
  wire[10:0] T892;
  wire[10:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[1:0] T897;
  wire[1:0] T898;
  wire[1:0] T899;
  wire[2:0] T900;
  wire[2:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[1:0] T905;
  wire[1:0] T906;
  wire[1:0] T907;
  wire[2:0] T908;
  wire[2:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[1:0] T913;
  wire[1:0] T914;
  wire[1:0] T915;
  wire[2:0] T916;
  wire[2:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire[1:0] T922;
  wire[1:0] T923;
  wire[2:0] T924;
  wire[2:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[3:0] T929;
  wire[3:0] T930;
  wire[3:0] T931;
  wire[10:0] T932;
  wire[10:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[1:0] T937;
  wire[1:0] T938;
  wire[1:0] T939;
  wire[2:0] T940;
  wire[2:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[1:0] T945;
  wire[1:0] T946;
  wire[1:0] T947;
  wire[2:0] T948;
  wire[2:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[1:0] T953;
  wire[1:0] T954;
  wire[1:0] T955;
  wire[2:0] T956;
  wire[2:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[1:0] T961;
  wire[1:0] T962;
  wire[1:0] T963;
  wire[2:0] T964;
  wire[2:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[3:0] T969;
  wire[3:0] T970;
  wire[3:0] T971;
  wire[10:0] T972;
  wire[10:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[1:0] T977;
  wire[1:0] T978;
  wire[1:0] T979;
  wire[2:0] T980;
  wire[2:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[1:0] T985;
  wire[1:0] T986;
  wire[1:0] T987;
  wire[2:0] T988;
  wire[2:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[1:0] T993;
  wire[1:0] T994;
  wire[1:0] T995;
  wire[2:0] T996;
  wire[2:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire[3:0] T1009;
  wire[3:0] T1010;
  wire[3:0] T1011;
  wire[10:0] T1012;
  wire[10:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire[3:0] T1049;
  wire[3:0] T1050;
  wire[3:0] T1051;
  wire[10:0] T1052;
  wire[10:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[3:0] T1089;
  wire[3:0] T1090;
  wire[3:0] T1091;
  wire[10:0] T1092;
  wire[10:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire[1:0] T1100;
  wire[1:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[1:0] T1108;
  wire[1:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire[1:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[10:0] T1132;
  wire[10:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire[1:0] T1140;
  wire[1:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire[1:0] T1148;
  wire[1:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire[1:0] T1156;
  wire[1:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[3:0] T1169;
  wire[3:0] T1170;
  wire[3:0] T1171;
  wire[10:0] T1172;
  wire[10:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire[1:0] T1180;
  wire[1:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire[1:0] T1188;
  wire[1:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire[1:0] T1204;
  wire[1:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[10:0] T1212;
  wire[10:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire T1217;
  wire T1218;
  wire T1219;
  wire[1:0] T1220;
  wire[1:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire[1:0] T1228;
  wire[1:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire[1:0] T1236;
  wire[1:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire[1:0] T1244;
  wire[1:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire[3:0] T1249;
  wire[3:0] T1250;
  wire[3:0] T1251;
  wire[10:0] T1252;
  wire[10:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire T1257;
  wire T1258;
  wire T1259;
  wire[1:0] T1260;
  wire[1:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[1:0] T1268;
  wire[1:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[1:0] T1276;
  wire[1:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[10:0] T1292;
  wire[10:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire[1:0] T1308;
  wire[1:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire[3:0] T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[10:0] T1332;
  wire[10:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire[1:0] T1340;
  wire[1:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire[1:0] T1356;
  wire[1:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire[1:0] T1364;
  wire[1:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[10:0] T1372;
  wire[10:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire[1:0] T1380;
  wire[1:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire[1:0] T1388;
  wire[1:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[1:0] T1396;
  wire[1:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h6d/* 109*/:7'h63/* 99*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h78/* 120*/:7'h6e/* 110*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[8'h83/* 131*/:7'h79/* 121*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[8'h8e/* 142*/:8'h84/* 132*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[8'h99/* 153*/:8'h8f/* 143*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[8'ha4/* 164*/:8'h9a/* 154*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[8'haf/* 175*/:8'ha5/* 165*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[8'hba/* 186*/:8'hb0/* 176*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[8'hc5/* 197*/:8'hbb/* 187*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[8'hd0/* 208*/:8'hc6/* 198*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[8'hdb/* 219*/:8'hd1/* 209*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[8'he6/* 230*/:8'hdc/* 220*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[8'hf1/* 241*/:8'he7/* 231*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[8'hfc/* 252*/:8'hf2/* 242*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[9'h107/* 263*/:8'hfd/* 253*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[9'h112/* 274*/:9'h108/* 264*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[9'h11d/* 285*/:9'h113/* 275*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[9'h128/* 296*/:9'h11e/* 286*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[9'h133/* 307*/:9'h129/* 297*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[9'h13e/* 318*/:9'h134/* 308*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[9'h149/* 329*/:9'h13f/* 319*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[9'h154/* 340*/:9'h14a/* 330*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[9'h15f/* 351*/:9'h155/* 341*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[9'h16a/* 362*/:9'h160/* 352*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[9'h175/* 373*/:9'h16b/* 363*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[9'h180/* 384*/:9'h176/* 374*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[9'h18b/* 395*/:9'h181/* 385*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[9'h196/* 406*/:9'h18c/* 396*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[9'h1ac/* 428*/:9'h1a2/* 418*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[9'h1b7/* 439*/:9'h1ad/* 429*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[9'h1ba/* 442*/:9'h1b8/* 440*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[8'ha5/* 165*/:8'ha2/* 162*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[9'h1c5/* 453*/:9'h1bb/* 443*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[9'h1c8/* 456*/:9'h1c6/* 454*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[9'h1cb/* 459*/:9'h1c9/* 457*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[9'h1ce/* 462*/:9'h1cc/* 460*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[9'h1d1/* 465*/:9'h1cf/* 463*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[8'hb1/* 177*/:8'hae/* 174*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[9'h1dc/* 476*/:9'h1d2/* 466*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[9'h1df/* 479*/:9'h1dd/* 477*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[9'h1e2/* 482*/:9'h1e0/* 480*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[9'h1e5/* 485*/:9'h1e3/* 483*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[9'h1e8/* 488*/:9'h1e6/* 486*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[8'hbd/* 189*/:8'hba/* 186*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[9'h1f3/* 499*/:9'h1e9/* 489*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[9'h1f6/* 502*/:9'h1f4/* 500*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[8'hc1/* 193*/:8'hc0/* 192*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[9'h1f9/* 505*/:9'h1f7/* 503*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[8'hc3/* 195*/:8'hc2/* 194*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[9'h1fc/* 508*/:9'h1fa/* 506*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[9'h1ff/* 511*/:9'h1fd/* 509*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'hc9/* 201*/:8'hc6/* 198*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[10'h20a/* 522*/:10'h200/* 512*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[10'h20d/* 525*/:10'h20b/* 523*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[10'h210/* 528*/:10'h20e/* 526*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[10'h213/* 531*/:10'h211/* 529*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[10'h216/* 534*/:10'h214/* 532*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'hd5/* 213*/:8'hd2/* 210*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[10'h221/* 545*/:10'h217/* 535*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'hd7/* 215*/:8'hd6/* 214*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[10'h224/* 548*/:10'h222/* 546*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[10'h227/* 551*/:10'h225/* 549*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'hdb/* 219*/:8'hda/* 218*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[10'h22a/* 554*/:10'h228/* 552*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[10'h22d/* 557*/:10'h22b/* 555*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'he1/* 225*/:8'hde/* 222*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[10'h238/* 568*/:10'h22e/* 558*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'he3/* 227*/:8'he2/* 226*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[10'h23b/* 571*/:10'h239/* 569*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'he5/* 229*/:8'he4/* 228*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[10'h23e/* 574*/:10'h23c/* 572*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'he7/* 231*/:8'he6/* 230*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[10'h241/* 577*/:10'h23f/* 575*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'he9/* 233*/:8'he8/* 232*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[10'h244/* 580*/:10'h242/* 578*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'hed/* 237*/:8'hea/* 234*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[10'h24f/* 591*/:10'h245/* 581*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'hef/* 239*/:8'hee/* 238*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[10'h252/* 594*/:10'h250/* 592*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[10'h255/* 597*/:10'h253/* 595*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'hf3/* 243*/:8'hf2/* 242*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[10'h258/* 600*/:10'h256/* 598*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'hf5/* 245*/:8'hf4/* 244*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[10'h25b/* 603*/:10'h259/* 601*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'hf9/* 249*/:8'hf6/* 246*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[10'h266/* 614*/:10'h25c/* 604*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'hfb/* 251*/:8'hfa/* 250*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[10'h269/* 617*/:10'h267/* 615*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'hfd/* 253*/:8'hfc/* 252*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[10'h26c/* 620*/:10'h26a/* 618*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'hff/* 255*/:8'hfe/* 254*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[10'h26f/* 623*/:10'h26d/* 621*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[9'h101/* 257*/:9'h100/* 256*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[10'h272/* 626*/:10'h270/* 624*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[9'h105/* 261*/:9'h102/* 258*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[10'h27d/* 637*/:10'h273/* 627*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[9'h107/* 263*/:9'h106/* 262*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[10'h280/* 640*/:10'h27e/* 638*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[9'h109/* 265*/:9'h108/* 264*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[10'h283/* 643*/:10'h281/* 641*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[10'h286/* 646*/:10'h284/* 644*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[10'h289/* 649*/:10'h287/* 647*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[9'h111/* 273*/:9'h10e/* 270*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[10'h294/* 660*/:10'h28a/* 650*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[9'h113/* 275*/:9'h112/* 274*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[10'h297/* 663*/:10'h295/* 661*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[9'h115/* 277*/:9'h114/* 276*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[10'h29a/* 666*/:10'h298/* 664*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[9'h117/* 279*/:9'h116/* 278*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[10'h29d/* 669*/:10'h29b/* 667*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[9'h118/* 280*/:9'h118/* 280*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[10'h29f/* 671*/:10'h29e/* 670*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[9'h11c/* 284*/:9'h119/* 281*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[10'h2aa/* 682*/:10'h2a0/* 672*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[9'h11d/* 285*/:9'h11d/* 285*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[10'h2ac/* 684*/:10'h2ab/* 683*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[9'h11e/* 286*/:9'h11e/* 286*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[10'h2ae/* 686*/:10'h2ad/* 685*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[9'h11f/* 287*/:9'h11f/* 287*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[10'h2b0/* 688*/:10'h2af/* 687*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[9'h120/* 288*/:9'h120/* 288*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[10'h2b2/* 690*/:10'h2b1/* 689*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[9'h124/* 292*/:9'h121/* 289*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[10'h2bd/* 701*/:10'h2b3/* 691*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[9'h125/* 293*/:9'h125/* 293*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[10'h2bf/* 703*/:10'h2be/* 702*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[9'h126/* 294*/:9'h126/* 294*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[10'h2c1/* 705*/:10'h2c0/* 704*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[9'h127/* 295*/:9'h127/* 295*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[10'h2c3/* 707*/:10'h2c2/* 706*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[9'h128/* 296*/:9'h128/* 296*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[10'h2c5/* 709*/:10'h2c4/* 708*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[9'h12c/* 300*/:9'h129/* 297*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[10'h2d0/* 720*/:10'h2c6/* 710*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[9'h12d/* 301*/:9'h12d/* 301*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[10'h2d2/* 722*/:10'h2d1/* 721*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[9'h12e/* 302*/:9'h12e/* 302*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[10'h2d4/* 724*/:10'h2d3/* 723*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[9'h12f/* 303*/:9'h12f/* 303*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[10'h2d6/* 726*/:10'h2d5/* 725*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[9'h130/* 304*/:9'h130/* 304*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[10'h2d8/* 728*/:10'h2d7/* 727*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[9'h134/* 308*/:9'h131/* 305*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[10'h2e3/* 739*/:10'h2d9/* 729*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[9'h135/* 309*/:9'h135/* 309*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[10'h2e5/* 741*/:10'h2e4/* 740*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[9'h136/* 310*/:9'h136/* 310*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h2e7/* 743*/:10'h2e6/* 742*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[9'h137/* 311*/:9'h137/* 311*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h2e9/* 745*/:10'h2e8/* 744*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[9'h138/* 312*/:9'h138/* 312*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h2eb/* 747*/:10'h2ea/* 746*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[9'h13c/* 316*/:9'h139/* 313*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h2f6/* 758*/:10'h2ec/* 748*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[9'h13d/* 317*/:9'h13d/* 317*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h2f8/* 760*/:10'h2f7/* 759*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[9'h13e/* 318*/:9'h13e/* 318*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h2fa/* 762*/:10'h2f9/* 761*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h13f/* 319*/:9'h13f/* 319*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h2fc/* 764*/:10'h2fb/* 763*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h140/* 320*/:9'h140/* 320*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h2fe/* 766*/:10'h2fd/* 765*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h144/* 324*/:9'h141/* 321*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h309/* 777*/:10'h2ff/* 767*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h145/* 325*/:9'h145/* 325*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h30b/* 779*/:10'h30a/* 778*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h146/* 326*/:9'h146/* 326*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h30d/* 781*/:10'h30c/* 780*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h147/* 327*/:9'h147/* 327*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h30f/* 783*/:10'h30e/* 782*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h148/* 328*/:9'h148/* 328*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h311/* 785*/:10'h310/* 784*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h14c/* 332*/:9'h149/* 329*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h31c/* 796*/:10'h312/* 786*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h14d/* 333*/:9'h14d/* 333*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h31e/* 798*/:10'h31d/* 797*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h14e/* 334*/:9'h14e/* 334*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h320/* 800*/:10'h31f/* 799*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h14f/* 335*/:9'h14f/* 335*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h322/* 802*/:10'h321/* 801*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h150/* 336*/:9'h150/* 336*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h324/* 804*/:10'h323/* 803*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h154/* 340*/:9'h151/* 337*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h32f/* 815*/:10'h325/* 805*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h155/* 341*/:9'h155/* 341*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h331/* 817*/:10'h330/* 816*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h156/* 342*/:9'h156/* 342*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h333/* 819*/:10'h332/* 818*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h157/* 343*/:9'h157/* 343*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h335/* 821*/:10'h334/* 820*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h337/* 823*/:10'h336/* 822*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h15c/* 348*/:9'h159/* 345*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h342/* 834*/:10'h338/* 824*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h15d/* 349*/:9'h15d/* 349*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h344/* 836*/:10'h343/* 835*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h15e/* 350*/:9'h15e/* 350*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h346/* 838*/:10'h345/* 837*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h15f/* 351*/:9'h15f/* 351*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h348/* 840*/:10'h347/* 839*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h160/* 352*/:9'h160/* 352*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h34a/* 842*/:10'h349/* 841*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h164/* 356*/:9'h161/* 353*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h355/* 853*/:10'h34b/* 843*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h165/* 357*/:9'h165/* 357*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h357/* 855*/:10'h356/* 854*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h166/* 358*/:9'h166/* 358*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h359/* 857*/:10'h358/* 856*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h35a/* 858*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_11(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_9 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_10(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [859:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[10:0] T284;
  wire[10:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[10:0] T292;
  wire[10:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[10:0] T300;
  wire[10:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[10:0] T308;
  wire[10:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[10:0] T316;
  wire[10:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[10:0] T324;
  wire[10:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[10:0] T332;
  wire[10:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[10:0] T340;
  wire[10:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[10:0] T348;
  wire[10:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[10:0] T356;
  wire[10:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[10:0] T364;
  wire[10:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[10:0] T372;
  wire[10:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[10:0] T380;
  wire[10:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[10:0] T388;
  wire[10:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[10:0] T396;
  wire[10:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[10:0] T404;
  wire[10:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[10:0] T412;
  wire[10:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[10:0] T420;
  wire[10:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[10:0] T428;
  wire[10:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[3:0] T433;
  wire[3:0] T434;
  wire[3:0] T435;
  wire[10:0] T436;
  wire[10:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[3:0] T441;
  wire[3:0] T442;
  wire[3:0] T443;
  wire[10:0] T444;
  wire[10:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[3:0] T449;
  wire[3:0] T450;
  wire[3:0] T451;
  wire[10:0] T452;
  wire[10:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[10:0] T460;
  wire[10:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[10:0] T468;
  wire[10:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[3:0] T473;
  wire[3:0] T474;
  wire[3:0] T475;
  wire[10:0] T476;
  wire[10:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[3:0] T481;
  wire[3:0] T482;
  wire[3:0] T483;
  wire[10:0] T484;
  wire[10:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[10:0] T492;
  wire[10:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[10:0] T500;
  wire[10:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[10:0] T508;
  wire[10:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[10:0] T516;
  wire[10:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[3:0] T521;
  wire[3:0] T522;
  wire[3:0] T523;
  wire[10:0] T524;
  wire[10:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[10:0] T532;
  wire[10:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[10:0] T540;
  wire[10:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[10:0] T548;
  wire[10:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[3:0] T553;
  wire[3:0] T554;
  wire[3:0] T555;
  wire[10:0] T556;
  wire[10:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[3:0] T561;
  wire[3:0] T562;
  wire[3:0] T563;
  wire[10:0] T564;
  wire[10:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[3:0] T569;
  wire[3:0] T570;
  wire[3:0] T571;
  wire[10:0] T572;
  wire[10:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[10:0] T580;
  wire[10:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[10:0] T588;
  wire[10:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[3:0] T593;
  wire[3:0] T594;
  wire[3:0] T595;
  wire[10:0] T596;
  wire[10:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[3:0] T617;
  wire[3:0] T618;
  wire[3:0] T619;
  wire[10:0] T620;
  wire[10:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[3:0] T657;
  wire[3:0] T658;
  wire[3:0] T659;
  wire[10:0] T660;
  wire[10:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire[1:0] T681;
  wire[1:0] T682;
  wire[1:0] T683;
  wire[2:0] T684;
  wire[2:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire[1:0] T689;
  wire[1:0] T690;
  wire[1:0] T691;
  wire[2:0] T692;
  wire[2:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire[3:0] T697;
  wire[3:0] T698;
  wire[3:0] T699;
  wire[10:0] T700;
  wire[10:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire[1:0] T705;
  wire[1:0] T706;
  wire[1:0] T707;
  wire[2:0] T708;
  wire[2:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire[1:0] T713;
  wire[1:0] T714;
  wire[1:0] T715;
  wire[2:0] T716;
  wire[2:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire[1:0] T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[2:0] T724;
  wire[2:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire[1:0] T729;
  wire[1:0] T730;
  wire[1:0] T731;
  wire[2:0] T732;
  wire[2:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire[3:0] T737;
  wire[3:0] T738;
  wire[3:0] T739;
  wire[10:0] T740;
  wire[10:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire[1:0] T745;
  wire[1:0] T746;
  wire[1:0] T747;
  wire[2:0] T748;
  wire[2:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire[1:0] T753;
  wire[1:0] T754;
  wire[1:0] T755;
  wire[2:0] T756;
  wire[2:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[3:0] T777;
  wire[3:0] T778;
  wire[3:0] T779;
  wire[10:0] T780;
  wire[10:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[1:0] T793;
  wire[1:0] T794;
  wire[1:0] T795;
  wire[2:0] T796;
  wire[2:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire[1:0] T801;
  wire[1:0] T802;
  wire[1:0] T803;
  wire[2:0] T804;
  wire[2:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[1:0] T809;
  wire[1:0] T810;
  wire[1:0] T811;
  wire[2:0] T812;
  wire[2:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[3:0] T817;
  wire[3:0] T818;
  wire[3:0] T819;
  wire[10:0] T820;
  wire[10:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[1:0] T825;
  wire[1:0] T826;
  wire[1:0] T827;
  wire[2:0] T828;
  wire[2:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[1:0] T833;
  wire[1:0] T834;
  wire[1:0] T835;
  wire[2:0] T836;
  wire[2:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire[1:0] T841;
  wire[1:0] T842;
  wire[1:0] T843;
  wire[2:0] T844;
  wire[2:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire[1:0] T849;
  wire[1:0] T850;
  wire[1:0] T851;
  wire[2:0] T852;
  wire[2:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire[3:0] T857;
  wire[3:0] T858;
  wire[3:0] T859;
  wire[10:0] T860;
  wire[10:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire[1:0] T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[2:0] T868;
  wire[2:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire[1:0] T873;
  wire[1:0] T874;
  wire[1:0] T875;
  wire[2:0] T876;
  wire[2:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire[1:0] T881;
  wire[1:0] T882;
  wire[1:0] T883;
  wire[2:0] T884;
  wire[2:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire[1:0] T889;
  wire[1:0] T890;
  wire[1:0] T891;
  wire[2:0] T892;
  wire[2:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire[3:0] T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[10:0] T900;
  wire[10:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire[1:0] T905;
  wire[1:0] T906;
  wire[1:0] T907;
  wire[2:0] T908;
  wire[2:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire[1:0] T913;
  wire[1:0] T914;
  wire[1:0] T915;
  wire[2:0] T916;
  wire[2:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire[1:0] T922;
  wire[1:0] T923;
  wire[2:0] T924;
  wire[2:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[2:0] T932;
  wire[2:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[3:0] T937;
  wire[3:0] T938;
  wire[3:0] T939;
  wire[10:0] T940;
  wire[10:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[1:0] T945;
  wire[1:0] T946;
  wire[1:0] T947;
  wire[2:0] T948;
  wire[2:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[1:0] T953;
  wire[1:0] T954;
  wire[1:0] T955;
  wire[2:0] T956;
  wire[2:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[1:0] T961;
  wire[1:0] T962;
  wire[1:0] T963;
  wire[2:0] T964;
  wire[2:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[1:0] T969;
  wire[1:0] T970;
  wire[1:0] T971;
  wire[2:0] T972;
  wire[2:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[3:0] T977;
  wire[3:0] T978;
  wire[3:0] T979;
  wire[10:0] T980;
  wire[10:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[1:0] T985;
  wire[1:0] T986;
  wire[1:0] T987;
  wire[2:0] T988;
  wire[2:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[1:0] T993;
  wire[1:0] T994;
  wire[1:0] T995;
  wire[2:0] T996;
  wire[2:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire[3:0] T1017;
  wire[3:0] T1018;
  wire[3:0] T1019;
  wire[10:0] T1020;
  wire[10:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire[3:0] T1057;
  wire[3:0] T1058;
  wire[3:0] T1059;
  wire[10:0] T1060;
  wire[10:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire[1:0] T1084;
  wire[1:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire[1:0] T1092;
  wire[1:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[10:0] T1100;
  wire[10:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[1:0] T1108;
  wire[1:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire T1113;
  wire T1114;
  wire T1115;
  wire[1:0] T1116;
  wire[1:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[1:0] T1124;
  wire[1:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[1:0] T1132;
  wire[1:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[3:0] T1137;
  wire[3:0] T1138;
  wire[3:0] T1139;
  wire[10:0] T1140;
  wire[10:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire T1145;
  wire T1146;
  wire T1147;
  wire[1:0] T1148;
  wire[1:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire T1153;
  wire T1154;
  wire T1155;
  wire[1:0] T1156;
  wire[1:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire[1:0] T1164;
  wire[1:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire T1170;
  wire T1171;
  wire[1:0] T1172;
  wire[1:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[10:0] T1180;
  wire[10:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire T1185;
  wire T1186;
  wire T1187;
  wire[1:0] T1188;
  wire[1:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire[1:0] T1196;
  wire[1:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire[1:0] T1204;
  wire[1:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire T1209;
  wire T1210;
  wire T1211;
  wire[1:0] T1212;
  wire[1:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[3:0] T1217;
  wire[3:0] T1218;
  wire[3:0] T1219;
  wire[10:0] T1220;
  wire[10:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire[1:0] T1228;
  wire[1:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire[1:0] T1236;
  wire[1:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire[1:0] T1244;
  wire[1:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[1:0] T1252;
  wire[1:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[10:0] T1260;
  wire[10:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[1:0] T1268;
  wire[1:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[1:0] T1276;
  wire[1:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire T1289;
  wire T1290;
  wire T1291;
  wire[1:0] T1292;
  wire[1:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire[3:0] T1297;
  wire[3:0] T1298;
  wire[3:0] T1299;
  wire[10:0] T1300;
  wire[10:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire[1:0] T1308;
  wire[1:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire[1:0] T1324;
  wire[1:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[10:0] T1340;
  wire[10:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire T1353;
  wire T1354;
  wire T1355;
  wire[1:0] T1356;
  wire[1:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire[1:0] T1364;
  wire[1:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire[1:0] T1372;
  wire[1:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire[3:0] T1377;
  wire[3:0] T1378;
  wire[3:0] T1379;
  wire[10:0] T1380;
  wire[10:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire[1:0] T1388;
  wire[1:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[1:0] T1396;
  wire[1:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[4'ha/* 10*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h15/* 21*/:4'hb/* 11*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[6'h20/* 32*/:5'h16/* 22*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h2b/* 43*/:6'h21/* 33*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h36/* 54*/:6'h2c/* 44*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[7'h41/* 65*/:6'h37/* 55*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[7'h4c/* 76*/:7'h42/* 66*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[7'h57/* 87*/:7'h4d/* 77*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h62/* 98*/:7'h58/* 88*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h6d/* 109*/:7'h63/* 99*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h78/* 120*/:7'h6e/* 110*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[8'h83/* 131*/:7'h79/* 121*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[8'h8e/* 142*/:8'h84/* 132*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[8'h99/* 153*/:8'h8f/* 143*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[8'ha4/* 164*/:8'h9a/* 154*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[8'haf/* 175*/:8'ha5/* 165*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[8'hba/* 186*/:8'hb0/* 176*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[8'hc5/* 197*/:8'hbb/* 187*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[8'hd0/* 208*/:8'hc6/* 198*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[8'hdb/* 219*/:8'hd1/* 209*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[8'he6/* 230*/:8'hdc/* 220*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[8'hf1/* 241*/:8'he7/* 231*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[8'hfc/* 252*/:8'hf2/* 242*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[9'h107/* 263*/:8'hfd/* 253*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[9'h112/* 274*/:9'h108/* 264*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[9'h11d/* 285*/:9'h113/* 275*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[9'h128/* 296*/:9'h11e/* 286*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[9'h133/* 307*/:9'h129/* 297*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[9'h13e/* 318*/:9'h134/* 308*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[9'h149/* 329*/:9'h13f/* 319*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[9'h154/* 340*/:9'h14a/* 330*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[9'h15f/* 351*/:9'h155/* 341*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[9'h16a/* 362*/:9'h160/* 352*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[9'h175/* 373*/:9'h16b/* 363*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[9'h180/* 384*/:9'h176/* 374*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[9'h18b/* 395*/:9'h181/* 385*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[9'h196/* 406*/:9'h18c/* 396*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[9'h1a1/* 417*/:9'h197/* 407*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[9'h1ac/* 428*/:9'h1a2/* 418*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[9'h1b7/* 439*/:9'h1ad/* 429*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[9'h1ba/* 442*/:9'h1b8/* 440*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[9'h1bd/* 445*/:9'h1bb/* 443*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[8'ha7/* 167*/:8'ha4/* 164*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[9'h1c8/* 456*/:9'h1be/* 446*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[9'h1cb/* 459*/:9'h1c9/* 457*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[9'h1ce/* 462*/:9'h1cc/* 460*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[9'h1d1/* 465*/:9'h1cf/* 463*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[9'h1d4/* 468*/:9'h1d2/* 466*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[8'hb3/* 179*/:8'hb0/* 176*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[9'h1df/* 479*/:9'h1d5/* 469*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[8'hb5/* 181*/:8'hb4/* 180*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[9'h1e2/* 482*/:9'h1e0/* 480*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[8'hb7/* 183*/:8'hb6/* 182*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[9'h1e5/* 485*/:9'h1e3/* 483*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[8'hb9/* 185*/:8'hb8/* 184*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[9'h1e8/* 488*/:9'h1e6/* 486*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[8'hbb/* 187*/:8'hba/* 186*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[9'h1eb/* 491*/:9'h1e9/* 489*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[8'hbf/* 191*/:8'hbc/* 188*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[9'h1f6/* 502*/:9'h1ec/* 492*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[8'hc1/* 193*/:8'hc0/* 192*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[9'h1f9/* 505*/:9'h1f7/* 503*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[8'hc3/* 195*/:8'hc2/* 194*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[9'h1fc/* 508*/:9'h1fa/* 506*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[9'h1ff/* 511*/:9'h1fd/* 509*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[10'h202/* 514*/:10'h200/* 512*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'hcb/* 203*/:8'hc8/* 200*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[10'h20d/* 525*/:10'h203/* 515*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[10'h210/* 528*/:10'h20e/* 526*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[10'h213/* 531*/:10'h211/* 529*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[10'h216/* 534*/:10'h214/* 532*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'hd3/* 211*/:8'hd2/* 210*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[10'h219/* 537*/:10'h217/* 535*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'hd7/* 215*/:8'hd4/* 212*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[10'h224/* 548*/:10'h21a/* 538*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'hd9/* 217*/:8'hd8/* 216*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[10'h227/* 551*/:10'h225/* 549*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'hdb/* 219*/:8'hda/* 218*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[10'h22a/* 554*/:10'h228/* 552*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[10'h22d/* 557*/:10'h22b/* 555*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[10'h230/* 560*/:10'h22e/* 558*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'he3/* 227*/:8'he0/* 224*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[10'h23b/* 571*/:10'h231/* 561*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'he5/* 229*/:8'he4/* 228*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[10'h23e/* 574*/:10'h23c/* 572*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'he7/* 231*/:8'he6/* 230*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[10'h241/* 577*/:10'h23f/* 575*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'he9/* 233*/:8'he8/* 232*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[10'h244/* 580*/:10'h242/* 578*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'heb/* 235*/:8'hea/* 234*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[10'h247/* 583*/:10'h245/* 581*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'hef/* 239*/:8'hec/* 236*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[10'h252/* 594*/:10'h248/* 584*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'hf1/* 241*/:8'hf0/* 240*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[10'h255/* 597*/:10'h253/* 595*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'hf3/* 243*/:8'hf2/* 242*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[10'h258/* 600*/:10'h256/* 598*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'hf5/* 245*/:8'hf4/* 244*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[10'h25b/* 603*/:10'h259/* 601*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'hf7/* 247*/:8'hf6/* 246*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[10'h25e/* 606*/:10'h25c/* 604*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'hfb/* 251*/:8'hf8/* 248*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[10'h269/* 617*/:10'h25f/* 607*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'hfd/* 253*/:8'hfc/* 252*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[10'h26c/* 620*/:10'h26a/* 618*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'hff/* 255*/:8'hfe/* 254*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[10'h26f/* 623*/:10'h26d/* 621*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[9'h101/* 257*/:9'h100/* 256*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[10'h272/* 626*/:10'h270/* 624*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[9'h103/* 259*/:9'h102/* 258*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[10'h275/* 629*/:10'h273/* 627*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[9'h107/* 263*/:9'h104/* 260*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[10'h280/* 640*/:10'h276/* 630*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[9'h109/* 265*/:9'h108/* 264*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[10'h283/* 643*/:10'h281/* 641*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[10'h286/* 646*/:10'h284/* 644*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[9'h10d/* 269*/:9'h10c/* 268*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[10'h289/* 649*/:10'h287/* 647*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[9'h10f/* 271*/:9'h10e/* 270*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[10'h28c/* 652*/:10'h28a/* 650*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[9'h113/* 275*/:9'h110/* 272*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[10'h297/* 663*/:10'h28d/* 653*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[9'h115/* 277*/:9'h114/* 276*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[10'h29a/* 666*/:10'h298/* 664*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[9'h117/* 279*/:9'h116/* 278*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[10'h29d/* 669*/:10'h29b/* 667*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[9'h118/* 280*/:9'h118/* 280*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[10'h29f/* 671*/:10'h29e/* 670*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[9'h119/* 281*/:9'h119/* 281*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[10'h2a1/* 673*/:10'h2a0/* 672*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[9'h11d/* 285*/:9'h11a/* 282*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[10'h2ac/* 684*/:10'h2a2/* 674*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[9'h11e/* 286*/:9'h11e/* 286*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[10'h2ae/* 686*/:10'h2ad/* 685*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[9'h11f/* 287*/:9'h11f/* 287*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[10'h2b0/* 688*/:10'h2af/* 687*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[9'h120/* 288*/:9'h120/* 288*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[10'h2b2/* 690*/:10'h2b1/* 689*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[9'h121/* 289*/:9'h121/* 289*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[10'h2b4/* 692*/:10'h2b3/* 691*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[9'h125/* 293*/:9'h122/* 290*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[10'h2bf/* 703*/:10'h2b5/* 693*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[9'h126/* 294*/:9'h126/* 294*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[10'h2c1/* 705*/:10'h2c0/* 704*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[9'h127/* 295*/:9'h127/* 295*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[10'h2c3/* 707*/:10'h2c2/* 706*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[9'h128/* 296*/:9'h128/* 296*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[10'h2c5/* 709*/:10'h2c4/* 708*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[9'h129/* 297*/:9'h129/* 297*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[10'h2c7/* 711*/:10'h2c6/* 710*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[9'h12d/* 301*/:9'h12a/* 298*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[10'h2d2/* 722*/:10'h2c8/* 712*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[9'h12e/* 302*/:9'h12e/* 302*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[10'h2d4/* 724*/:10'h2d3/* 723*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[9'h12f/* 303*/:9'h12f/* 303*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[10'h2d6/* 726*/:10'h2d5/* 725*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[9'h130/* 304*/:9'h130/* 304*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[10'h2d8/* 728*/:10'h2d7/* 727*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[9'h131/* 305*/:9'h131/* 305*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[10'h2da/* 730*/:10'h2d9/* 729*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[9'h135/* 309*/:9'h132/* 306*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[10'h2e5/* 741*/:10'h2db/* 731*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[9'h136/* 310*/:9'h136/* 310*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h2e7/* 743*/:10'h2e6/* 742*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[9'h137/* 311*/:9'h137/* 311*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h2e9/* 745*/:10'h2e8/* 744*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[9'h138/* 312*/:9'h138/* 312*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h2eb/* 747*/:10'h2ea/* 746*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[9'h139/* 313*/:9'h139/* 313*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h2ed/* 749*/:10'h2ec/* 748*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[9'h13d/* 317*/:9'h13a/* 314*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h2f8/* 760*/:10'h2ee/* 750*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[9'h13e/* 318*/:9'h13e/* 318*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h2fa/* 762*/:10'h2f9/* 761*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h13f/* 319*/:9'h13f/* 319*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h2fc/* 764*/:10'h2fb/* 763*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h140/* 320*/:9'h140/* 320*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h2fe/* 766*/:10'h2fd/* 765*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h141/* 321*/:9'h141/* 321*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h300/* 768*/:10'h2ff/* 767*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h145/* 325*/:9'h142/* 322*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h30b/* 779*/:10'h301/* 769*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h146/* 326*/:9'h146/* 326*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h30d/* 781*/:10'h30c/* 780*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h147/* 327*/:9'h147/* 327*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h30f/* 783*/:10'h30e/* 782*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h148/* 328*/:9'h148/* 328*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h311/* 785*/:10'h310/* 784*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h313/* 787*/:10'h312/* 786*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h14d/* 333*/:9'h14a/* 330*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h31e/* 798*/:10'h314/* 788*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h14e/* 334*/:9'h14e/* 334*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h320/* 800*/:10'h31f/* 799*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h14f/* 335*/:9'h14f/* 335*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h322/* 802*/:10'h321/* 801*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h150/* 336*/:9'h150/* 336*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h324/* 804*/:10'h323/* 803*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h151/* 337*/:9'h151/* 337*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h326/* 806*/:10'h325/* 805*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h155/* 341*/:9'h152/* 338*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h331/* 817*/:10'h327/* 807*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h156/* 342*/:9'h156/* 342*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h333/* 819*/:10'h332/* 818*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h157/* 343*/:9'h157/* 343*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h335/* 821*/:10'h334/* 820*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h337/* 823*/:10'h336/* 822*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h159/* 345*/:9'h159/* 345*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h339/* 825*/:10'h338/* 824*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h15d/* 349*/:9'h15a/* 346*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h344/* 836*/:10'h33a/* 826*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h15e/* 350*/:9'h15e/* 350*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h346/* 838*/:10'h345/* 837*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h15f/* 351*/:9'h15f/* 351*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h348/* 840*/:10'h347/* 839*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h160/* 352*/:9'h160/* 352*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h34a/* 842*/:10'h349/* 841*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h161/* 353*/:9'h161/* 353*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h34c/* 844*/:10'h34b/* 843*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h165/* 357*/:9'h162/* 354*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h357/* 855*/:10'h34d/* 845*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h166/* 358*/:9'h166/* 358*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h359/* 857*/:10'h358/* 856*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h35b/* 859*/:10'h35a/* 858*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_12(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [859:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {7'h0/* 0*/, 1'h1/* 1*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_10 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module sbcb_sp_11(
    input [527:0] io_ipin_in,
    input [131:0] io_ipin_config,
    input [779:0] io_chanxy_in,
    input [359:0] io_chanxy_config,
    output[32:0] io_ipin_out,
    output[139:0] io_chanxy_out);

  wire[139:0] T0;
  wire[139:0] T1;
  wire[138:0] T2;
  wire[138:0] T3;
  wire[137:0] T4;
  wire[137:0] T5;
  wire[136:0] T6;
  wire[136:0] T7;
  wire[135:0] T8;
  wire[135:0] T9;
  wire[134:0] T10;
  wire[134:0] T11;
  wire[133:0] T12;
  wire[133:0] T13;
  wire[132:0] T14;
  wire[132:0] T15;
  wire[131:0] T16;
  wire[131:0] T17;
  wire[130:0] T18;
  wire[130:0] T19;
  wire[129:0] T20;
  wire[129:0] T21;
  wire[128:0] T22;
  wire[128:0] T23;
  wire[127:0] T24;
  wire[127:0] T25;
  wire[126:0] T26;
  wire[126:0] T27;
  wire[125:0] T28;
  wire[125:0] T29;
  wire[124:0] T30;
  wire[124:0] T31;
  wire[123:0] T32;
  wire[123:0] T33;
  wire[122:0] T34;
  wire[122:0] T35;
  wire[121:0] T36;
  wire[121:0] T37;
  wire[120:0] T38;
  wire[120:0] T39;
  wire[119:0] T40;
  wire[119:0] T41;
  wire[118:0] T42;
  wire[118:0] T43;
  wire[117:0] T44;
  wire[117:0] T45;
  wire[116:0] T46;
  wire[116:0] T47;
  wire[115:0] T48;
  wire[115:0] T49;
  wire[114:0] T50;
  wire[114:0] T51;
  wire[113:0] T52;
  wire[113:0] T53;
  wire[112:0] T54;
  wire[112:0] T55;
  wire[111:0] T56;
  wire[111:0] T57;
  wire[110:0] T58;
  wire[110:0] T59;
  wire[109:0] T60;
  wire[109:0] T61;
  wire[108:0] T62;
  wire[108:0] T63;
  wire[107:0] T64;
  wire[107:0] T65;
  wire[106:0] T66;
  wire[106:0] T67;
  wire[105:0] T68;
  wire[105:0] T69;
  wire[104:0] T70;
  wire[104:0] T71;
  wire[103:0] T72;
  wire[103:0] T73;
  wire[102:0] T74;
  wire[102:0] T75;
  wire[101:0] T76;
  wire[101:0] T77;
  wire[100:0] T78;
  wire[100:0] T79;
  wire[99:0] T80;
  wire[99:0] T81;
  wire[98:0] T82;
  wire[98:0] T83;
  wire[97:0] T84;
  wire[97:0] T85;
  wire[96:0] T86;
  wire[96:0] T87;
  wire[95:0] T88;
  wire[95:0] T89;
  wire[94:0] T90;
  wire[94:0] T91;
  wire[93:0] T92;
  wire[93:0] T93;
  wire[92:0] T94;
  wire[92:0] T95;
  wire[91:0] T96;
  wire[91:0] T97;
  wire[90:0] T98;
  wire[90:0] T99;
  wire[89:0] T100;
  wire[89:0] T101;
  wire[88:0] T102;
  wire[88:0] T103;
  wire[87:0] T104;
  wire[87:0] T105;
  wire[86:0] T106;
  wire[86:0] T107;
  wire[85:0] T108;
  wire[85:0] T109;
  wire[84:0] T110;
  wire[84:0] T111;
  wire[83:0] T112;
  wire[83:0] T113;
  wire[82:0] T114;
  wire[82:0] T115;
  wire[81:0] T116;
  wire[81:0] T117;
  wire[80:0] T118;
  wire[80:0] T119;
  wire[79:0] T120;
  wire[79:0] T121;
  wire[78:0] T122;
  wire[78:0] T123;
  wire[77:0] T124;
  wire[77:0] T125;
  wire[76:0] T126;
  wire[76:0] T127;
  wire[75:0] T128;
  wire[75:0] T129;
  wire[74:0] T130;
  wire[74:0] T131;
  wire[73:0] T132;
  wire[73:0] T133;
  wire[72:0] T134;
  wire[72:0] T135;
  wire[71:0] T136;
  wire[71:0] T137;
  wire[70:0] T138;
  wire[70:0] T139;
  wire[69:0] T140;
  wire[69:0] T141;
  wire[68:0] T142;
  wire[68:0] T143;
  wire[67:0] T144;
  wire[67:0] T145;
  wire[66:0] T146;
  wire[66:0] T147;
  wire[65:0] T148;
  wire[65:0] T149;
  wire[64:0] T150;
  wire[64:0] T151;
  wire[63:0] T152;
  wire[63:0] T153;
  wire[62:0] T154;
  wire[62:0] T155;
  wire[61:0] T156;
  wire[61:0] T157;
  wire[60:0] T158;
  wire[60:0] T159;
  wire[59:0] T160;
  wire[59:0] T161;
  wire[58:0] T162;
  wire[58:0] T163;
  wire[57:0] T164;
  wire[57:0] T165;
  wire[56:0] T166;
  wire[56:0] T167;
  wire[55:0] T168;
  wire[55:0] T169;
  wire[54:0] T170;
  wire[54:0] T171;
  wire[53:0] T172;
  wire[53:0] T173;
  wire[52:0] T174;
  wire[52:0] T175;
  wire[51:0] T176;
  wire[51:0] T177;
  wire[50:0] T178;
  wire[50:0] T179;
  wire[49:0] T180;
  wire[49:0] T181;
  wire[48:0] T182;
  wire[48:0] T183;
  wire[47:0] T184;
  wire[47:0] T185;
  wire[46:0] T186;
  wire[46:0] T187;
  wire[45:0] T188;
  wire[45:0] T189;
  wire[44:0] T190;
  wire[44:0] T191;
  wire[43:0] T192;
  wire[43:0] T193;
  wire[42:0] T194;
  wire[42:0] T195;
  wire[41:0] T196;
  wire[41:0] T197;
  wire[40:0] T198;
  wire[40:0] T199;
  wire[39:0] T200;
  wire[39:0] T201;
  wire[38:0] T202;
  wire[38:0] T203;
  wire[37:0] T204;
  wire[37:0] T205;
  wire[36:0] T206;
  wire[36:0] T207;
  wire[35:0] T208;
  wire[35:0] T209;
  wire[34:0] T210;
  wire[34:0] T211;
  wire[33:0] T212;
  wire[33:0] T213;
  wire[32:0] T214;
  wire[32:0] T215;
  wire[31:0] T216;
  wire[31:0] T217;
  wire[30:0] T218;
  wire[30:0] T219;
  wire[29:0] T220;
  wire[29:0] T221;
  wire[28:0] T222;
  wire[28:0] T223;
  wire[27:0] T224;
  wire[27:0] T225;
  wire[26:0] T226;
  wire[26:0] T227;
  wire[25:0] T228;
  wire[25:0] T229;
  wire[24:0] T230;
  wire[24:0] T231;
  wire[23:0] T232;
  wire[23:0] T233;
  wire[22:0] T234;
  wire[22:0] T235;
  wire[21:0] T236;
  wire[21:0] T237;
  wire[20:0] T238;
  wire[20:0] T239;
  wire[19:0] T240;
  wire[19:0] T241;
  wire[18:0] T242;
  wire[18:0] T243;
  wire[17:0] T244;
  wire[17:0] T245;
  wire[16:0] T246;
  wire[16:0] T247;
  wire[15:0] T248;
  wire[15:0] T249;
  wire[14:0] T250;
  wire[14:0] T251;
  wire[13:0] T252;
  wire[13:0] T253;
  wire[12:0] T254;
  wire[12:0] T255;
  wire[11:0] T256;
  wire[11:0] T257;
  wire[10:0] T258;
  wire[10:0] T259;
  wire[9:0] T260;
  wire[9:0] T261;
  wire[8:0] T262;
  wire[8:0] T263;
  wire[7:0] T264;
  wire[7:0] T265;
  wire[6:0] T266;
  wire[6:0] T267;
  wire[5:0] T268;
  wire[5:0] T269;
  wire[4:0] T270;
  wire[4:0] T271;
  wire[3:0] T272;
  wire[3:0] T273;
  wire[2:0] T274;
  wire[2:0] T275;
  wire[1:0] T276;
  wire[1:0] T277;
  wire T278;
  wire T279;
  wire T280;
  wire[3:0] T281;
  wire[3:0] T282;
  wire[3:0] T283;
  wire[8:0] T284;
  wire[8:0] T285;
  wire T286;
  wire T287;
  wire T288;
  wire[3:0] T289;
  wire[3:0] T290;
  wire[3:0] T291;
  wire[8:0] T292;
  wire[8:0] T293;
  wire T294;
  wire T295;
  wire T296;
  wire[3:0] T297;
  wire[3:0] T298;
  wire[3:0] T299;
  wire[8:0] T300;
  wire[8:0] T301;
  wire T302;
  wire T303;
  wire T304;
  wire[3:0] T305;
  wire[3:0] T306;
  wire[3:0] T307;
  wire[8:0] T308;
  wire[8:0] T309;
  wire T310;
  wire T311;
  wire T312;
  wire[3:0] T313;
  wire[3:0] T314;
  wire[3:0] T315;
  wire[8:0] T316;
  wire[8:0] T317;
  wire T318;
  wire T319;
  wire T320;
  wire[3:0] T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[8:0] T324;
  wire[8:0] T325;
  wire T326;
  wire T327;
  wire T328;
  wire[3:0] T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire[8:0] T332;
  wire[8:0] T333;
  wire T334;
  wire T335;
  wire T336;
  wire[3:0] T337;
  wire[3:0] T338;
  wire[3:0] T339;
  wire[8:0] T340;
  wire[8:0] T341;
  wire T342;
  wire T343;
  wire T344;
  wire[3:0] T345;
  wire[3:0] T346;
  wire[3:0] T347;
  wire[8:0] T348;
  wire[8:0] T349;
  wire T350;
  wire T351;
  wire T352;
  wire[3:0] T353;
  wire[3:0] T354;
  wire[3:0] T355;
  wire[8:0] T356;
  wire[8:0] T357;
  wire T358;
  wire T359;
  wire T360;
  wire[3:0] T361;
  wire[3:0] T362;
  wire[3:0] T363;
  wire[8:0] T364;
  wire[8:0] T365;
  wire T366;
  wire T367;
  wire T368;
  wire[3:0] T369;
  wire[3:0] T370;
  wire[3:0] T371;
  wire[8:0] T372;
  wire[8:0] T373;
  wire T374;
  wire T375;
  wire T376;
  wire[3:0] T377;
  wire[3:0] T378;
  wire[3:0] T379;
  wire[8:0] T380;
  wire[8:0] T381;
  wire T382;
  wire T383;
  wire T384;
  wire[3:0] T385;
  wire[3:0] T386;
  wire[3:0] T387;
  wire[8:0] T388;
  wire[8:0] T389;
  wire T390;
  wire T391;
  wire T392;
  wire[3:0] T393;
  wire[3:0] T394;
  wire[3:0] T395;
  wire[8:0] T396;
  wire[8:0] T397;
  wire T398;
  wire T399;
  wire T400;
  wire[3:0] T401;
  wire[3:0] T402;
  wire[3:0] T403;
  wire[8:0] T404;
  wire[8:0] T405;
  wire T406;
  wire T407;
  wire T408;
  wire[3:0] T409;
  wire[3:0] T410;
  wire[3:0] T411;
  wire[8:0] T412;
  wire[8:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire[3:0] T417;
  wire[3:0] T418;
  wire[3:0] T419;
  wire[8:0] T420;
  wire[8:0] T421;
  wire T422;
  wire T423;
  wire T424;
  wire[3:0] T425;
  wire[3:0] T426;
  wire[3:0] T427;
  wire[8:0] T428;
  wire[8:0] T429;
  wire T430;
  wire T431;
  wire T432;
  wire[3:0] T433;
  wire[3:0] T434;
  wire[3:0] T435;
  wire[8:0] T436;
  wire[8:0] T437;
  wire T438;
  wire T439;
  wire T440;
  wire[3:0] T441;
  wire[3:0] T442;
  wire[3:0] T443;
  wire[8:0] T444;
  wire[8:0] T445;
  wire T446;
  wire T447;
  wire T448;
  wire[3:0] T449;
  wire[3:0] T450;
  wire[3:0] T451;
  wire[8:0] T452;
  wire[8:0] T453;
  wire T454;
  wire T455;
  wire T456;
  wire[3:0] T457;
  wire[3:0] T458;
  wire[3:0] T459;
  wire[8:0] T460;
  wire[8:0] T461;
  wire T462;
  wire T463;
  wire T464;
  wire[3:0] T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[8:0] T468;
  wire[8:0] T469;
  wire T470;
  wire T471;
  wire T472;
  wire[3:0] T473;
  wire[3:0] T474;
  wire[3:0] T475;
  wire[8:0] T476;
  wire[8:0] T477;
  wire T478;
  wire T479;
  wire T480;
  wire[3:0] T481;
  wire[3:0] T482;
  wire[3:0] T483;
  wire[8:0] T484;
  wire[8:0] T485;
  wire T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[3:0] T490;
  wire[3:0] T491;
  wire[8:0] T492;
  wire[8:0] T493;
  wire T494;
  wire T495;
  wire T496;
  wire[3:0] T497;
  wire[3:0] T498;
  wire[3:0] T499;
  wire[8:0] T500;
  wire[8:0] T501;
  wire T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[3:0] T506;
  wire[3:0] T507;
  wire[8:0] T508;
  wire[8:0] T509;
  wire T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire[3:0] T514;
  wire[3:0] T515;
  wire[8:0] T516;
  wire[8:0] T517;
  wire T518;
  wire T519;
  wire T520;
  wire[3:0] T521;
  wire[3:0] T522;
  wire[3:0] T523;
  wire[8:0] T524;
  wire[8:0] T525;
  wire T526;
  wire T527;
  wire T528;
  wire[3:0] T529;
  wire[3:0] T530;
  wire[3:0] T531;
  wire[8:0] T532;
  wire[8:0] T533;
  wire T534;
  wire T535;
  wire T536;
  wire[3:0] T537;
  wire[3:0] T538;
  wire[3:0] T539;
  wire[8:0] T540;
  wire[8:0] T541;
  wire T542;
  wire T543;
  wire T544;
  wire[3:0] T545;
  wire[3:0] T546;
  wire[3:0] T547;
  wire[8:0] T548;
  wire[8:0] T549;
  wire T550;
  wire T551;
  wire T552;
  wire[3:0] T553;
  wire[3:0] T554;
  wire[3:0] T555;
  wire[8:0] T556;
  wire[8:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire[3:0] T561;
  wire[3:0] T562;
  wire[3:0] T563;
  wire[8:0] T564;
  wire[8:0] T565;
  wire T566;
  wire T567;
  wire T568;
  wire[3:0] T569;
  wire[3:0] T570;
  wire[3:0] T571;
  wire[8:0] T572;
  wire[8:0] T573;
  wire T574;
  wire T575;
  wire T576;
  wire[3:0] T577;
  wire[3:0] T578;
  wire[3:0] T579;
  wire[8:0] T580;
  wire[8:0] T581;
  wire T582;
  wire T583;
  wire T584;
  wire[3:0] T585;
  wire[3:0] T586;
  wire[3:0] T587;
  wire[8:0] T588;
  wire[8:0] T589;
  wire T590;
  wire T591;
  wire T592;
  wire[3:0] T593;
  wire[3:0] T594;
  wire[3:0] T595;
  wire[8:0] T596;
  wire[8:0] T597;
  wire T598;
  wire T599;
  wire T600;
  wire[1:0] T601;
  wire[1:0] T602;
  wire[1:0] T603;
  wire[2:0] T604;
  wire[2:0] T605;
  wire T606;
  wire T607;
  wire T608;
  wire[1:0] T609;
  wire[1:0] T610;
  wire[1:0] T611;
  wire[2:0] T612;
  wire[2:0] T613;
  wire T614;
  wire T615;
  wire T616;
  wire[1:0] T617;
  wire[1:0] T618;
  wire[1:0] T619;
  wire[2:0] T620;
  wire[2:0] T621;
  wire T622;
  wire T623;
  wire T624;
  wire[1:0] T625;
  wire[1:0] T626;
  wire[1:0] T627;
  wire[2:0] T628;
  wire[2:0] T629;
  wire T630;
  wire T631;
  wire T632;
  wire[1:0] T633;
  wire[1:0] T634;
  wire[1:0] T635;
  wire[2:0] T636;
  wire[2:0] T637;
  wire T638;
  wire T639;
  wire T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[2:0] T644;
  wire[2:0] T645;
  wire T646;
  wire T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[1:0] T651;
  wire[2:0] T652;
  wire[2:0] T653;
  wire T654;
  wire T655;
  wire T656;
  wire[1:0] T657;
  wire[1:0] T658;
  wire[1:0] T659;
  wire[2:0] T660;
  wire[2:0] T661;
  wire T662;
  wire T663;
  wire T664;
  wire[1:0] T665;
  wire[1:0] T666;
  wire[1:0] T667;
  wire[2:0] T668;
  wire[2:0] T669;
  wire T670;
  wire T671;
  wire T672;
  wire[1:0] T673;
  wire[1:0] T674;
  wire[1:0] T675;
  wire[2:0] T676;
  wire[2:0] T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire[1:0] T684;
  wire[1:0] T685;
  wire T686;
  wire T687;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[1:0] T692;
  wire[1:0] T693;
  wire T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[1:0] T700;
  wire[1:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire[1:0] T708;
  wire[1:0] T709;
  wire T710;
  wire T711;
  wire T712;
  wire T713;
  wire T714;
  wire T715;
  wire[1:0] T716;
  wire[1:0] T717;
  wire T718;
  wire T719;
  wire T720;
  wire T721;
  wire T722;
  wire T723;
  wire[1:0] T724;
  wire[1:0] T725;
  wire T726;
  wire T727;
  wire T728;
  wire T729;
  wire T730;
  wire T731;
  wire[1:0] T732;
  wire[1:0] T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire T738;
  wire T739;
  wire[1:0] T740;
  wire[1:0] T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire[1:0] T748;
  wire[1:0] T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire[1:0] T756;
  wire[1:0] T757;
  wire T758;
  wire T759;
  wire T760;
  wire[1:0] T761;
  wire[1:0] T762;
  wire[1:0] T763;
  wire[2:0] T764;
  wire[2:0] T765;
  wire T766;
  wire T767;
  wire T768;
  wire[1:0] T769;
  wire[1:0] T770;
  wire[1:0] T771;
  wire[2:0] T772;
  wire[2:0] T773;
  wire T774;
  wire T775;
  wire T776;
  wire[1:0] T777;
  wire[1:0] T778;
  wire[1:0] T779;
  wire[2:0] T780;
  wire[2:0] T781;
  wire T782;
  wire T783;
  wire T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[2:0] T788;
  wire[2:0] T789;
  wire T790;
  wire T791;
  wire T792;
  wire[1:0] T793;
  wire[1:0] T794;
  wire[1:0] T795;
  wire[2:0] T796;
  wire[2:0] T797;
  wire T798;
  wire T799;
  wire T800;
  wire[1:0] T801;
  wire[1:0] T802;
  wire[1:0] T803;
  wire[2:0] T804;
  wire[2:0] T805;
  wire T806;
  wire T807;
  wire T808;
  wire[1:0] T809;
  wire[1:0] T810;
  wire[1:0] T811;
  wire[2:0] T812;
  wire[2:0] T813;
  wire T814;
  wire T815;
  wire T816;
  wire[1:0] T817;
  wire[1:0] T818;
  wire[1:0] T819;
  wire[2:0] T820;
  wire[2:0] T821;
  wire T822;
  wire T823;
  wire T824;
  wire[1:0] T825;
  wire[1:0] T826;
  wire[1:0] T827;
  wire[2:0] T828;
  wire[2:0] T829;
  wire T830;
  wire T831;
  wire T832;
  wire[1:0] T833;
  wire[1:0] T834;
  wire[1:0] T835;
  wire[2:0] T836;
  wire[2:0] T837;
  wire T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[1:0] T844;
  wire[1:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire[1:0] T852;
  wire[1:0] T853;
  wire T854;
  wire T855;
  wire T856;
  wire T857;
  wire T858;
  wire T859;
  wire[1:0] T860;
  wire[1:0] T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire[1:0] T868;
  wire[1:0] T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire[1:0] T876;
  wire[1:0] T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire[1:0] T884;
  wire[1:0] T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire[1:0] T892;
  wire[1:0] T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire[1:0] T900;
  wire[1:0] T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire[1:0] T908;
  wire[1:0] T909;
  wire T910;
  wire T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire[1:0] T916;
  wire[1:0] T917;
  wire T918;
  wire T919;
  wire T920;
  wire[1:0] T921;
  wire[1:0] T922;
  wire[1:0] T923;
  wire[2:0] T924;
  wire[2:0] T925;
  wire T926;
  wire T927;
  wire T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[2:0] T932;
  wire[2:0] T933;
  wire T934;
  wire T935;
  wire T936;
  wire[1:0] T937;
  wire[1:0] T938;
  wire[1:0] T939;
  wire[2:0] T940;
  wire[2:0] T941;
  wire T942;
  wire T943;
  wire T944;
  wire[1:0] T945;
  wire[1:0] T946;
  wire[1:0] T947;
  wire[2:0] T948;
  wire[2:0] T949;
  wire T950;
  wire T951;
  wire T952;
  wire[1:0] T953;
  wire[1:0] T954;
  wire[1:0] T955;
  wire[2:0] T956;
  wire[2:0] T957;
  wire T958;
  wire T959;
  wire T960;
  wire[1:0] T961;
  wire[1:0] T962;
  wire[1:0] T963;
  wire[2:0] T964;
  wire[2:0] T965;
  wire T966;
  wire T967;
  wire T968;
  wire[1:0] T969;
  wire[1:0] T970;
  wire[1:0] T971;
  wire[2:0] T972;
  wire[2:0] T973;
  wire T974;
  wire T975;
  wire T976;
  wire[1:0] T977;
  wire[1:0] T978;
  wire[1:0] T979;
  wire[2:0] T980;
  wire[2:0] T981;
  wire T982;
  wire T983;
  wire T984;
  wire[1:0] T985;
  wire[1:0] T986;
  wire[1:0] T987;
  wire[2:0] T988;
  wire[2:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire[1:0] T993;
  wire[1:0] T994;
  wire[1:0] T995;
  wire[2:0] T996;
  wire[2:0] T997;
  wire T998;
  wire T999;
  wire T1000;
  wire T1001;
  wire T1002;
  wire T1003;
  wire[1:0] T1004;
  wire[1:0] T1005;
  wire T1006;
  wire T1007;
  wire T1008;
  wire T1009;
  wire T1010;
  wire T1011;
  wire[1:0] T1012;
  wire[1:0] T1013;
  wire T1014;
  wire T1015;
  wire T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire[1:0] T1020;
  wire[1:0] T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire T1026;
  wire T1027;
  wire[1:0] T1028;
  wire[1:0] T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire[1:0] T1036;
  wire[1:0] T1037;
  wire T1038;
  wire T1039;
  wire T1040;
  wire T1041;
  wire T1042;
  wire T1043;
  wire[1:0] T1044;
  wire[1:0] T1045;
  wire T1046;
  wire T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire[1:0] T1052;
  wire[1:0] T1053;
  wire T1054;
  wire T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire[1:0] T1060;
  wire[1:0] T1061;
  wire T1062;
  wire T1063;
  wire T1064;
  wire T1065;
  wire T1066;
  wire T1067;
  wire[1:0] T1068;
  wire[1:0] T1069;
  wire T1070;
  wire T1071;
  wire T1072;
  wire T1073;
  wire T1074;
  wire T1075;
  wire[1:0] T1076;
  wire[1:0] T1077;
  wire T1078;
  wire T1079;
  wire T1080;
  wire[3:0] T1081;
  wire[3:0] T1082;
  wire[3:0] T1083;
  wire[10:0] T1084;
  wire[10:0] T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire[1:0] T1089;
  wire[1:0] T1090;
  wire[1:0] T1091;
  wire[2:0] T1092;
  wire[2:0] T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire[3:0] T1097;
  wire[3:0] T1098;
  wire[3:0] T1099;
  wire[10:0] T1100;
  wire[10:0] T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire[1:0] T1105;
  wire[1:0] T1106;
  wire[1:0] T1107;
  wire[2:0] T1108;
  wire[2:0] T1109;
  wire T1110;
  wire T1111;
  wire T1112;
  wire[3:0] T1113;
  wire[3:0] T1114;
  wire[3:0] T1115;
  wire[10:0] T1116;
  wire[10:0] T1117;
  wire T1118;
  wire T1119;
  wire T1120;
  wire[1:0] T1121;
  wire[1:0] T1122;
  wire[1:0] T1123;
  wire[2:0] T1124;
  wire[2:0] T1125;
  wire T1126;
  wire T1127;
  wire T1128;
  wire[3:0] T1129;
  wire[3:0] T1130;
  wire[3:0] T1131;
  wire[10:0] T1132;
  wire[10:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire[1:0] T1137;
  wire[1:0] T1138;
  wire[1:0] T1139;
  wire[2:0] T1140;
  wire[2:0] T1141;
  wire T1142;
  wire T1143;
  wire T1144;
  wire[3:0] T1145;
  wire[3:0] T1146;
  wire[3:0] T1147;
  wire[10:0] T1148;
  wire[10:0] T1149;
  wire T1150;
  wire T1151;
  wire T1152;
  wire[1:0] T1153;
  wire[1:0] T1154;
  wire[1:0] T1155;
  wire[2:0] T1156;
  wire[2:0] T1157;
  wire T1158;
  wire T1159;
  wire T1160;
  wire[3:0] T1161;
  wire[3:0] T1162;
  wire[3:0] T1163;
  wire[10:0] T1164;
  wire[10:0] T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire[1:0] T1169;
  wire[1:0] T1170;
  wire[1:0] T1171;
  wire[2:0] T1172;
  wire[2:0] T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire[3:0] T1177;
  wire[3:0] T1178;
  wire[3:0] T1179;
  wire[10:0] T1180;
  wire[10:0] T1181;
  wire T1182;
  wire T1183;
  wire T1184;
  wire[1:0] T1185;
  wire[1:0] T1186;
  wire[1:0] T1187;
  wire[2:0] T1188;
  wire[2:0] T1189;
  wire T1190;
  wire T1191;
  wire T1192;
  wire[3:0] T1193;
  wire[3:0] T1194;
  wire[3:0] T1195;
  wire[10:0] T1196;
  wire[10:0] T1197;
  wire T1198;
  wire T1199;
  wire T1200;
  wire[1:0] T1201;
  wire[1:0] T1202;
  wire[1:0] T1203;
  wire[2:0] T1204;
  wire[2:0] T1205;
  wire T1206;
  wire T1207;
  wire T1208;
  wire[3:0] T1209;
  wire[3:0] T1210;
  wire[3:0] T1211;
  wire[10:0] T1212;
  wire[10:0] T1213;
  wire T1214;
  wire T1215;
  wire T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[2:0] T1220;
  wire[2:0] T1221;
  wire T1222;
  wire T1223;
  wire T1224;
  wire[3:0] T1225;
  wire[3:0] T1226;
  wire[3:0] T1227;
  wire[10:0] T1228;
  wire[10:0] T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire[1:0] T1233;
  wire[1:0] T1234;
  wire[1:0] T1235;
  wire[2:0] T1236;
  wire[2:0] T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire[3:0] T1241;
  wire[3:0] T1242;
  wire[3:0] T1243;
  wire[10:0] T1244;
  wire[10:0] T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[1:0] T1252;
  wire[1:0] T1253;
  wire T1254;
  wire T1255;
  wire T1256;
  wire[3:0] T1257;
  wire[3:0] T1258;
  wire[3:0] T1259;
  wire[10:0] T1260;
  wire[10:0] T1261;
  wire T1262;
  wire T1263;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[1:0] T1268;
  wire[1:0] T1269;
  wire T1270;
  wire T1271;
  wire T1272;
  wire[3:0] T1273;
  wire[3:0] T1274;
  wire[3:0] T1275;
  wire[10:0] T1276;
  wire[10:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire[1:0] T1284;
  wire[1:0] T1285;
  wire T1286;
  wire T1287;
  wire T1288;
  wire[3:0] T1289;
  wire[3:0] T1290;
  wire[3:0] T1291;
  wire[10:0] T1292;
  wire[10:0] T1293;
  wire T1294;
  wire T1295;
  wire T1296;
  wire T1297;
  wire T1298;
  wire T1299;
  wire[1:0] T1300;
  wire[1:0] T1301;
  wire T1302;
  wire T1303;
  wire T1304;
  wire[3:0] T1305;
  wire[3:0] T1306;
  wire[3:0] T1307;
  wire[10:0] T1308;
  wire[10:0] T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire T1314;
  wire T1315;
  wire[1:0] T1316;
  wire[1:0] T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire[3:0] T1321;
  wire[3:0] T1322;
  wire[3:0] T1323;
  wire[10:0] T1324;
  wire[10:0] T1325;
  wire T1326;
  wire T1327;
  wire T1328;
  wire T1329;
  wire T1330;
  wire T1331;
  wire[1:0] T1332;
  wire[1:0] T1333;
  wire T1334;
  wire T1335;
  wire T1336;
  wire[3:0] T1337;
  wire[3:0] T1338;
  wire[3:0] T1339;
  wire[10:0] T1340;
  wire[10:0] T1341;
  wire T1342;
  wire T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire[1:0] T1348;
  wire[1:0] T1349;
  wire T1350;
  wire T1351;
  wire T1352;
  wire[3:0] T1353;
  wire[3:0] T1354;
  wire[3:0] T1355;
  wire[10:0] T1356;
  wire[10:0] T1357;
  wire T1358;
  wire T1359;
  wire T1360;
  wire T1361;
  wire T1362;
  wire T1363;
  wire[1:0] T1364;
  wire[1:0] T1365;
  wire T1366;
  wire T1367;
  wire T1368;
  wire[3:0] T1369;
  wire[3:0] T1370;
  wire[3:0] T1371;
  wire[10:0] T1372;
  wire[10:0] T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire[1:0] T1380;
  wire[1:0] T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire[3:0] T1385;
  wire[3:0] T1386;
  wire[3:0] T1387;
  wire[10:0] T1388;
  wire[10:0] T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[1:0] T1396;
  wire[1:0] T1397;
  wire[32:0] T1398;
  wire[32:0] T1399;
  wire[31:0] T1400;
  wire[31:0] T1401;
  wire[30:0] T1402;
  wire[30:0] T1403;
  wire[29:0] T1404;
  wire[29:0] T1405;
  wire[28:0] T1406;
  wire[28:0] T1407;
  wire[27:0] T1408;
  wire[27:0] T1409;
  wire[26:0] T1410;
  wire[26:0] T1411;
  wire[25:0] T1412;
  wire[25:0] T1413;
  wire[24:0] T1414;
  wire[24:0] T1415;
  wire[23:0] T1416;
  wire[23:0] T1417;
  wire[22:0] T1418;
  wire[22:0] T1419;
  wire[21:0] T1420;
  wire[21:0] T1421;
  wire[20:0] T1422;
  wire[20:0] T1423;
  wire[19:0] T1424;
  wire[19:0] T1425;
  wire[18:0] T1426;
  wire[18:0] T1427;
  wire[17:0] T1428;
  wire[17:0] T1429;
  wire[16:0] T1430;
  wire[16:0] T1431;
  wire[15:0] T1432;
  wire[15:0] T1433;
  wire[14:0] T1434;
  wire[14:0] T1435;
  wire[13:0] T1436;
  wire[13:0] T1437;
  wire[12:0] T1438;
  wire[12:0] T1439;
  wire[11:0] T1440;
  wire[11:0] T1441;
  wire[10:0] T1442;
  wire[10:0] T1443;
  wire[9:0] T1444;
  wire[9:0] T1445;
  wire[8:0] T1446;
  wire[8:0] T1447;
  wire[7:0] T1448;
  wire[7:0] T1449;
  wire[6:0] T1450;
  wire[6:0] T1451;
  wire[5:0] T1452;
  wire[5:0] T1453;
  wire[4:0] T1454;
  wire[4:0] T1455;
  wire[3:0] T1456;
  wire[3:0] T1457;
  wire[2:0] T1458;
  wire[2:0] T1459;
  wire[1:0] T1460;
  wire[1:0] T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire[3:0] T1465;
  wire[3:0] T1466;
  wire[3:0] T1467;
  wire[15:0] T1468;
  wire[15:0] T1469;
  wire T1470;
  wire T1471;
  wire T1472;
  wire[3:0] T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[15:0] T1476;
  wire[15:0] T1477;
  wire T1478;
  wire T1479;
  wire T1480;
  wire[3:0] T1481;
  wire[3:0] T1482;
  wire[3:0] T1483;
  wire[15:0] T1484;
  wire[15:0] T1485;
  wire T1486;
  wire T1487;
  wire T1488;
  wire[3:0] T1489;
  wire[3:0] T1490;
  wire[3:0] T1491;
  wire[15:0] T1492;
  wire[15:0] T1493;
  wire T1494;
  wire T1495;
  wire T1496;
  wire[3:0] T1497;
  wire[3:0] T1498;
  wire[3:0] T1499;
  wire[15:0] T1500;
  wire[15:0] T1501;
  wire T1502;
  wire T1503;
  wire T1504;
  wire[3:0] T1505;
  wire[3:0] T1506;
  wire[3:0] T1507;
  wire[15:0] T1508;
  wire[15:0] T1509;
  wire T1510;
  wire T1511;
  wire T1512;
  wire[3:0] T1513;
  wire[3:0] T1514;
  wire[3:0] T1515;
  wire[15:0] T1516;
  wire[15:0] T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire[3:0] T1521;
  wire[3:0] T1522;
  wire[3:0] T1523;
  wire[15:0] T1524;
  wire[15:0] T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire[3:0] T1529;
  wire[3:0] T1530;
  wire[3:0] T1531;
  wire[15:0] T1532;
  wire[15:0] T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire[3:0] T1537;
  wire[3:0] T1538;
  wire[3:0] T1539;
  wire[15:0] T1540;
  wire[15:0] T1541;
  wire T1542;
  wire T1543;
  wire T1544;
  wire[3:0] T1545;
  wire[3:0] T1546;
  wire[3:0] T1547;
  wire[15:0] T1548;
  wire[15:0] T1549;
  wire T1550;
  wire T1551;
  wire T1552;
  wire[3:0] T1553;
  wire[3:0] T1554;
  wire[3:0] T1555;
  wire[15:0] T1556;
  wire[15:0] T1557;
  wire T1558;
  wire T1559;
  wire T1560;
  wire[3:0] T1561;
  wire[3:0] T1562;
  wire[3:0] T1563;
  wire[15:0] T1564;
  wire[15:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire[3:0] T1569;
  wire[3:0] T1570;
  wire[3:0] T1571;
  wire[15:0] T1572;
  wire[15:0] T1573;
  wire T1574;
  wire T1575;
  wire T1576;
  wire[3:0] T1577;
  wire[3:0] T1578;
  wire[3:0] T1579;
  wire[15:0] T1580;
  wire[15:0] T1581;
  wire T1582;
  wire T1583;
  wire T1584;
  wire[3:0] T1585;
  wire[3:0] T1586;
  wire[3:0] T1587;
  wire[15:0] T1588;
  wire[15:0] T1589;
  wire T1590;
  wire T1591;
  wire T1592;
  wire[3:0] T1593;
  wire[3:0] T1594;
  wire[3:0] T1595;
  wire[15:0] T1596;
  wire[15:0] T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire[3:0] T1601;
  wire[3:0] T1602;
  wire[3:0] T1603;
  wire[15:0] T1604;
  wire[15:0] T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire[3:0] T1609;
  wire[3:0] T1610;
  wire[3:0] T1611;
  wire[15:0] T1612;
  wire[15:0] T1613;
  wire T1614;
  wire T1615;
  wire T1616;
  wire[3:0] T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[15:0] T1620;
  wire[15:0] T1621;
  wire T1622;
  wire T1623;
  wire T1624;
  wire[3:0] T1625;
  wire[3:0] T1626;
  wire[3:0] T1627;
  wire[15:0] T1628;
  wire[15:0] T1629;
  wire T1630;
  wire T1631;
  wire T1632;
  wire[3:0] T1633;
  wire[3:0] T1634;
  wire[3:0] T1635;
  wire[15:0] T1636;
  wire[15:0] T1637;
  wire T1638;
  wire T1639;
  wire T1640;
  wire[3:0] T1641;
  wire[3:0] T1642;
  wire[3:0] T1643;
  wire[15:0] T1644;
  wire[15:0] T1645;
  wire T1646;
  wire T1647;
  wire T1648;
  wire[3:0] T1649;
  wire[3:0] T1650;
  wire[3:0] T1651;
  wire[15:0] T1652;
  wire[15:0] T1653;
  wire T1654;
  wire T1655;
  wire T1656;
  wire[3:0] T1657;
  wire[3:0] T1658;
  wire[3:0] T1659;
  wire[15:0] T1660;
  wire[15:0] T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire[3:0] T1665;
  wire[3:0] T1666;
  wire[3:0] T1667;
  wire[15:0] T1668;
  wire[15:0] T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire[3:0] T1673;
  wire[3:0] T1674;
  wire[3:0] T1675;
  wire[15:0] T1676;
  wire[15:0] T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire[3:0] T1681;
  wire[3:0] T1682;
  wire[3:0] T1683;
  wire[15:0] T1684;
  wire[15:0] T1685;
  wire T1686;
  wire T1687;
  wire T1688;
  wire[3:0] T1689;
  wire[3:0] T1690;
  wire[3:0] T1691;
  wire[15:0] T1692;
  wire[15:0] T1693;
  wire T1694;
  wire T1695;
  wire T1696;
  wire[3:0] T1697;
  wire[3:0] T1698;
  wire[3:0] T1699;
  wire[15:0] T1700;
  wire[15:0] T1701;
  wire T1702;
  wire T1703;
  wire T1704;
  wire[3:0] T1705;
  wire[3:0] T1706;
  wire[3:0] T1707;
  wire[15:0] T1708;
  wire[15:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire[3:0] T1713;
  wire[3:0] T1714;
  wire[3:0] T1715;
  wire[15:0] T1716;
  wire[15:0] T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire[3:0] T1721;
  wire[3:0] T1722;
  wire[3:0] T1723;
  wire[15:0] T1724;
  wire[15:0] T1725;

  assign io_chanxy_out = T0;
  assign T0 = T1;
  assign T1 = {T1390, T2};
  assign T2 = T3;
  assign T3 = {T1382, T4};
  assign T4 = T5;
  assign T5 = {T1374, T6};
  assign T6 = T7;
  assign T7 = {T1366, T8};
  assign T8 = T9;
  assign T9 = {T1358, T10};
  assign T10 = T11;
  assign T11 = {T1350, T12};
  assign T12 = T13;
  assign T13 = {T1342, T14};
  assign T14 = T15;
  assign T15 = {T1334, T16};
  assign T16 = T17;
  assign T17 = {T1326, T18};
  assign T18 = T19;
  assign T19 = {T1318, T20};
  assign T20 = T21;
  assign T21 = {T1310, T22};
  assign T22 = T23;
  assign T23 = {T1302, T24};
  assign T24 = T25;
  assign T25 = {T1294, T26};
  assign T26 = T27;
  assign T27 = {T1286, T28};
  assign T28 = T29;
  assign T29 = {T1278, T30};
  assign T30 = T31;
  assign T31 = {T1270, T32};
  assign T32 = T33;
  assign T33 = {T1262, T34};
  assign T34 = T35;
  assign T35 = {T1254, T36};
  assign T36 = T37;
  assign T37 = {T1246, T38};
  assign T38 = T39;
  assign T39 = {T1238, T40};
  assign T40 = T41;
  assign T41 = {T1230, T42};
  assign T42 = T43;
  assign T43 = {T1222, T44};
  assign T44 = T45;
  assign T45 = {T1214, T46};
  assign T46 = T47;
  assign T47 = {T1206, T48};
  assign T48 = T49;
  assign T49 = {T1198, T50};
  assign T50 = T51;
  assign T51 = {T1190, T52};
  assign T52 = T53;
  assign T53 = {T1182, T54};
  assign T54 = T55;
  assign T55 = {T1174, T56};
  assign T56 = T57;
  assign T57 = {T1166, T58};
  assign T58 = T59;
  assign T59 = {T1158, T60};
  assign T60 = T61;
  assign T61 = {T1150, T62};
  assign T62 = T63;
  assign T63 = {T1142, T64};
  assign T64 = T65;
  assign T65 = {T1134, T66};
  assign T66 = T67;
  assign T67 = {T1126, T68};
  assign T68 = T69;
  assign T69 = {T1118, T70};
  assign T70 = T71;
  assign T71 = {T1110, T72};
  assign T72 = T73;
  assign T73 = {T1102, T74};
  assign T74 = T75;
  assign T75 = {T1094, T76};
  assign T76 = T77;
  assign T77 = {T1086, T78};
  assign T78 = T79;
  assign T79 = {T1078, T80};
  assign T80 = T81;
  assign T81 = {T1070, T82};
  assign T82 = T83;
  assign T83 = {T1062, T84};
  assign T84 = T85;
  assign T85 = {T1054, T86};
  assign T86 = T87;
  assign T87 = {T1046, T88};
  assign T88 = T89;
  assign T89 = {T1038, T90};
  assign T90 = T91;
  assign T91 = {T1030, T92};
  assign T92 = T93;
  assign T93 = {T1022, T94};
  assign T94 = T95;
  assign T95 = {T1014, T96};
  assign T96 = T97;
  assign T97 = {T1006, T98};
  assign T98 = T99;
  assign T99 = {T998, T100};
  assign T100 = T101;
  assign T101 = {T990, T102};
  assign T102 = T103;
  assign T103 = {T982, T104};
  assign T104 = T105;
  assign T105 = {T974, T106};
  assign T106 = T107;
  assign T107 = {T966, T108};
  assign T108 = T109;
  assign T109 = {T958, T110};
  assign T110 = T111;
  assign T111 = {T950, T112};
  assign T112 = T113;
  assign T113 = {T942, T114};
  assign T114 = T115;
  assign T115 = {T934, T116};
  assign T116 = T117;
  assign T117 = {T926, T118};
  assign T118 = T119;
  assign T119 = {T918, T120};
  assign T120 = T121;
  assign T121 = {T910, T122};
  assign T122 = T123;
  assign T123 = {T902, T124};
  assign T124 = T125;
  assign T125 = {T894, T126};
  assign T126 = T127;
  assign T127 = {T886, T128};
  assign T128 = T129;
  assign T129 = {T878, T130};
  assign T130 = T131;
  assign T131 = {T870, T132};
  assign T132 = T133;
  assign T133 = {T862, T134};
  assign T134 = T135;
  assign T135 = {T854, T136};
  assign T136 = T137;
  assign T137 = {T846, T138};
  assign T138 = T139;
  assign T139 = {T838, T140};
  assign T140 = T141;
  assign T141 = {T830, T142};
  assign T142 = T143;
  assign T143 = {T822, T144};
  assign T144 = T145;
  assign T145 = {T814, T146};
  assign T146 = T147;
  assign T147 = {T806, T148};
  assign T148 = T149;
  assign T149 = {T798, T150};
  assign T150 = T151;
  assign T151 = {T790, T152};
  assign T152 = T153;
  assign T153 = {T782, T154};
  assign T154 = T155;
  assign T155 = {T774, T156};
  assign T156 = T157;
  assign T157 = {T766, T158};
  assign T158 = T159;
  assign T159 = {T758, T160};
  assign T160 = T161;
  assign T161 = {T750, T162};
  assign T162 = T163;
  assign T163 = {T742, T164};
  assign T164 = T165;
  assign T165 = {T734, T166};
  assign T166 = T167;
  assign T167 = {T726, T168};
  assign T168 = T169;
  assign T169 = {T718, T170};
  assign T170 = T171;
  assign T171 = {T710, T172};
  assign T172 = T173;
  assign T173 = {T702, T174};
  assign T174 = T175;
  assign T175 = {T694, T176};
  assign T176 = T177;
  assign T177 = {T686, T178};
  assign T178 = T179;
  assign T179 = {T678, T180};
  assign T180 = T181;
  assign T181 = {T670, T182};
  assign T182 = T183;
  assign T183 = {T662, T184};
  assign T184 = T185;
  assign T185 = {T654, T186};
  assign T186 = T187;
  assign T187 = {T646, T188};
  assign T188 = T189;
  assign T189 = {T638, T190};
  assign T190 = T191;
  assign T191 = {T630, T192};
  assign T192 = T193;
  assign T193 = {T622, T194};
  assign T194 = T195;
  assign T195 = {T614, T196};
  assign T196 = T197;
  assign T197 = {T606, T198};
  assign T198 = T199;
  assign T199 = {T598, T200};
  assign T200 = T201;
  assign T201 = {T590, T202};
  assign T202 = T203;
  assign T203 = {T582, T204};
  assign T204 = T205;
  assign T205 = {T574, T206};
  assign T206 = T207;
  assign T207 = {T566, T208};
  assign T208 = T209;
  assign T209 = {T558, T210};
  assign T210 = T211;
  assign T211 = {T550, T212};
  assign T212 = T213;
  assign T213 = {T542, T214};
  assign T214 = T215;
  assign T215 = {T534, T216};
  assign T216 = T217;
  assign T217 = {T526, T218};
  assign T218 = T219;
  assign T219 = {T518, T220};
  assign T220 = T221;
  assign T221 = {T510, T222};
  assign T222 = T223;
  assign T223 = {T502, T224};
  assign T224 = T225;
  assign T225 = {T494, T226};
  assign T226 = T227;
  assign T227 = {T486, T228};
  assign T228 = T229;
  assign T229 = {T478, T230};
  assign T230 = T231;
  assign T231 = {T470, T232};
  assign T232 = T233;
  assign T233 = {T462, T234};
  assign T234 = T235;
  assign T235 = {T454, T236};
  assign T236 = T237;
  assign T237 = {T446, T238};
  assign T238 = T239;
  assign T239 = {T438, T240};
  assign T240 = T241;
  assign T241 = {T430, T242};
  assign T242 = T243;
  assign T243 = {T422, T244};
  assign T244 = T245;
  assign T245 = {T414, T246};
  assign T246 = T247;
  assign T247 = {T406, T248};
  assign T248 = T249;
  assign T249 = {T398, T250};
  assign T250 = T251;
  assign T251 = {T390, T252};
  assign T252 = T253;
  assign T253 = {T382, T254};
  assign T254 = T255;
  assign T255 = {T374, T256};
  assign T256 = T257;
  assign T257 = {T366, T258};
  assign T258 = T259;
  assign T259 = {T358, T260};
  assign T260 = T261;
  assign T261 = {T350, T262};
  assign T262 = T263;
  assign T263 = {T342, T264};
  assign T264 = T265;
  assign T265 = {T334, T266};
  assign T266 = T267;
  assign T267 = {T326, T268};
  assign T268 = T269;
  assign T269 = {T318, T270};
  assign T270 = T271;
  assign T271 = {T310, T272};
  assign T272 = T273;
  assign T273 = {T302, T274};
  assign T274 = T275;
  assign T275 = {T294, T276};
  assign T276 = T277;
  assign T277 = {T286, T278};
  assign T278 = T279;
  assign T279 = T280;
  assign T280 = T284[T281];
  assign T281 = T282;
  assign T282 = T283;
  assign T283 = io_chanxy_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T284 = T285;
  assign T285 = io_chanxy_in[4'h8/* 8*/:1'h0/* 0*/];
  assign T286 = T287;
  assign T287 = T288;
  assign T288 = T292[T289];
  assign T289 = T290;
  assign T290 = T291;
  assign T291 = io_chanxy_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T292 = T293;
  assign T293 = io_chanxy_in[5'h11/* 17*/:4'h9/* 9*/];
  assign T294 = T295;
  assign T295 = T296;
  assign T296 = T300[T297];
  assign T297 = T298;
  assign T298 = T299;
  assign T299 = io_chanxy_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T300 = T301;
  assign T301 = io_chanxy_in[5'h1a/* 26*/:5'h12/* 18*/];
  assign T302 = T303;
  assign T303 = T304;
  assign T304 = T308[T305];
  assign T305 = T306;
  assign T306 = T307;
  assign T307 = io_chanxy_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T308 = T309;
  assign T309 = io_chanxy_in[6'h23/* 35*/:5'h1b/* 27*/];
  assign T310 = T311;
  assign T311 = T312;
  assign T312 = T316[T313];
  assign T313 = T314;
  assign T314 = T315;
  assign T315 = io_chanxy_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T316 = T317;
  assign T317 = io_chanxy_in[6'h2c/* 44*/:6'h24/* 36*/];
  assign T318 = T319;
  assign T319 = T320;
  assign T320 = T324[T321];
  assign T321 = T322;
  assign T322 = T323;
  assign T323 = io_chanxy_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T324 = T325;
  assign T325 = io_chanxy_in[6'h35/* 53*/:6'h2d/* 45*/];
  assign T326 = T327;
  assign T327 = T328;
  assign T328 = T332[T329];
  assign T329 = T330;
  assign T330 = T331;
  assign T331 = io_chanxy_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T332 = T333;
  assign T333 = io_chanxy_in[6'h3e/* 62*/:6'h36/* 54*/];
  assign T334 = T335;
  assign T335 = T336;
  assign T336 = T340[T337];
  assign T337 = T338;
  assign T338 = T339;
  assign T339 = io_chanxy_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T340 = T341;
  assign T341 = io_chanxy_in[7'h47/* 71*/:6'h3f/* 63*/];
  assign T342 = T343;
  assign T343 = T344;
  assign T344 = T348[T345];
  assign T345 = T346;
  assign T346 = T347;
  assign T347 = io_chanxy_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T348 = T349;
  assign T349 = io_chanxy_in[7'h50/* 80*/:7'h48/* 72*/];
  assign T350 = T351;
  assign T351 = T352;
  assign T352 = T356[T353];
  assign T353 = T354;
  assign T354 = T355;
  assign T355 = io_chanxy_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T356 = T357;
  assign T357 = io_chanxy_in[7'h59/* 89*/:7'h51/* 81*/];
  assign T358 = T359;
  assign T359 = T360;
  assign T360 = T364[T361];
  assign T361 = T362;
  assign T362 = T363;
  assign T363 = io_chanxy_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T364 = T365;
  assign T365 = io_chanxy_in[7'h62/* 98*/:7'h5a/* 90*/];
  assign T366 = T367;
  assign T367 = T368;
  assign T368 = T372[T369];
  assign T369 = T370;
  assign T370 = T371;
  assign T371 = io_chanxy_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T372 = T373;
  assign T373 = io_chanxy_in[7'h6b/* 107*/:7'h63/* 99*/];
  assign T374 = T375;
  assign T375 = T376;
  assign T376 = T380[T377];
  assign T377 = T378;
  assign T378 = T379;
  assign T379 = io_chanxy_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T380 = T381;
  assign T381 = io_chanxy_in[7'h74/* 116*/:7'h6c/* 108*/];
  assign T382 = T383;
  assign T383 = T384;
  assign T384 = T388[T385];
  assign T385 = T386;
  assign T386 = T387;
  assign T387 = io_chanxy_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T388 = T389;
  assign T389 = io_chanxy_in[7'h7d/* 125*/:7'h75/* 117*/];
  assign T390 = T391;
  assign T391 = T392;
  assign T392 = T396[T393];
  assign T393 = T394;
  assign T394 = T395;
  assign T395 = io_chanxy_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T396 = T397;
  assign T397 = io_chanxy_in[8'h86/* 134*/:7'h7e/* 126*/];
  assign T398 = T399;
  assign T399 = T400;
  assign T400 = T404[T401];
  assign T401 = T402;
  assign T402 = T403;
  assign T403 = io_chanxy_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T404 = T405;
  assign T405 = io_chanxy_in[8'h8f/* 143*/:8'h87/* 135*/];
  assign T406 = T407;
  assign T407 = T408;
  assign T408 = T412[T409];
  assign T409 = T410;
  assign T410 = T411;
  assign T411 = io_chanxy_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T412 = T413;
  assign T413 = io_chanxy_in[8'h98/* 152*/:8'h90/* 144*/];
  assign T414 = T415;
  assign T415 = T416;
  assign T416 = T420[T417];
  assign T417 = T418;
  assign T418 = T419;
  assign T419 = io_chanxy_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T420 = T421;
  assign T421 = io_chanxy_in[8'ha1/* 161*/:8'h99/* 153*/];
  assign T422 = T423;
  assign T423 = T424;
  assign T424 = T428[T425];
  assign T425 = T426;
  assign T426 = T427;
  assign T427 = io_chanxy_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T428 = T429;
  assign T429 = io_chanxy_in[8'haa/* 170*/:8'ha2/* 162*/];
  assign T430 = T431;
  assign T431 = T432;
  assign T432 = T436[T433];
  assign T433 = T434;
  assign T434 = T435;
  assign T435 = io_chanxy_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T436 = T437;
  assign T437 = io_chanxy_in[8'hb3/* 179*/:8'hab/* 171*/];
  assign T438 = T439;
  assign T439 = T440;
  assign T440 = T444[T441];
  assign T441 = T442;
  assign T442 = T443;
  assign T443 = io_chanxy_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T444 = T445;
  assign T445 = io_chanxy_in[8'hbc/* 188*/:8'hb4/* 180*/];
  assign T446 = T447;
  assign T447 = T448;
  assign T448 = T452[T449];
  assign T449 = T450;
  assign T450 = T451;
  assign T451 = io_chanxy_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T452 = T453;
  assign T453 = io_chanxy_in[8'hc5/* 197*/:8'hbd/* 189*/];
  assign T454 = T455;
  assign T455 = T456;
  assign T456 = T460[T457];
  assign T457 = T458;
  assign T458 = T459;
  assign T459 = io_chanxy_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T460 = T461;
  assign T461 = io_chanxy_in[8'hce/* 206*/:8'hc6/* 198*/];
  assign T462 = T463;
  assign T463 = T464;
  assign T464 = T468[T465];
  assign T465 = T466;
  assign T466 = T467;
  assign T467 = io_chanxy_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T468 = T469;
  assign T469 = io_chanxy_in[8'hd7/* 215*/:8'hcf/* 207*/];
  assign T470 = T471;
  assign T471 = T472;
  assign T472 = T476[T473];
  assign T473 = T474;
  assign T474 = T475;
  assign T475 = io_chanxy_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T476 = T477;
  assign T477 = io_chanxy_in[8'he0/* 224*/:8'hd8/* 216*/];
  assign T478 = T479;
  assign T479 = T480;
  assign T480 = T484[T481];
  assign T481 = T482;
  assign T482 = T483;
  assign T483 = io_chanxy_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T484 = T485;
  assign T485 = io_chanxy_in[8'he9/* 233*/:8'he1/* 225*/];
  assign T486 = T487;
  assign T487 = T488;
  assign T488 = T492[T489];
  assign T489 = T490;
  assign T490 = T491;
  assign T491 = io_chanxy_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T492 = T493;
  assign T493 = io_chanxy_in[8'hf2/* 242*/:8'hea/* 234*/];
  assign T494 = T495;
  assign T495 = T496;
  assign T496 = T500[T497];
  assign T497 = T498;
  assign T498 = T499;
  assign T499 = io_chanxy_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T500 = T501;
  assign T501 = io_chanxy_in[8'hfb/* 251*/:8'hf3/* 243*/];
  assign T502 = T503;
  assign T503 = T504;
  assign T504 = T508[T505];
  assign T505 = T506;
  assign T506 = T507;
  assign T507 = io_chanxy_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T508 = T509;
  assign T509 = io_chanxy_in[9'h104/* 260*/:8'hfc/* 252*/];
  assign T510 = T511;
  assign T511 = T512;
  assign T512 = T516[T513];
  assign T513 = T514;
  assign T514 = T515;
  assign T515 = io_chanxy_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T516 = T517;
  assign T517 = io_chanxy_in[9'h10d/* 269*/:9'h105/* 261*/];
  assign T518 = T519;
  assign T519 = T520;
  assign T520 = T524[T521];
  assign T521 = T522;
  assign T522 = T523;
  assign T523 = io_chanxy_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T524 = T525;
  assign T525 = io_chanxy_in[9'h116/* 278*/:9'h10e/* 270*/];
  assign T526 = T527;
  assign T527 = T528;
  assign T528 = T532[T529];
  assign T529 = T530;
  assign T530 = T531;
  assign T531 = io_chanxy_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T532 = T533;
  assign T533 = io_chanxy_in[9'h11f/* 287*/:9'h117/* 279*/];
  assign T534 = T535;
  assign T535 = T536;
  assign T536 = T540[T537];
  assign T537 = T538;
  assign T538 = T539;
  assign T539 = io_chanxy_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T540 = T541;
  assign T541 = io_chanxy_in[9'h128/* 296*/:9'h120/* 288*/];
  assign T542 = T543;
  assign T543 = T544;
  assign T544 = T548[T545];
  assign T545 = T546;
  assign T546 = T547;
  assign T547 = io_chanxy_config[8'h87/* 135*/:8'h84/* 132*/];
  assign T548 = T549;
  assign T549 = io_chanxy_in[9'h131/* 305*/:9'h129/* 297*/];
  assign T550 = T551;
  assign T551 = T552;
  assign T552 = T556[T553];
  assign T553 = T554;
  assign T554 = T555;
  assign T555 = io_chanxy_config[8'h8b/* 139*/:8'h88/* 136*/];
  assign T556 = T557;
  assign T557 = io_chanxy_in[9'h13a/* 314*/:9'h132/* 306*/];
  assign T558 = T559;
  assign T559 = T560;
  assign T560 = T564[T561];
  assign T561 = T562;
  assign T562 = T563;
  assign T563 = io_chanxy_config[8'h8f/* 143*/:8'h8c/* 140*/];
  assign T564 = T565;
  assign T565 = io_chanxy_in[9'h143/* 323*/:9'h13b/* 315*/];
  assign T566 = T567;
  assign T567 = T568;
  assign T568 = T572[T569];
  assign T569 = T570;
  assign T570 = T571;
  assign T571 = io_chanxy_config[8'h93/* 147*/:8'h90/* 144*/];
  assign T572 = T573;
  assign T573 = io_chanxy_in[9'h14c/* 332*/:9'h144/* 324*/];
  assign T574 = T575;
  assign T575 = T576;
  assign T576 = T580[T577];
  assign T577 = T578;
  assign T578 = T579;
  assign T579 = io_chanxy_config[8'h97/* 151*/:8'h94/* 148*/];
  assign T580 = T581;
  assign T581 = io_chanxy_in[9'h155/* 341*/:9'h14d/* 333*/];
  assign T582 = T583;
  assign T583 = T584;
  assign T584 = T588[T585];
  assign T585 = T586;
  assign T586 = T587;
  assign T587 = io_chanxy_config[8'h9b/* 155*/:8'h98/* 152*/];
  assign T588 = T589;
  assign T589 = io_chanxy_in[9'h15e/* 350*/:9'h156/* 342*/];
  assign T590 = T591;
  assign T591 = T592;
  assign T592 = T596[T593];
  assign T593 = T594;
  assign T594 = T595;
  assign T595 = io_chanxy_config[8'h9f/* 159*/:8'h9c/* 156*/];
  assign T596 = T597;
  assign T597 = io_chanxy_in[9'h167/* 359*/:9'h15f/* 351*/];
  assign T598 = T599;
  assign T599 = T600;
  assign T600 = T604[T601];
  assign T601 = T602;
  assign T602 = T603;
  assign T603 = io_chanxy_config[8'ha1/* 161*/:8'ha0/* 160*/];
  assign T604 = T605;
  assign T605 = io_chanxy_in[9'h16a/* 362*/:9'h168/* 360*/];
  assign T606 = T607;
  assign T607 = T608;
  assign T608 = T612[T609];
  assign T609 = T610;
  assign T610 = T611;
  assign T611 = io_chanxy_config[8'ha3/* 163*/:8'ha2/* 162*/];
  assign T612 = T613;
  assign T613 = io_chanxy_in[9'h16d/* 365*/:9'h16b/* 363*/];
  assign T614 = T615;
  assign T615 = T616;
  assign T616 = T620[T617];
  assign T617 = T618;
  assign T618 = T619;
  assign T619 = io_chanxy_config[8'ha5/* 165*/:8'ha4/* 164*/];
  assign T620 = T621;
  assign T621 = io_chanxy_in[9'h170/* 368*/:9'h16e/* 366*/];
  assign T622 = T623;
  assign T623 = T624;
  assign T624 = T628[T625];
  assign T625 = T626;
  assign T626 = T627;
  assign T627 = io_chanxy_config[8'ha7/* 167*/:8'ha6/* 166*/];
  assign T628 = T629;
  assign T629 = io_chanxy_in[9'h173/* 371*/:9'h171/* 369*/];
  assign T630 = T631;
  assign T631 = T632;
  assign T632 = T636[T633];
  assign T633 = T634;
  assign T634 = T635;
  assign T635 = io_chanxy_config[8'ha9/* 169*/:8'ha8/* 168*/];
  assign T636 = T637;
  assign T637 = io_chanxy_in[9'h176/* 374*/:9'h174/* 372*/];
  assign T638 = T639;
  assign T639 = T640;
  assign T640 = T644[T641];
  assign T641 = T642;
  assign T642 = T643;
  assign T643 = io_chanxy_config[8'hab/* 171*/:8'haa/* 170*/];
  assign T644 = T645;
  assign T645 = io_chanxy_in[9'h179/* 377*/:9'h177/* 375*/];
  assign T646 = T647;
  assign T647 = T648;
  assign T648 = T652[T649];
  assign T649 = T650;
  assign T650 = T651;
  assign T651 = io_chanxy_config[8'had/* 173*/:8'hac/* 172*/];
  assign T652 = T653;
  assign T653 = io_chanxy_in[9'h17c/* 380*/:9'h17a/* 378*/];
  assign T654 = T655;
  assign T655 = T656;
  assign T656 = T660[T657];
  assign T657 = T658;
  assign T658 = T659;
  assign T659 = io_chanxy_config[8'haf/* 175*/:8'hae/* 174*/];
  assign T660 = T661;
  assign T661 = io_chanxy_in[9'h17f/* 383*/:9'h17d/* 381*/];
  assign T662 = T663;
  assign T663 = T664;
  assign T664 = T668[T665];
  assign T665 = T666;
  assign T666 = T667;
  assign T667 = io_chanxy_config[8'hb1/* 177*/:8'hb0/* 176*/];
  assign T668 = T669;
  assign T669 = io_chanxy_in[9'h182/* 386*/:9'h180/* 384*/];
  assign T670 = T671;
  assign T671 = T672;
  assign T672 = T676[T673];
  assign T673 = T674;
  assign T674 = T675;
  assign T675 = io_chanxy_config[8'hb3/* 179*/:8'hb2/* 178*/];
  assign T676 = T677;
  assign T677 = io_chanxy_in[9'h185/* 389*/:9'h183/* 387*/];
  assign T678 = T679;
  assign T679 = T680;
  assign T680 = T684[T681];
  assign T681 = T682;
  assign T682 = T683;
  assign T683 = io_chanxy_config[8'hb4/* 180*/:8'hb4/* 180*/];
  assign T684 = T685;
  assign T685 = io_chanxy_in[9'h187/* 391*/:9'h186/* 390*/];
  assign T686 = T687;
  assign T687 = T688;
  assign T688 = T692[T689];
  assign T689 = T690;
  assign T690 = T691;
  assign T691 = io_chanxy_config[8'hb5/* 181*/:8'hb5/* 181*/];
  assign T692 = T693;
  assign T693 = io_chanxy_in[9'h189/* 393*/:9'h188/* 392*/];
  assign T694 = T695;
  assign T695 = T696;
  assign T696 = T700[T697];
  assign T697 = T698;
  assign T698 = T699;
  assign T699 = io_chanxy_config[8'hb6/* 182*/:8'hb6/* 182*/];
  assign T700 = T701;
  assign T701 = io_chanxy_in[9'h18b/* 395*/:9'h18a/* 394*/];
  assign T702 = T703;
  assign T703 = T704;
  assign T704 = T708[T705];
  assign T705 = T706;
  assign T706 = T707;
  assign T707 = io_chanxy_config[8'hb7/* 183*/:8'hb7/* 183*/];
  assign T708 = T709;
  assign T709 = io_chanxy_in[9'h18d/* 397*/:9'h18c/* 396*/];
  assign T710 = T711;
  assign T711 = T712;
  assign T712 = T716[T713];
  assign T713 = T714;
  assign T714 = T715;
  assign T715 = io_chanxy_config[8'hb8/* 184*/:8'hb8/* 184*/];
  assign T716 = T717;
  assign T717 = io_chanxy_in[9'h18f/* 399*/:9'h18e/* 398*/];
  assign T718 = T719;
  assign T719 = T720;
  assign T720 = T724[T721];
  assign T721 = T722;
  assign T722 = T723;
  assign T723 = io_chanxy_config[8'hb9/* 185*/:8'hb9/* 185*/];
  assign T724 = T725;
  assign T725 = io_chanxy_in[9'h191/* 401*/:9'h190/* 400*/];
  assign T726 = T727;
  assign T727 = T728;
  assign T728 = T732[T729];
  assign T729 = T730;
  assign T730 = T731;
  assign T731 = io_chanxy_config[8'hba/* 186*/:8'hba/* 186*/];
  assign T732 = T733;
  assign T733 = io_chanxy_in[9'h193/* 403*/:9'h192/* 402*/];
  assign T734 = T735;
  assign T735 = T736;
  assign T736 = T740[T737];
  assign T737 = T738;
  assign T738 = T739;
  assign T739 = io_chanxy_config[8'hbb/* 187*/:8'hbb/* 187*/];
  assign T740 = T741;
  assign T741 = io_chanxy_in[9'h195/* 405*/:9'h194/* 404*/];
  assign T742 = T743;
  assign T743 = T744;
  assign T744 = T748[T745];
  assign T745 = T746;
  assign T746 = T747;
  assign T747 = io_chanxy_config[8'hbc/* 188*/:8'hbc/* 188*/];
  assign T748 = T749;
  assign T749 = io_chanxy_in[9'h197/* 407*/:9'h196/* 406*/];
  assign T750 = T751;
  assign T751 = T752;
  assign T752 = T756[T753];
  assign T753 = T754;
  assign T754 = T755;
  assign T755 = io_chanxy_config[8'hbd/* 189*/:8'hbd/* 189*/];
  assign T756 = T757;
  assign T757 = io_chanxy_in[9'h199/* 409*/:9'h198/* 408*/];
  assign T758 = T759;
  assign T759 = T760;
  assign T760 = T764[T761];
  assign T761 = T762;
  assign T762 = T763;
  assign T763 = io_chanxy_config[8'hbf/* 191*/:8'hbe/* 190*/];
  assign T764 = T765;
  assign T765 = io_chanxy_in[9'h19c/* 412*/:9'h19a/* 410*/];
  assign T766 = T767;
  assign T767 = T768;
  assign T768 = T772[T769];
  assign T769 = T770;
  assign T770 = T771;
  assign T771 = io_chanxy_config[8'hc1/* 193*/:8'hc0/* 192*/];
  assign T772 = T773;
  assign T773 = io_chanxy_in[9'h19f/* 415*/:9'h19d/* 413*/];
  assign T774 = T775;
  assign T775 = T776;
  assign T776 = T780[T777];
  assign T777 = T778;
  assign T778 = T779;
  assign T779 = io_chanxy_config[8'hc3/* 195*/:8'hc2/* 194*/];
  assign T780 = T781;
  assign T781 = io_chanxy_in[9'h1a2/* 418*/:9'h1a0/* 416*/];
  assign T782 = T783;
  assign T783 = T784;
  assign T784 = T788[T785];
  assign T785 = T786;
  assign T786 = T787;
  assign T787 = io_chanxy_config[8'hc5/* 197*/:8'hc4/* 196*/];
  assign T788 = T789;
  assign T789 = io_chanxy_in[9'h1a5/* 421*/:9'h1a3/* 419*/];
  assign T790 = T791;
  assign T791 = T792;
  assign T792 = T796[T793];
  assign T793 = T794;
  assign T794 = T795;
  assign T795 = io_chanxy_config[8'hc7/* 199*/:8'hc6/* 198*/];
  assign T796 = T797;
  assign T797 = io_chanxy_in[9'h1a8/* 424*/:9'h1a6/* 422*/];
  assign T798 = T799;
  assign T799 = T800;
  assign T800 = T804[T801];
  assign T801 = T802;
  assign T802 = T803;
  assign T803 = io_chanxy_config[8'hc9/* 201*/:8'hc8/* 200*/];
  assign T804 = T805;
  assign T805 = io_chanxy_in[9'h1ab/* 427*/:9'h1a9/* 425*/];
  assign T806 = T807;
  assign T807 = T808;
  assign T808 = T812[T809];
  assign T809 = T810;
  assign T810 = T811;
  assign T811 = io_chanxy_config[8'hcb/* 203*/:8'hca/* 202*/];
  assign T812 = T813;
  assign T813 = io_chanxy_in[9'h1ae/* 430*/:9'h1ac/* 428*/];
  assign T814 = T815;
  assign T815 = T816;
  assign T816 = T820[T817];
  assign T817 = T818;
  assign T818 = T819;
  assign T819 = io_chanxy_config[8'hcd/* 205*/:8'hcc/* 204*/];
  assign T820 = T821;
  assign T821 = io_chanxy_in[9'h1b1/* 433*/:9'h1af/* 431*/];
  assign T822 = T823;
  assign T823 = T824;
  assign T824 = T828[T825];
  assign T825 = T826;
  assign T826 = T827;
  assign T827 = io_chanxy_config[8'hcf/* 207*/:8'hce/* 206*/];
  assign T828 = T829;
  assign T829 = io_chanxy_in[9'h1b4/* 436*/:9'h1b2/* 434*/];
  assign T830 = T831;
  assign T831 = T832;
  assign T832 = T836[T833];
  assign T833 = T834;
  assign T834 = T835;
  assign T835 = io_chanxy_config[8'hd1/* 209*/:8'hd0/* 208*/];
  assign T836 = T837;
  assign T837 = io_chanxy_in[9'h1b7/* 439*/:9'h1b5/* 437*/];
  assign T838 = T839;
  assign T839 = T840;
  assign T840 = T844[T841];
  assign T841 = T842;
  assign T842 = T843;
  assign T843 = io_chanxy_config[8'hd2/* 210*/:8'hd2/* 210*/];
  assign T844 = T845;
  assign T845 = io_chanxy_in[9'h1b9/* 441*/:9'h1b8/* 440*/];
  assign T846 = T847;
  assign T847 = T848;
  assign T848 = T852[T849];
  assign T849 = T850;
  assign T850 = T851;
  assign T851 = io_chanxy_config[8'hd3/* 211*/:8'hd3/* 211*/];
  assign T852 = T853;
  assign T853 = io_chanxy_in[9'h1bb/* 443*/:9'h1ba/* 442*/];
  assign T854 = T855;
  assign T855 = T856;
  assign T856 = T860[T857];
  assign T857 = T858;
  assign T858 = T859;
  assign T859 = io_chanxy_config[8'hd4/* 212*/:8'hd4/* 212*/];
  assign T860 = T861;
  assign T861 = io_chanxy_in[9'h1bd/* 445*/:9'h1bc/* 444*/];
  assign T862 = T863;
  assign T863 = T864;
  assign T864 = T868[T865];
  assign T865 = T866;
  assign T866 = T867;
  assign T867 = io_chanxy_config[8'hd5/* 213*/:8'hd5/* 213*/];
  assign T868 = T869;
  assign T869 = io_chanxy_in[9'h1bf/* 447*/:9'h1be/* 446*/];
  assign T870 = T871;
  assign T871 = T872;
  assign T872 = T876[T873];
  assign T873 = T874;
  assign T874 = T875;
  assign T875 = io_chanxy_config[8'hd6/* 214*/:8'hd6/* 214*/];
  assign T876 = T877;
  assign T877 = io_chanxy_in[9'h1c1/* 449*/:9'h1c0/* 448*/];
  assign T878 = T879;
  assign T879 = T880;
  assign T880 = T884[T881];
  assign T881 = T882;
  assign T882 = T883;
  assign T883 = io_chanxy_config[8'hd7/* 215*/:8'hd7/* 215*/];
  assign T884 = T885;
  assign T885 = io_chanxy_in[9'h1c3/* 451*/:9'h1c2/* 450*/];
  assign T886 = T887;
  assign T887 = T888;
  assign T888 = T892[T889];
  assign T889 = T890;
  assign T890 = T891;
  assign T891 = io_chanxy_config[8'hd8/* 216*/:8'hd8/* 216*/];
  assign T892 = T893;
  assign T893 = io_chanxy_in[9'h1c5/* 453*/:9'h1c4/* 452*/];
  assign T894 = T895;
  assign T895 = T896;
  assign T896 = T900[T897];
  assign T897 = T898;
  assign T898 = T899;
  assign T899 = io_chanxy_config[8'hd9/* 217*/:8'hd9/* 217*/];
  assign T900 = T901;
  assign T901 = io_chanxy_in[9'h1c7/* 455*/:9'h1c6/* 454*/];
  assign T902 = T903;
  assign T903 = T904;
  assign T904 = T908[T905];
  assign T905 = T906;
  assign T906 = T907;
  assign T907 = io_chanxy_config[8'hda/* 218*/:8'hda/* 218*/];
  assign T908 = T909;
  assign T909 = io_chanxy_in[9'h1c9/* 457*/:9'h1c8/* 456*/];
  assign T910 = T911;
  assign T911 = T912;
  assign T912 = T916[T913];
  assign T913 = T914;
  assign T914 = T915;
  assign T915 = io_chanxy_config[8'hdb/* 219*/:8'hdb/* 219*/];
  assign T916 = T917;
  assign T917 = io_chanxy_in[9'h1cb/* 459*/:9'h1ca/* 458*/];
  assign T918 = T919;
  assign T919 = T920;
  assign T920 = T924[T921];
  assign T921 = T922;
  assign T922 = T923;
  assign T923 = io_chanxy_config[8'hdd/* 221*/:8'hdc/* 220*/];
  assign T924 = T925;
  assign T925 = io_chanxy_in[9'h1ce/* 462*/:9'h1cc/* 460*/];
  assign T926 = T927;
  assign T927 = T928;
  assign T928 = T932[T929];
  assign T929 = T930;
  assign T930 = T931;
  assign T931 = io_chanxy_config[8'hdf/* 223*/:8'hde/* 222*/];
  assign T932 = T933;
  assign T933 = io_chanxy_in[9'h1d1/* 465*/:9'h1cf/* 463*/];
  assign T934 = T935;
  assign T935 = T936;
  assign T936 = T940[T937];
  assign T937 = T938;
  assign T938 = T939;
  assign T939 = io_chanxy_config[8'he1/* 225*/:8'he0/* 224*/];
  assign T940 = T941;
  assign T941 = io_chanxy_in[9'h1d4/* 468*/:9'h1d2/* 466*/];
  assign T942 = T943;
  assign T943 = T944;
  assign T944 = T948[T945];
  assign T945 = T946;
  assign T946 = T947;
  assign T947 = io_chanxy_config[8'he3/* 227*/:8'he2/* 226*/];
  assign T948 = T949;
  assign T949 = io_chanxy_in[9'h1d7/* 471*/:9'h1d5/* 469*/];
  assign T950 = T951;
  assign T951 = T952;
  assign T952 = T956[T953];
  assign T953 = T954;
  assign T954 = T955;
  assign T955 = io_chanxy_config[8'he5/* 229*/:8'he4/* 228*/];
  assign T956 = T957;
  assign T957 = io_chanxy_in[9'h1da/* 474*/:9'h1d8/* 472*/];
  assign T958 = T959;
  assign T959 = T960;
  assign T960 = T964[T961];
  assign T961 = T962;
  assign T962 = T963;
  assign T963 = io_chanxy_config[8'he7/* 231*/:8'he6/* 230*/];
  assign T964 = T965;
  assign T965 = io_chanxy_in[9'h1dd/* 477*/:9'h1db/* 475*/];
  assign T966 = T967;
  assign T967 = T968;
  assign T968 = T972[T969];
  assign T969 = T970;
  assign T970 = T971;
  assign T971 = io_chanxy_config[8'he9/* 233*/:8'he8/* 232*/];
  assign T972 = T973;
  assign T973 = io_chanxy_in[9'h1e0/* 480*/:9'h1de/* 478*/];
  assign T974 = T975;
  assign T975 = T976;
  assign T976 = T980[T977];
  assign T977 = T978;
  assign T978 = T979;
  assign T979 = io_chanxy_config[8'heb/* 235*/:8'hea/* 234*/];
  assign T980 = T981;
  assign T981 = io_chanxy_in[9'h1e3/* 483*/:9'h1e1/* 481*/];
  assign T982 = T983;
  assign T983 = T984;
  assign T984 = T988[T985];
  assign T985 = T986;
  assign T986 = T987;
  assign T987 = io_chanxy_config[8'hed/* 237*/:8'hec/* 236*/];
  assign T988 = T989;
  assign T989 = io_chanxy_in[9'h1e6/* 486*/:9'h1e4/* 484*/];
  assign T990 = T991;
  assign T991 = T992;
  assign T992 = T996[T993];
  assign T993 = T994;
  assign T994 = T995;
  assign T995 = io_chanxy_config[8'hef/* 239*/:8'hee/* 238*/];
  assign T996 = T997;
  assign T997 = io_chanxy_in[9'h1e9/* 489*/:9'h1e7/* 487*/];
  assign T998 = T999;
  assign T999 = T1000;
  assign T1000 = T1004[T1001];
  assign T1001 = T1002;
  assign T1002 = T1003;
  assign T1003 = io_chanxy_config[8'hf0/* 240*/:8'hf0/* 240*/];
  assign T1004 = T1005;
  assign T1005 = io_chanxy_in[9'h1eb/* 491*/:9'h1ea/* 490*/];
  assign T1006 = T1007;
  assign T1007 = T1008;
  assign T1008 = T1012[T1009];
  assign T1009 = T1010;
  assign T1010 = T1011;
  assign T1011 = io_chanxy_config[8'hf1/* 241*/:8'hf1/* 241*/];
  assign T1012 = T1013;
  assign T1013 = io_chanxy_in[9'h1ed/* 493*/:9'h1ec/* 492*/];
  assign T1014 = T1015;
  assign T1015 = T1016;
  assign T1016 = T1020[T1017];
  assign T1017 = T1018;
  assign T1018 = T1019;
  assign T1019 = io_chanxy_config[8'hf2/* 242*/:8'hf2/* 242*/];
  assign T1020 = T1021;
  assign T1021 = io_chanxy_in[9'h1ef/* 495*/:9'h1ee/* 494*/];
  assign T1022 = T1023;
  assign T1023 = T1024;
  assign T1024 = T1028[T1025];
  assign T1025 = T1026;
  assign T1026 = T1027;
  assign T1027 = io_chanxy_config[8'hf3/* 243*/:8'hf3/* 243*/];
  assign T1028 = T1029;
  assign T1029 = io_chanxy_in[9'h1f1/* 497*/:9'h1f0/* 496*/];
  assign T1030 = T1031;
  assign T1031 = T1032;
  assign T1032 = T1036[T1033];
  assign T1033 = T1034;
  assign T1034 = T1035;
  assign T1035 = io_chanxy_config[8'hf4/* 244*/:8'hf4/* 244*/];
  assign T1036 = T1037;
  assign T1037 = io_chanxy_in[9'h1f3/* 499*/:9'h1f2/* 498*/];
  assign T1038 = T1039;
  assign T1039 = T1040;
  assign T1040 = T1044[T1041];
  assign T1041 = T1042;
  assign T1042 = T1043;
  assign T1043 = io_chanxy_config[8'hf5/* 245*/:8'hf5/* 245*/];
  assign T1044 = T1045;
  assign T1045 = io_chanxy_in[9'h1f5/* 501*/:9'h1f4/* 500*/];
  assign T1046 = T1047;
  assign T1047 = T1048;
  assign T1048 = T1052[T1049];
  assign T1049 = T1050;
  assign T1050 = T1051;
  assign T1051 = io_chanxy_config[8'hf6/* 246*/:8'hf6/* 246*/];
  assign T1052 = T1053;
  assign T1053 = io_chanxy_in[9'h1f7/* 503*/:9'h1f6/* 502*/];
  assign T1054 = T1055;
  assign T1055 = T1056;
  assign T1056 = T1060[T1057];
  assign T1057 = T1058;
  assign T1058 = T1059;
  assign T1059 = io_chanxy_config[8'hf7/* 247*/:8'hf7/* 247*/];
  assign T1060 = T1061;
  assign T1061 = io_chanxy_in[9'h1f9/* 505*/:9'h1f8/* 504*/];
  assign T1062 = T1063;
  assign T1063 = T1064;
  assign T1064 = T1068[T1065];
  assign T1065 = T1066;
  assign T1066 = T1067;
  assign T1067 = io_chanxy_config[8'hf8/* 248*/:8'hf8/* 248*/];
  assign T1068 = T1069;
  assign T1069 = io_chanxy_in[9'h1fb/* 507*/:9'h1fa/* 506*/];
  assign T1070 = T1071;
  assign T1071 = T1072;
  assign T1072 = T1076[T1073];
  assign T1073 = T1074;
  assign T1074 = T1075;
  assign T1075 = io_chanxy_config[8'hf9/* 249*/:8'hf9/* 249*/];
  assign T1076 = T1077;
  assign T1077 = io_chanxy_in[9'h1fd/* 509*/:9'h1fc/* 508*/];
  assign T1078 = T1079;
  assign T1079 = T1080;
  assign T1080 = T1084[T1081];
  assign T1081 = T1082;
  assign T1082 = T1083;
  assign T1083 = io_chanxy_config[8'hfd/* 253*/:8'hfa/* 250*/];
  assign T1084 = T1085;
  assign T1085 = io_chanxy_in[10'h208/* 520*/:9'h1fe/* 510*/];
  assign T1086 = T1087;
  assign T1087 = T1088;
  assign T1088 = T1092[T1089];
  assign T1089 = T1090;
  assign T1090 = T1091;
  assign T1091 = io_chanxy_config[8'hff/* 255*/:8'hfe/* 254*/];
  assign T1092 = T1093;
  assign T1093 = io_chanxy_in[10'h20b/* 523*/:10'h209/* 521*/];
  assign T1094 = T1095;
  assign T1095 = T1096;
  assign T1096 = T1100[T1097];
  assign T1097 = T1098;
  assign T1098 = T1099;
  assign T1099 = io_chanxy_config[9'h103/* 259*/:9'h100/* 256*/];
  assign T1100 = T1101;
  assign T1101 = io_chanxy_in[10'h216/* 534*/:10'h20c/* 524*/];
  assign T1102 = T1103;
  assign T1103 = T1104;
  assign T1104 = T1108[T1105];
  assign T1105 = T1106;
  assign T1106 = T1107;
  assign T1107 = io_chanxy_config[9'h105/* 261*/:9'h104/* 260*/];
  assign T1108 = T1109;
  assign T1109 = io_chanxy_in[10'h219/* 537*/:10'h217/* 535*/];
  assign T1110 = T1111;
  assign T1111 = T1112;
  assign T1112 = T1116[T1113];
  assign T1113 = T1114;
  assign T1114 = T1115;
  assign T1115 = io_chanxy_config[9'h109/* 265*/:9'h106/* 262*/];
  assign T1116 = T1117;
  assign T1117 = io_chanxy_in[10'h224/* 548*/:10'h21a/* 538*/];
  assign T1118 = T1119;
  assign T1119 = T1120;
  assign T1120 = T1124[T1121];
  assign T1121 = T1122;
  assign T1122 = T1123;
  assign T1123 = io_chanxy_config[9'h10b/* 267*/:9'h10a/* 266*/];
  assign T1124 = T1125;
  assign T1125 = io_chanxy_in[10'h227/* 551*/:10'h225/* 549*/];
  assign T1126 = T1127;
  assign T1127 = T1128;
  assign T1128 = T1132[T1129];
  assign T1129 = T1130;
  assign T1130 = T1131;
  assign T1131 = io_chanxy_config[9'h10f/* 271*/:9'h10c/* 268*/];
  assign T1132 = T1133;
  assign T1133 = io_chanxy_in[10'h232/* 562*/:10'h228/* 552*/];
  assign T1134 = T1135;
  assign T1135 = T1136;
  assign T1136 = T1140[T1137];
  assign T1137 = T1138;
  assign T1138 = T1139;
  assign T1139 = io_chanxy_config[9'h111/* 273*/:9'h110/* 272*/];
  assign T1140 = T1141;
  assign T1141 = io_chanxy_in[10'h235/* 565*/:10'h233/* 563*/];
  assign T1142 = T1143;
  assign T1143 = T1144;
  assign T1144 = T1148[T1145];
  assign T1145 = T1146;
  assign T1146 = T1147;
  assign T1147 = io_chanxy_config[9'h115/* 277*/:9'h112/* 274*/];
  assign T1148 = T1149;
  assign T1149 = io_chanxy_in[10'h240/* 576*/:10'h236/* 566*/];
  assign T1150 = T1151;
  assign T1151 = T1152;
  assign T1152 = T1156[T1153];
  assign T1153 = T1154;
  assign T1154 = T1155;
  assign T1155 = io_chanxy_config[9'h117/* 279*/:9'h116/* 278*/];
  assign T1156 = T1157;
  assign T1157 = io_chanxy_in[10'h243/* 579*/:10'h241/* 577*/];
  assign T1158 = T1159;
  assign T1159 = T1160;
  assign T1160 = T1164[T1161];
  assign T1161 = T1162;
  assign T1162 = T1163;
  assign T1163 = io_chanxy_config[9'h11b/* 283*/:9'h118/* 280*/];
  assign T1164 = T1165;
  assign T1165 = io_chanxy_in[10'h24e/* 590*/:10'h244/* 580*/];
  assign T1166 = T1167;
  assign T1167 = T1168;
  assign T1168 = T1172[T1169];
  assign T1169 = T1170;
  assign T1170 = T1171;
  assign T1171 = io_chanxy_config[9'h11d/* 285*/:9'h11c/* 284*/];
  assign T1172 = T1173;
  assign T1173 = io_chanxy_in[10'h251/* 593*/:10'h24f/* 591*/];
  assign T1174 = T1175;
  assign T1175 = T1176;
  assign T1176 = T1180[T1177];
  assign T1177 = T1178;
  assign T1178 = T1179;
  assign T1179 = io_chanxy_config[9'h121/* 289*/:9'h11e/* 286*/];
  assign T1180 = T1181;
  assign T1181 = io_chanxy_in[10'h25c/* 604*/:10'h252/* 594*/];
  assign T1182 = T1183;
  assign T1183 = T1184;
  assign T1184 = T1188[T1185];
  assign T1185 = T1186;
  assign T1186 = T1187;
  assign T1187 = io_chanxy_config[9'h123/* 291*/:9'h122/* 290*/];
  assign T1188 = T1189;
  assign T1189 = io_chanxy_in[10'h25f/* 607*/:10'h25d/* 605*/];
  assign T1190 = T1191;
  assign T1191 = T1192;
  assign T1192 = T1196[T1193];
  assign T1193 = T1194;
  assign T1194 = T1195;
  assign T1195 = io_chanxy_config[9'h127/* 295*/:9'h124/* 292*/];
  assign T1196 = T1197;
  assign T1197 = io_chanxy_in[10'h26a/* 618*/:10'h260/* 608*/];
  assign T1198 = T1199;
  assign T1199 = T1200;
  assign T1200 = T1204[T1201];
  assign T1201 = T1202;
  assign T1202 = T1203;
  assign T1203 = io_chanxy_config[9'h129/* 297*/:9'h128/* 296*/];
  assign T1204 = T1205;
  assign T1205 = io_chanxy_in[10'h26d/* 621*/:10'h26b/* 619*/];
  assign T1206 = T1207;
  assign T1207 = T1208;
  assign T1208 = T1212[T1209];
  assign T1209 = T1210;
  assign T1210 = T1211;
  assign T1211 = io_chanxy_config[9'h12d/* 301*/:9'h12a/* 298*/];
  assign T1212 = T1213;
  assign T1213 = io_chanxy_in[10'h278/* 632*/:10'h26e/* 622*/];
  assign T1214 = T1215;
  assign T1215 = T1216;
  assign T1216 = T1220[T1217];
  assign T1217 = T1218;
  assign T1218 = T1219;
  assign T1219 = io_chanxy_config[9'h12f/* 303*/:9'h12e/* 302*/];
  assign T1220 = T1221;
  assign T1221 = io_chanxy_in[10'h27b/* 635*/:10'h279/* 633*/];
  assign T1222 = T1223;
  assign T1223 = T1224;
  assign T1224 = T1228[T1225];
  assign T1225 = T1226;
  assign T1226 = T1227;
  assign T1227 = io_chanxy_config[9'h133/* 307*/:9'h130/* 304*/];
  assign T1228 = T1229;
  assign T1229 = io_chanxy_in[10'h286/* 646*/:10'h27c/* 636*/];
  assign T1230 = T1231;
  assign T1231 = T1232;
  assign T1232 = T1236[T1233];
  assign T1233 = T1234;
  assign T1234 = T1235;
  assign T1235 = io_chanxy_config[9'h135/* 309*/:9'h134/* 308*/];
  assign T1236 = T1237;
  assign T1237 = io_chanxy_in[10'h289/* 649*/:10'h287/* 647*/];
  assign T1238 = T1239;
  assign T1239 = T1240;
  assign T1240 = T1244[T1241];
  assign T1241 = T1242;
  assign T1242 = T1243;
  assign T1243 = io_chanxy_config[9'h139/* 313*/:9'h136/* 310*/];
  assign T1244 = T1245;
  assign T1245 = io_chanxy_in[10'h294/* 660*/:10'h28a/* 650*/];
  assign T1246 = T1247;
  assign T1247 = T1248;
  assign T1248 = T1252[T1249];
  assign T1249 = T1250;
  assign T1250 = T1251;
  assign T1251 = io_chanxy_config[9'h13a/* 314*/:9'h13a/* 314*/];
  assign T1252 = T1253;
  assign T1253 = io_chanxy_in[10'h296/* 662*/:10'h295/* 661*/];
  assign T1254 = T1255;
  assign T1255 = T1256;
  assign T1256 = T1260[T1257];
  assign T1257 = T1258;
  assign T1258 = T1259;
  assign T1259 = io_chanxy_config[9'h13e/* 318*/:9'h13b/* 315*/];
  assign T1260 = T1261;
  assign T1261 = io_chanxy_in[10'h2a1/* 673*/:10'h297/* 663*/];
  assign T1262 = T1263;
  assign T1263 = T1264;
  assign T1264 = T1268[T1265];
  assign T1265 = T1266;
  assign T1266 = T1267;
  assign T1267 = io_chanxy_config[9'h13f/* 319*/:9'h13f/* 319*/];
  assign T1268 = T1269;
  assign T1269 = io_chanxy_in[10'h2a3/* 675*/:10'h2a2/* 674*/];
  assign T1270 = T1271;
  assign T1271 = T1272;
  assign T1272 = T1276[T1273];
  assign T1273 = T1274;
  assign T1274 = T1275;
  assign T1275 = io_chanxy_config[9'h143/* 323*/:9'h140/* 320*/];
  assign T1276 = T1277;
  assign T1277 = io_chanxy_in[10'h2ae/* 686*/:10'h2a4/* 676*/];
  assign T1278 = T1279;
  assign T1279 = T1280;
  assign T1280 = T1284[T1281];
  assign T1281 = T1282;
  assign T1282 = T1283;
  assign T1283 = io_chanxy_config[9'h144/* 324*/:9'h144/* 324*/];
  assign T1284 = T1285;
  assign T1285 = io_chanxy_in[10'h2b0/* 688*/:10'h2af/* 687*/];
  assign T1286 = T1287;
  assign T1287 = T1288;
  assign T1288 = T1292[T1289];
  assign T1289 = T1290;
  assign T1290 = T1291;
  assign T1291 = io_chanxy_config[9'h148/* 328*/:9'h145/* 325*/];
  assign T1292 = T1293;
  assign T1293 = io_chanxy_in[10'h2bb/* 699*/:10'h2b1/* 689*/];
  assign T1294 = T1295;
  assign T1295 = T1296;
  assign T1296 = T1300[T1297];
  assign T1297 = T1298;
  assign T1298 = T1299;
  assign T1299 = io_chanxy_config[9'h149/* 329*/:9'h149/* 329*/];
  assign T1300 = T1301;
  assign T1301 = io_chanxy_in[10'h2bd/* 701*/:10'h2bc/* 700*/];
  assign T1302 = T1303;
  assign T1303 = T1304;
  assign T1304 = T1308[T1305];
  assign T1305 = T1306;
  assign T1306 = T1307;
  assign T1307 = io_chanxy_config[9'h14d/* 333*/:9'h14a/* 330*/];
  assign T1308 = T1309;
  assign T1309 = io_chanxy_in[10'h2c8/* 712*/:10'h2be/* 702*/];
  assign T1310 = T1311;
  assign T1311 = T1312;
  assign T1312 = T1316[T1313];
  assign T1313 = T1314;
  assign T1314 = T1315;
  assign T1315 = io_chanxy_config[9'h14e/* 334*/:9'h14e/* 334*/];
  assign T1316 = T1317;
  assign T1317 = io_chanxy_in[10'h2ca/* 714*/:10'h2c9/* 713*/];
  assign T1318 = T1319;
  assign T1319 = T1320;
  assign T1320 = T1324[T1321];
  assign T1321 = T1322;
  assign T1322 = T1323;
  assign T1323 = io_chanxy_config[9'h152/* 338*/:9'h14f/* 335*/];
  assign T1324 = T1325;
  assign T1325 = io_chanxy_in[10'h2d5/* 725*/:10'h2cb/* 715*/];
  assign T1326 = T1327;
  assign T1327 = T1328;
  assign T1328 = T1332[T1329];
  assign T1329 = T1330;
  assign T1330 = T1331;
  assign T1331 = io_chanxy_config[9'h153/* 339*/:9'h153/* 339*/];
  assign T1332 = T1333;
  assign T1333 = io_chanxy_in[10'h2d7/* 727*/:10'h2d6/* 726*/];
  assign T1334 = T1335;
  assign T1335 = T1336;
  assign T1336 = T1340[T1337];
  assign T1337 = T1338;
  assign T1338 = T1339;
  assign T1339 = io_chanxy_config[9'h157/* 343*/:9'h154/* 340*/];
  assign T1340 = T1341;
  assign T1341 = io_chanxy_in[10'h2e2/* 738*/:10'h2d8/* 728*/];
  assign T1342 = T1343;
  assign T1343 = T1344;
  assign T1344 = T1348[T1345];
  assign T1345 = T1346;
  assign T1346 = T1347;
  assign T1347 = io_chanxy_config[9'h158/* 344*/:9'h158/* 344*/];
  assign T1348 = T1349;
  assign T1349 = io_chanxy_in[10'h2e4/* 740*/:10'h2e3/* 739*/];
  assign T1350 = T1351;
  assign T1351 = T1352;
  assign T1352 = T1356[T1353];
  assign T1353 = T1354;
  assign T1354 = T1355;
  assign T1355 = io_chanxy_config[9'h15c/* 348*/:9'h159/* 345*/];
  assign T1356 = T1357;
  assign T1357 = io_chanxy_in[10'h2ef/* 751*/:10'h2e5/* 741*/];
  assign T1358 = T1359;
  assign T1359 = T1360;
  assign T1360 = T1364[T1361];
  assign T1361 = T1362;
  assign T1362 = T1363;
  assign T1363 = io_chanxy_config[9'h15d/* 349*/:9'h15d/* 349*/];
  assign T1364 = T1365;
  assign T1365 = io_chanxy_in[10'h2f1/* 753*/:10'h2f0/* 752*/];
  assign T1366 = T1367;
  assign T1367 = T1368;
  assign T1368 = T1372[T1369];
  assign T1369 = T1370;
  assign T1370 = T1371;
  assign T1371 = io_chanxy_config[9'h161/* 353*/:9'h15e/* 350*/];
  assign T1372 = T1373;
  assign T1373 = io_chanxy_in[10'h2fc/* 764*/:10'h2f2/* 754*/];
  assign T1374 = T1375;
  assign T1375 = T1376;
  assign T1376 = T1380[T1377];
  assign T1377 = T1378;
  assign T1378 = T1379;
  assign T1379 = io_chanxy_config[9'h162/* 354*/:9'h162/* 354*/];
  assign T1380 = T1381;
  assign T1381 = io_chanxy_in[10'h2fe/* 766*/:10'h2fd/* 765*/];
  assign T1382 = T1383;
  assign T1383 = T1384;
  assign T1384 = T1388[T1385];
  assign T1385 = T1386;
  assign T1386 = T1387;
  assign T1387 = io_chanxy_config[9'h166/* 358*/:9'h163/* 355*/];
  assign T1388 = T1389;
  assign T1389 = io_chanxy_in[10'h309/* 777*/:10'h2ff/* 767*/];
  assign T1390 = T1391;
  assign T1391 = T1392;
  assign T1392 = T1396[T1393];
  assign T1393 = T1394;
  assign T1394 = T1395;
  assign T1395 = io_chanxy_config[9'h167/* 359*/:9'h167/* 359*/];
  assign T1396 = T1397;
  assign T1397 = io_chanxy_in[10'h30b/* 779*/:10'h30a/* 778*/];
  assign io_ipin_out = T1398;
  assign T1398 = T1399;
  assign T1399 = {T1718, T1400};
  assign T1400 = T1401;
  assign T1401 = {T1710, T1402};
  assign T1402 = T1403;
  assign T1403 = {T1702, T1404};
  assign T1404 = T1405;
  assign T1405 = {T1694, T1406};
  assign T1406 = T1407;
  assign T1407 = {T1686, T1408};
  assign T1408 = T1409;
  assign T1409 = {T1678, T1410};
  assign T1410 = T1411;
  assign T1411 = {T1670, T1412};
  assign T1412 = T1413;
  assign T1413 = {T1662, T1414};
  assign T1414 = T1415;
  assign T1415 = {T1654, T1416};
  assign T1416 = T1417;
  assign T1417 = {T1646, T1418};
  assign T1418 = T1419;
  assign T1419 = {T1638, T1420};
  assign T1420 = T1421;
  assign T1421 = {T1630, T1422};
  assign T1422 = T1423;
  assign T1423 = {T1622, T1424};
  assign T1424 = T1425;
  assign T1425 = {T1614, T1426};
  assign T1426 = T1427;
  assign T1427 = {T1606, T1428};
  assign T1428 = T1429;
  assign T1429 = {T1598, T1430};
  assign T1430 = T1431;
  assign T1431 = {T1590, T1432};
  assign T1432 = T1433;
  assign T1433 = {T1582, T1434};
  assign T1434 = T1435;
  assign T1435 = {T1574, T1436};
  assign T1436 = T1437;
  assign T1437 = {T1566, T1438};
  assign T1438 = T1439;
  assign T1439 = {T1558, T1440};
  assign T1440 = T1441;
  assign T1441 = {T1550, T1442};
  assign T1442 = T1443;
  assign T1443 = {T1542, T1444};
  assign T1444 = T1445;
  assign T1445 = {T1534, T1446};
  assign T1446 = T1447;
  assign T1447 = {T1526, T1448};
  assign T1448 = T1449;
  assign T1449 = {T1518, T1450};
  assign T1450 = T1451;
  assign T1451 = {T1510, T1452};
  assign T1452 = T1453;
  assign T1453 = {T1502, T1454};
  assign T1454 = T1455;
  assign T1455 = {T1494, T1456};
  assign T1456 = T1457;
  assign T1457 = {T1486, T1458};
  assign T1458 = T1459;
  assign T1459 = {T1478, T1460};
  assign T1460 = T1461;
  assign T1461 = {T1470, T1462};
  assign T1462 = T1463;
  assign T1463 = T1464;
  assign T1464 = T1468[T1465];
  assign T1465 = T1466;
  assign T1466 = T1467;
  assign T1467 = io_ipin_config[2'h3/* 3*/:1'h0/* 0*/];
  assign T1468 = T1469;
  assign T1469 = io_ipin_in[4'hf/* 15*/:1'h0/* 0*/];
  assign T1470 = T1471;
  assign T1471 = T1472;
  assign T1472 = T1476[T1473];
  assign T1473 = T1474;
  assign T1474 = T1475;
  assign T1475 = io_ipin_config[3'h7/* 7*/:3'h4/* 4*/];
  assign T1476 = T1477;
  assign T1477 = io_ipin_in[5'h1f/* 31*/:5'h10/* 16*/];
  assign T1478 = T1479;
  assign T1479 = T1480;
  assign T1480 = T1484[T1481];
  assign T1481 = T1482;
  assign T1482 = T1483;
  assign T1483 = io_ipin_config[4'hb/* 11*/:4'h8/* 8*/];
  assign T1484 = T1485;
  assign T1485 = io_ipin_in[6'h2f/* 47*/:6'h20/* 32*/];
  assign T1486 = T1487;
  assign T1487 = T1488;
  assign T1488 = T1492[T1489];
  assign T1489 = T1490;
  assign T1490 = T1491;
  assign T1491 = io_ipin_config[4'hf/* 15*/:4'hc/* 12*/];
  assign T1492 = T1493;
  assign T1493 = io_ipin_in[6'h3f/* 63*/:6'h30/* 48*/];
  assign T1494 = T1495;
  assign T1495 = T1496;
  assign T1496 = T1500[T1497];
  assign T1497 = T1498;
  assign T1498 = T1499;
  assign T1499 = io_ipin_config[5'h13/* 19*/:5'h10/* 16*/];
  assign T1500 = T1501;
  assign T1501 = io_ipin_in[7'h4f/* 79*/:7'h40/* 64*/];
  assign T1502 = T1503;
  assign T1503 = T1504;
  assign T1504 = T1508[T1505];
  assign T1505 = T1506;
  assign T1506 = T1507;
  assign T1507 = io_ipin_config[5'h17/* 23*/:5'h14/* 20*/];
  assign T1508 = T1509;
  assign T1509 = io_ipin_in[7'h5f/* 95*/:7'h50/* 80*/];
  assign T1510 = T1511;
  assign T1511 = T1512;
  assign T1512 = T1516[T1513];
  assign T1513 = T1514;
  assign T1514 = T1515;
  assign T1515 = io_ipin_config[5'h1b/* 27*/:5'h18/* 24*/];
  assign T1516 = T1517;
  assign T1517 = io_ipin_in[7'h6f/* 111*/:7'h60/* 96*/];
  assign T1518 = T1519;
  assign T1519 = T1520;
  assign T1520 = T1524[T1521];
  assign T1521 = T1522;
  assign T1522 = T1523;
  assign T1523 = io_ipin_config[5'h1f/* 31*/:5'h1c/* 28*/];
  assign T1524 = T1525;
  assign T1525 = io_ipin_in[7'h7f/* 127*/:7'h70/* 112*/];
  assign T1526 = T1527;
  assign T1527 = T1528;
  assign T1528 = T1532[T1529];
  assign T1529 = T1530;
  assign T1530 = T1531;
  assign T1531 = io_ipin_config[6'h23/* 35*/:6'h20/* 32*/];
  assign T1532 = T1533;
  assign T1533 = io_ipin_in[8'h8f/* 143*/:8'h80/* 128*/];
  assign T1534 = T1535;
  assign T1535 = T1536;
  assign T1536 = T1540[T1537];
  assign T1537 = T1538;
  assign T1538 = T1539;
  assign T1539 = io_ipin_config[6'h27/* 39*/:6'h24/* 36*/];
  assign T1540 = T1541;
  assign T1541 = io_ipin_in[8'h9f/* 159*/:8'h90/* 144*/];
  assign T1542 = T1543;
  assign T1543 = T1544;
  assign T1544 = T1548[T1545];
  assign T1545 = T1546;
  assign T1546 = T1547;
  assign T1547 = io_ipin_config[6'h2b/* 43*/:6'h28/* 40*/];
  assign T1548 = T1549;
  assign T1549 = io_ipin_in[8'haf/* 175*/:8'ha0/* 160*/];
  assign T1550 = T1551;
  assign T1551 = T1552;
  assign T1552 = T1556[T1553];
  assign T1553 = T1554;
  assign T1554 = T1555;
  assign T1555 = io_ipin_config[6'h2f/* 47*/:6'h2c/* 44*/];
  assign T1556 = T1557;
  assign T1557 = io_ipin_in[8'hbf/* 191*/:8'hb0/* 176*/];
  assign T1558 = T1559;
  assign T1559 = T1560;
  assign T1560 = T1564[T1561];
  assign T1561 = T1562;
  assign T1562 = T1563;
  assign T1563 = io_ipin_config[6'h33/* 51*/:6'h30/* 48*/];
  assign T1564 = T1565;
  assign T1565 = io_ipin_in[8'hcf/* 207*/:8'hc0/* 192*/];
  assign T1566 = T1567;
  assign T1567 = T1568;
  assign T1568 = T1572[T1569];
  assign T1569 = T1570;
  assign T1570 = T1571;
  assign T1571 = io_ipin_config[6'h37/* 55*/:6'h34/* 52*/];
  assign T1572 = T1573;
  assign T1573 = io_ipin_in[8'hdf/* 223*/:8'hd0/* 208*/];
  assign T1574 = T1575;
  assign T1575 = T1576;
  assign T1576 = T1580[T1577];
  assign T1577 = T1578;
  assign T1578 = T1579;
  assign T1579 = io_ipin_config[6'h3b/* 59*/:6'h38/* 56*/];
  assign T1580 = T1581;
  assign T1581 = io_ipin_in[8'hef/* 239*/:8'he0/* 224*/];
  assign T1582 = T1583;
  assign T1583 = T1584;
  assign T1584 = T1588[T1585];
  assign T1585 = T1586;
  assign T1586 = T1587;
  assign T1587 = io_ipin_config[6'h3f/* 63*/:6'h3c/* 60*/];
  assign T1588 = T1589;
  assign T1589 = io_ipin_in[8'hff/* 255*/:8'hf0/* 240*/];
  assign T1590 = T1591;
  assign T1591 = T1592;
  assign T1592 = T1596[T1593];
  assign T1593 = T1594;
  assign T1594 = T1595;
  assign T1595 = io_ipin_config[7'h43/* 67*/:7'h40/* 64*/];
  assign T1596 = T1597;
  assign T1597 = io_ipin_in[9'h10f/* 271*/:9'h100/* 256*/];
  assign T1598 = T1599;
  assign T1599 = T1600;
  assign T1600 = T1604[T1601];
  assign T1601 = T1602;
  assign T1602 = T1603;
  assign T1603 = io_ipin_config[7'h47/* 71*/:7'h44/* 68*/];
  assign T1604 = T1605;
  assign T1605 = io_ipin_in[9'h11f/* 287*/:9'h110/* 272*/];
  assign T1606 = T1607;
  assign T1607 = T1608;
  assign T1608 = T1612[T1609];
  assign T1609 = T1610;
  assign T1610 = T1611;
  assign T1611 = io_ipin_config[7'h4b/* 75*/:7'h48/* 72*/];
  assign T1612 = T1613;
  assign T1613 = io_ipin_in[9'h12f/* 303*/:9'h120/* 288*/];
  assign T1614 = T1615;
  assign T1615 = T1616;
  assign T1616 = T1620[T1617];
  assign T1617 = T1618;
  assign T1618 = T1619;
  assign T1619 = io_ipin_config[7'h4f/* 79*/:7'h4c/* 76*/];
  assign T1620 = T1621;
  assign T1621 = io_ipin_in[9'h13f/* 319*/:9'h130/* 304*/];
  assign T1622 = T1623;
  assign T1623 = T1624;
  assign T1624 = T1628[T1625];
  assign T1625 = T1626;
  assign T1626 = T1627;
  assign T1627 = io_ipin_config[7'h53/* 83*/:7'h50/* 80*/];
  assign T1628 = T1629;
  assign T1629 = io_ipin_in[9'h14f/* 335*/:9'h140/* 320*/];
  assign T1630 = T1631;
  assign T1631 = T1632;
  assign T1632 = T1636[T1633];
  assign T1633 = T1634;
  assign T1634 = T1635;
  assign T1635 = io_ipin_config[7'h57/* 87*/:7'h54/* 84*/];
  assign T1636 = T1637;
  assign T1637 = io_ipin_in[9'h15f/* 351*/:9'h150/* 336*/];
  assign T1638 = T1639;
  assign T1639 = T1640;
  assign T1640 = T1644[T1641];
  assign T1641 = T1642;
  assign T1642 = T1643;
  assign T1643 = io_ipin_config[7'h5b/* 91*/:7'h58/* 88*/];
  assign T1644 = T1645;
  assign T1645 = io_ipin_in[9'h16f/* 367*/:9'h160/* 352*/];
  assign T1646 = T1647;
  assign T1647 = T1648;
  assign T1648 = T1652[T1649];
  assign T1649 = T1650;
  assign T1650 = T1651;
  assign T1651 = io_ipin_config[7'h5f/* 95*/:7'h5c/* 92*/];
  assign T1652 = T1653;
  assign T1653 = io_ipin_in[9'h17f/* 383*/:9'h170/* 368*/];
  assign T1654 = T1655;
  assign T1655 = T1656;
  assign T1656 = T1660[T1657];
  assign T1657 = T1658;
  assign T1658 = T1659;
  assign T1659 = io_ipin_config[7'h63/* 99*/:7'h60/* 96*/];
  assign T1660 = T1661;
  assign T1661 = io_ipin_in[9'h18f/* 399*/:9'h180/* 384*/];
  assign T1662 = T1663;
  assign T1663 = T1664;
  assign T1664 = T1668[T1665];
  assign T1665 = T1666;
  assign T1666 = T1667;
  assign T1667 = io_ipin_config[7'h67/* 103*/:7'h64/* 100*/];
  assign T1668 = T1669;
  assign T1669 = io_ipin_in[9'h19f/* 415*/:9'h190/* 400*/];
  assign T1670 = T1671;
  assign T1671 = T1672;
  assign T1672 = T1676[T1673];
  assign T1673 = T1674;
  assign T1674 = T1675;
  assign T1675 = io_ipin_config[7'h6b/* 107*/:7'h68/* 104*/];
  assign T1676 = T1677;
  assign T1677 = io_ipin_in[9'h1af/* 431*/:9'h1a0/* 416*/];
  assign T1678 = T1679;
  assign T1679 = T1680;
  assign T1680 = T1684[T1681];
  assign T1681 = T1682;
  assign T1682 = T1683;
  assign T1683 = io_ipin_config[7'h6f/* 111*/:7'h6c/* 108*/];
  assign T1684 = T1685;
  assign T1685 = io_ipin_in[9'h1bf/* 447*/:9'h1b0/* 432*/];
  assign T1686 = T1687;
  assign T1687 = T1688;
  assign T1688 = T1692[T1689];
  assign T1689 = T1690;
  assign T1690 = T1691;
  assign T1691 = io_ipin_config[7'h73/* 115*/:7'h70/* 112*/];
  assign T1692 = T1693;
  assign T1693 = io_ipin_in[9'h1cf/* 463*/:9'h1c0/* 448*/];
  assign T1694 = T1695;
  assign T1695 = T1696;
  assign T1696 = T1700[T1697];
  assign T1697 = T1698;
  assign T1698 = T1699;
  assign T1699 = io_ipin_config[7'h77/* 119*/:7'h74/* 116*/];
  assign T1700 = T1701;
  assign T1701 = io_ipin_in[9'h1df/* 479*/:9'h1d0/* 464*/];
  assign T1702 = T1703;
  assign T1703 = T1704;
  assign T1704 = T1708[T1705];
  assign T1705 = T1706;
  assign T1706 = T1707;
  assign T1707 = io_ipin_config[7'h7b/* 123*/:7'h78/* 120*/];
  assign T1708 = T1709;
  assign T1709 = io_ipin_in[9'h1ef/* 495*/:9'h1e0/* 480*/];
  assign T1710 = T1711;
  assign T1711 = T1712;
  assign T1712 = T1716[T1713];
  assign T1713 = T1714;
  assign T1714 = T1715;
  assign T1715 = io_ipin_config[7'h7f/* 127*/:7'h7c/* 124*/];
  assign T1716 = T1717;
  assign T1717 = io_ipin_in[9'h1ff/* 511*/:9'h1f0/* 496*/];
  assign T1718 = T1719;
  assign T1719 = T1720;
  assign T1720 = T1724[T1721];
  assign T1721 = T1722;
  assign T1722 = T1723;
  assign T1723 = io_ipin_config[8'h83/* 131*/:8'h80/* 128*/];
  assign T1724 = T1725;
  assign T1725 = io_ipin_in[10'h20f/* 527*/:10'h200/* 512*/];
endmodule

module lut_tile_sp_13(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [779:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h2/* 2*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_11 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_14(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [779:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {6'h0/* 0*/, 2'h3/* 3*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_11 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule

module lut_tile_sp_15(input clk, input reset,
    input  io_ff_en,
    input [31:0] io_configs_in,
    input [46:0] io_configs_en,
    input [527:0] io_ipin_in,
    input [779:0] io_chanxy_in,
    output[139:0] io_chanxy_out,
    output[9:0] io_opin_out,
    output[7:0] io_x_loc,
    output[7:0] io_y_loc);

  wire[359:0] T0;
  wire[1503:0] this_config_io_configs_out;
  wire[131:0] T1;
  wire[359:0] T2;
  wire[42:0] T3;
  wire[32:0] this_sbcb_io_ipin_out;
  wire[9:0] this_clb_io_clb_out;
  wire[9:0] T4;
  wire[639:0] T5;
  wire[59:0] this_xbar_io_xbar_out;
  wire[7:0] T6;
  wire[7:0] T7;
  wire[139:0] this_sbcb_io_chanxy_out;

  assign T0 = this_config_io_configs_out[11'h5dd/* 1501*/:11'h476/* 1142*/];
  assign T1 = this_config_io_configs_out[11'h475/* 1141*/:10'h3f2/* 1010*/];
  assign T2 = this_config_io_configs_out[10'h3f1/* 1009*/:10'h28a/* 650*/];
  assign T3 = {this_clb_io_clb_out, this_sbcb_io_ipin_out};
  assign T4 = this_config_io_configs_out[10'h289/* 649*/:10'h280/* 640*/];
  assign T5 = this_config_io_configs_out[10'h27f/* 639*/:1'h0/* 0*/];
  assign io_y_loc = T6;
  assign T6 = {5'h0/* 0*/, 3'h5/* 5*/};
  assign io_x_loc = T7;
  assign T7 = {5'h0/* 0*/, 3'h4/* 4*/};
  assign io_opin_out = this_clb_io_clb_out;
  assign io_chanxy_out = this_sbcb_io_chanxy_out;
  clb this_clb(.clk(clk), .reset(reset),
       .io_clb_in( this_xbar_io_xbar_out ),
       .io_clb_out( this_clb_io_clb_out ),
       .io_lut_configs( T5 ),
       .io_mux_configs( T4 ),
       .io_ff_en( io_ff_en ));
  xbar this_xbar(.clk(clk), .reset(reset),
       .io_xbar_in( T3 ),
       .io_xbar_out( this_xbar_io_xbar_out ),
       .io_mux_configs( T2 ));
    configs_latches_47 this_config(.clk(clk), .reset(reset),
       .io_d_in( io_configs_in ),
       .io_configs_out( this_config_io_configs_out ),
       .io_configs_en( io_configs_en ));
  sbcb_sp_11 this_sbcb(
       .io_ipin_in( io_ipin_in ),
       .io_ipin_config( T1 ),
       .io_chanxy_in( io_chanxy_in ),
       .io_chanxy_config( T0 ),
       .io_ipin_out( this_sbcb_io_ipin_out ),
       .io_chanxy_out( this_sbcb_io_chanxy_out ));
endmodule


